//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:23 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n700, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XOR2_X1   g001(.A(KEYINPUT95), .B(G36gat), .Z(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT94), .B(G29gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT15), .ZN(new_n206));
  NOR2_X1   g005(.A1(G29gat), .A2(G36gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT14), .ZN(new_n208));
  OR3_X1    g007(.A1(new_n205), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G43gat), .B(G50gat), .ZN(new_n210));
  OR2_X1    g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n206), .B1(new_n205), .B2(new_n208), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n212), .A3(new_n210), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G15gat), .B(G22gat), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT16), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n215), .B1(new_n216), .B2(G1gat), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(G1gat), .B2(new_n215), .ZN(new_n218));
  XOR2_X1   g017(.A(new_n218), .B(G8gat), .Z(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n214), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT17), .ZN(new_n222));
  OAI21_X1  g021(.A(new_n219), .B1(new_n214), .B2(new_n222), .ZN(new_n223));
  XOR2_X1   g022(.A(KEYINPUT96), .B(KEYINPUT17), .Z(new_n224));
  AOI21_X1  g023(.A(new_n224), .B1(new_n211), .B2(new_n213), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n202), .B(new_n221), .C1(new_n223), .C2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT18), .ZN(new_n227));
  OR2_X1    g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n227), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n214), .B(new_n220), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n202), .B(KEYINPUT13), .Z(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G169gat), .B(G197gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT93), .ZN(new_n235));
  INV_X1    g034(.A(G113gat), .ZN(new_n236));
  XNOR2_X1  g035(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n238));
  INV_X1    g037(.A(G141gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n237), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n241), .B(KEYINPUT12), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n233), .A2(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n228), .A2(new_n229), .A3(new_n232), .A4(new_n242), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n244), .A2(KEYINPUT97), .A3(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT97), .B1(new_n244), .B2(new_n245), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(G15gat), .B(G43gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT76), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT77), .ZN(new_n251));
  XOR2_X1   g050(.A(G71gat), .B(G99gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G134gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n254), .A2(G127gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(G127gat), .ZN(new_n258));
  INV_X1    g057(.A(G127gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(G134gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(new_n257), .B1(new_n261), .B2(new_n256), .ZN(new_n262));
  INV_X1    g061(.A(G120gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n236), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(G113gat), .A2(G120gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n266), .A2(KEYINPUT71), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT1), .B1(new_n266), .B2(KEYINPUT71), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n262), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT73), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT73), .B1(new_n258), .B2(new_n260), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AND2_X1   g072(.A1(G113gat), .A2(G120gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(G113gat), .A2(G120gat), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT72), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT72), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n264), .A2(new_n277), .A3(new_n265), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT74), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n273), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT73), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n259), .A2(G134gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(new_n255), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT73), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(KEYINPUT74), .B1(new_n283), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n270), .B1(new_n282), .B2(new_n289), .ZN(new_n290));
  OR2_X1    g089(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n291));
  NAND2_X1  g090(.A1(KEYINPUT68), .A2(KEYINPUT27), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n291), .A2(G183gat), .A3(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n294));
  XNOR2_X1  g093(.A(KEYINPUT67), .B(G183gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT27), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n293), .B(new_n294), .C1(new_n295), .C2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(G169gat), .A2(G176gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT66), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT26), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n302));
  NAND3_X1  g101(.A1(new_n300), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G169gat), .A2(G176gat), .ZN(new_n304));
  INV_X1    g103(.A(G169gat), .ZN(new_n305));
  INV_X1    g104(.A(G176gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n304), .B1(new_n307), .B2(KEYINPUT26), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  AND3_X1   g109(.A1(new_n297), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G190gat), .ZN(new_n312));
  INV_X1    g111(.A(G183gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT27), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n296), .A2(G183gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT69), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n314), .B2(new_n315), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n312), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT24), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n313), .A2(new_n312), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n304), .B1(KEYINPUT23), .B2(new_n298), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT65), .B1(new_n307), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT65), .ZN(new_n330));
  NOR3_X1   g129(.A1(new_n298), .A2(new_n330), .A3(KEYINPUT23), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n326), .B(new_n327), .C1(new_n329), .C2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n333));
  NAND2_X1  g132(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g133(.A(new_n323), .B(new_n324), .C1(new_n295), .C2(G190gat), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT25), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n304), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n307), .A2(KEYINPUT65), .A3(new_n328), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n330), .B1(new_n298), .B2(KEYINPUT23), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n300), .A2(KEYINPUT23), .A3(new_n302), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n335), .A2(new_n337), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n311), .A2(new_n321), .B1(new_n334), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n290), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n334), .A2(new_n342), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n303), .A2(new_n308), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n296), .A2(G183gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n313), .A2(KEYINPUT27), .ZN(new_n348));
  OAI21_X1  g147(.A(KEYINPUT69), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(G190gat), .B1(new_n349), .B2(new_n317), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  OAI211_X1 g150(.A(new_n346), .B(new_n297), .C1(new_n350), .C2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n281), .B1(new_n273), .B2(new_n280), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT1), .B1(new_n266), .B2(KEYINPUT72), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n288), .A2(KEYINPUT74), .A3(new_n355), .A4(new_n278), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n269), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(G227gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n344), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(KEYINPUT75), .B(KEYINPUT33), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n253), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n362), .B(KEYINPUT32), .C1(new_n253), .C2(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n361), .B1(new_n344), .B2(new_n358), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT34), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n368), .A2(KEYINPUT78), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT78), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n367), .B(new_n366), .C1(new_n370), .C2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT36), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n370), .A2(new_n366), .A3(new_n367), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT34), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n369), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n369), .A2(new_n378), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n366), .A2(new_n367), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  OR3_X1    g180(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT36), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(G155gat), .A2(G162gat), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT2), .ZN(new_n387));
  INV_X1    g186(.A(G148gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n239), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(G141gat), .A2(G148gat), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n387), .A2(new_n389), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G155gat), .B(G162gat), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT82), .B1(G155gat), .B2(G162gat), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n392), .B1(new_n391), .B2(new_n393), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n396));
  NOR3_X1   g195(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G141gat), .B(G148gat), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT2), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n399), .B1(G155gat), .B2(G162gat), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n393), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n392), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT3), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n397), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n385), .B1(new_n290), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n354), .A2(new_n356), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n395), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AND4_X1   g210(.A1(new_n408), .A2(new_n409), .A3(new_n270), .A4(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n408), .B1(new_n357), .B2(new_n411), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n407), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n290), .A2(new_n410), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n357), .A2(new_n411), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n417), .A2(KEYINPUT84), .A3(new_n418), .ZN(new_n419));
  OR3_X1    g218(.A1(new_n357), .A2(KEYINPUT84), .A3(new_n411), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n385), .A3(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n407), .B(KEYINPUT83), .C1(new_n412), .C2(new_n413), .ZN(new_n422));
  NAND4_X1  g221(.A1(new_n416), .A2(KEYINPUT5), .A3(new_n421), .A4(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n357), .A2(new_n408), .A3(new_n411), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n424), .A2(KEYINPUT85), .ZN(new_n425));
  INV_X1    g224(.A(new_n413), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT85), .ZN(new_n427));
  NAND4_X1  g226(.A1(new_n357), .A2(new_n427), .A3(new_n408), .A4(new_n411), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n425), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n429), .A2(new_n430), .A3(new_n407), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n423), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(G1gat), .B(G29gat), .ZN(new_n433));
  XNOR2_X1  g232(.A(new_n433), .B(KEYINPUT0), .ZN(new_n434));
  XNOR2_X1  g233(.A(G57gat), .B(G85gat), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n434), .B(new_n435), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n432), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n436), .A3(new_n431), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n432), .A2(KEYINPUT6), .A3(new_n437), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT86), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n436), .B1(new_n423), .B2(new_n431), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(KEYINPUT6), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n443), .A3(new_n446), .ZN(new_n447));
  XNOR2_X1  g246(.A(G8gat), .B(G36gat), .ZN(new_n448));
  XNOR2_X1  g247(.A(G64gat), .B(G92gat), .ZN(new_n449));
  XOR2_X1   g248(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND2_X1  g249(.A1(G226gat), .A2(G233gat), .ZN(new_n451));
  XOR2_X1   g250(.A(new_n451), .B(KEYINPUT81), .Z(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n343), .B2(KEYINPUT29), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n455));
  XNOR2_X1  g254(.A(G211gat), .B(G218gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT79), .ZN(new_n457));
  XNOR2_X1  g256(.A(G197gat), .B(G204gat), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT22), .ZN(new_n459));
  INV_X1    g258(.A(G211gat), .ZN(new_n460));
  INV_X1    g259(.A(G218gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT79), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n456), .B(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n463), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n455), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n466), .A2(new_n467), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n457), .A2(new_n463), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT80), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n353), .A2(new_n452), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n454), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n473), .B1(new_n454), .B2(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n450), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n469), .A2(new_n472), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT29), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n452), .B1(new_n353), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n343), .A2(new_n453), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n479), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n450), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n475), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n478), .A2(KEYINPUT30), .A3(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT30), .ZN(new_n487));
  OAI211_X1 g286(.A(new_n487), .B(new_n450), .C1(new_n476), .C2(new_n477), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n486), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n447), .A2(new_n489), .ZN(new_n490));
  XNOR2_X1  g289(.A(G78gat), .B(G106gat), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n405), .A2(KEYINPUT29), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n479), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n470), .A2(new_n471), .A3(new_n480), .ZN(new_n494));
  AND2_X1   g293(.A1(new_n494), .A2(new_n396), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(new_n411), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n491), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n491), .ZN(new_n498));
  OAI221_X1 g297(.A(new_n498), .B1(new_n495), .B2(new_n411), .C1(new_n479), .C2(new_n492), .ZN(new_n499));
  NAND2_X1  g298(.A1(G228gat), .A2(G233gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(G22gat), .ZN(new_n501));
  XOR2_X1   g300(.A(KEYINPUT31), .B(G50gat), .Z(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n497), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n497), .B2(new_n499), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n383), .B1(new_n490), .B2(new_n507), .ZN(new_n508));
  AND4_X1   g307(.A1(new_n445), .A2(new_n432), .A3(KEYINPUT6), .A4(new_n437), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n445), .B1(new_n444), .B2(KEYINPUT6), .ZN(new_n510));
  NOR2_X1   g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n432), .A2(KEYINPUT88), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT88), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n423), .A2(new_n513), .A3(new_n431), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n512), .A2(new_n437), .A3(new_n514), .ZN(new_n515));
  AND2_X1   g314(.A1(new_n440), .A2(new_n439), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n478), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT37), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n483), .A2(new_n475), .A3(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n483), .B2(new_n475), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n484), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n518), .B1(new_n522), .B2(KEYINPUT38), .ZN(new_n523));
  INV_X1    g322(.A(new_n521), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n483), .A2(new_n475), .A3(new_n519), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT89), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT38), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n526), .A2(new_n527), .A3(new_n528), .A4(new_n484), .ZN(new_n529));
  OAI211_X1 g328(.A(new_n528), .B(new_n484), .C1(new_n520), .C2(new_n521), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(KEYINPUT89), .ZN(new_n531));
  AND3_X1   g330(.A1(new_n523), .A2(new_n529), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n517), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n290), .A2(new_n406), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n384), .B1(new_n429), .B2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT39), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(new_n436), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n385), .B1(new_n419), .B2(new_n420), .ZN(new_n539));
  NOR3_X1   g338(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n489), .B1(new_n541), .B2(KEYINPUT40), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT40), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n543), .B1(new_n538), .B2(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT87), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n546), .B(new_n543), .C1(new_n538), .C2(new_n540), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n542), .A2(new_n545), .A3(new_n515), .A4(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n533), .A2(new_n548), .A3(new_n506), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n508), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n375), .A2(new_n507), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n447), .A2(new_n489), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT35), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n511), .A2(new_n517), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n377), .B2(new_n381), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n368), .A2(new_n371), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n370), .A2(new_n366), .A3(new_n367), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT90), .A3(new_n558), .ZN(new_n559));
  AND4_X1   g358(.A1(new_n489), .A2(new_n556), .A3(new_n506), .A4(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT35), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n554), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n553), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n550), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT91), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n550), .A2(KEYINPUT91), .A3(new_n563), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n248), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  XOR2_X1   g367(.A(G57gat), .B(G64gat), .Z(new_n569));
  INV_X1    g368(.A(KEYINPUT9), .ZN(new_n570));
  INV_X1    g369(.A(G71gat), .ZN(new_n571));
  INV_X1    g370(.A(G78gat), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  AOI22_X1  g373(.A1(new_n569), .A2(new_n573), .B1(new_n574), .B2(KEYINPUT98), .ZN(new_n575));
  INV_X1    g374(.A(new_n574), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT98), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n576), .A2(new_n569), .A3(new_n577), .A4(new_n573), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g380(.A1(new_n581), .A2(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  NOR2_X1   g383(.A1(new_n584), .A2(new_n259), .ZN(new_n585));
  INV_X1    g384(.A(new_n583), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n582), .B(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n587), .A2(G127gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT100), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n581), .B(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n220), .B1(new_n590), .B2(KEYINPUT21), .ZN(new_n591));
  OR3_X1    g390(.A1(new_n585), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n591), .B1(new_n585), .B2(new_n588), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT99), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(G155gat), .ZN(new_n596));
  XOR2_X1   g395(.A(G183gat), .B(G211gat), .Z(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  AND3_X1   g397(.A1(new_n592), .A2(new_n593), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n592), .B2(new_n593), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G85gat), .A2(G92gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(KEYINPUT7), .ZN(new_n603));
  NAND2_X1  g402(.A1(G99gat), .A2(G106gat), .ZN(new_n604));
  INV_X1    g403(.A(G85gat), .ZN(new_n605));
  INV_X1    g404(.A(G92gat), .ZN(new_n606));
  AOI22_X1  g405(.A1(KEYINPUT8), .A2(new_n604), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n214), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n610), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n214), .B2(new_n222), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n611), .B(new_n612), .C1(new_n614), .C2(new_n225), .ZN(new_n615));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n616), .B(KEYINPUT101), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n615), .B1(KEYINPUT102), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(KEYINPUT102), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n619), .B(new_n620), .Z(new_n621));
  AND2_X1   g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n618), .A2(new_n621), .ZN(new_n623));
  XNOR2_X1  g422(.A(G134gat), .B(G162gat), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT103), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n622), .B2(new_n623), .ZN(new_n628));
  INV_X1    g427(.A(G230gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n629), .A2(new_n360), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n581), .B1(KEYINPUT104), .B2(new_n609), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n631), .A2(new_n613), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n631), .A2(new_n613), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n590), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n634), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n639), .A2(new_n630), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(G176gat), .B(G204gat), .ZN(new_n642));
  XOR2_X1   g441(.A(new_n641), .B(new_n642), .Z(new_n643));
  NAND3_X1  g442(.A1(new_n638), .A2(new_n640), .A3(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n643), .B1(new_n638), .B2(new_n640), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g446(.A1(new_n601), .A2(new_n627), .A3(new_n628), .A4(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n568), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n447), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(G1gat), .Z(G1324gat));
  OAI21_X1  g451(.A(G8gat), .B1(new_n650), .B2(new_n489), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n653), .B(KEYINPUT106), .Z(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(new_n489), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT42), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT16), .B(G8gat), .Z(new_n657));
  AND4_X1   g456(.A1(KEYINPUT105), .A2(new_n655), .A3(new_n656), .A4(new_n657), .ZN(new_n658));
  OR3_X1    g457(.A1(new_n650), .A2(KEYINPUT105), .A3(new_n489), .ZN(new_n659));
  AOI22_X1  g458(.A1(new_n659), .A2(new_n656), .B1(new_n655), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n654), .B1(new_n658), .B2(new_n660), .ZN(G1325gat));
  INV_X1    g460(.A(new_n383), .ZN(new_n662));
  OAI21_X1  g461(.A(G15gat), .B1(new_n650), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n556), .A2(new_n559), .ZN(new_n664));
  OR2_X1    g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n663), .B1(new_n650), .B2(new_n665), .ZN(G1326gat));
  NOR2_X1   g465(.A1(new_n650), .A2(new_n506), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT43), .B(G22gat), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  INV_X1    g468(.A(new_n447), .ZN(new_n670));
  INV_X1    g469(.A(new_n647), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n601), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n627), .A2(new_n628), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n568), .A2(new_n670), .A3(new_n204), .A4(new_n676), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT45), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n566), .A2(new_n567), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n674), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT44), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n564), .A2(KEYINPUT107), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT107), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n550), .B2(new_n563), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n674), .A2(new_n685), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n682), .A2(new_n684), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n681), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n244), .A2(new_n245), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n673), .A2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n690), .A2(new_n447), .A3(new_n694), .ZN(new_n695));
  OAI21_X1  g494(.A(new_n678), .B1(new_n695), .B2(new_n204), .ZN(G1328gat));
  INV_X1    g495(.A(new_n489), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n568), .A2(new_n697), .A3(new_n203), .A4(new_n676), .ZN(new_n698));
  XOR2_X1   g497(.A(new_n698), .B(KEYINPUT46), .Z(new_n699));
  NOR3_X1   g498(.A1(new_n690), .A2(new_n489), .A3(new_n694), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n203), .ZN(G1329gat));
  NAND2_X1  g500(.A1(new_n568), .A2(new_n676), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(G43gat), .A3(new_n664), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n689), .A2(new_n383), .A3(new_n693), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n704), .B2(G43gat), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT47), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT47), .B(new_n703), .C1(new_n704), .C2(G43gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n707), .A2(new_n708), .ZN(G1330gat));
  INV_X1    g508(.A(KEYINPUT108), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n506), .B(new_n694), .C1(new_n681), .C2(new_n688), .ZN(new_n711));
  INV_X1    g510(.A(G50gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND4_X1  g512(.A1(new_n568), .A2(new_n712), .A3(new_n507), .A4(new_n676), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n714), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT48), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n713), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  OAI221_X1 g516(.A(new_n714), .B1(new_n710), .B2(KEYINPUT48), .C1(new_n711), .C2(new_n712), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1331gat));
  NAND4_X1  g518(.A1(new_n675), .A2(new_n692), .A3(new_n601), .A4(new_n671), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n682), .A2(new_n684), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n721), .A2(new_n670), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n697), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT49), .B(G64gat), .Z(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT109), .ZN(G1333gat));
  AOI21_X1  g527(.A(new_n571), .B1(new_n721), .B2(new_n383), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n664), .A2(G71gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n721), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g531(.A1(new_n721), .A2(new_n507), .ZN(new_n733));
  XNOR2_X1  g532(.A(KEYINPUT110), .B(G78gat), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n733), .B(new_n734), .ZN(G1335gat));
  INV_X1    g534(.A(new_n601), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(new_n692), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n647), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n689), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(G85gat), .B1(new_n739), .B2(new_n447), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n675), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n564), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(KEYINPUT51), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT51), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n564), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n671), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n670), .A2(new_n605), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n740), .B1(new_n747), .B2(new_n748), .ZN(G1336gat));
  INV_X1    g548(.A(KEYINPUT52), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n689), .A2(new_n697), .A3(new_n738), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n744), .A2(KEYINPUT111), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n742), .B(new_n752), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n489), .A2(G92gat), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n647), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n751), .A2(G92gat), .B1(new_n753), .B2(new_n756), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n751), .A2(G92gat), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT112), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n747), .B2(new_n755), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n746), .A2(KEYINPUT112), .A3(new_n671), .A4(new_n754), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n760), .A2(new_n750), .A3(new_n761), .ZN(new_n762));
  OAI22_X1  g561(.A1(new_n750), .A2(new_n757), .B1(new_n758), .B2(new_n762), .ZN(G1337gat));
  OAI21_X1  g562(.A(G99gat), .B1(new_n739), .B2(new_n662), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n664), .A2(G99gat), .A3(new_n647), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT113), .Z(new_n766));
  NAND2_X1  g565(.A1(new_n746), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(G1338gat));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n506), .A2(G106gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n743), .A2(new_n671), .A3(new_n745), .A4(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT116), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(new_n772), .B2(new_n771), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n685), .B1(new_n679), .B2(new_n674), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n507), .B(new_n738), .C1(new_n775), .C2(new_n687), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(G106gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n776), .A2(KEYINPUT114), .A3(G106gat), .ZN(new_n779));
  AOI21_X1  g578(.A(KEYINPUT114), .B1(new_n776), .B2(G106gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n647), .A2(G106gat), .A3(new_n506), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n753), .A2(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(KEYINPUT115), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n753), .A2(KEYINPUT115), .A3(new_n781), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n779), .A2(new_n780), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n778), .B1(new_n787), .B2(new_n769), .ZN(G1339gat));
  NOR2_X1   g587(.A1(new_n648), .A2(new_n691), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT117), .ZN(new_n790));
  XNOR2_X1  g589(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n635), .A2(new_n630), .A3(new_n636), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n638), .A2(KEYINPUT54), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT54), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n643), .B1(new_n637), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT55), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n793), .A2(KEYINPUT55), .A3(new_n795), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n644), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT118), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n798), .A2(KEYINPUT118), .A3(new_n644), .A4(new_n799), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n691), .A3(new_n803), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n223), .A2(new_n225), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n202), .B1(new_n805), .B2(new_n221), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n230), .A2(new_n231), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n241), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g607(.A1(new_n245), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n671), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n674), .B1(new_n804), .B2(new_n810), .ZN(new_n811));
  AND4_X1   g610(.A1(new_n674), .A2(new_n802), .A3(new_n803), .A4(new_n809), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n736), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n447), .B1(new_n791), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n560), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT97), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n691), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n244), .A2(KEYINPUT97), .A3(new_n245), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n236), .B1(new_n815), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g619(.A(new_n820), .B(KEYINPUT119), .Z(new_n821));
  AND3_X1   g620(.A1(new_n814), .A2(new_n489), .A3(new_n551), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n822), .A2(new_n236), .A3(new_n691), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(G1340gat));
  AOI21_X1  g623(.A(G120gat), .B1(new_n822), .B2(new_n671), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n647), .A2(new_n263), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n815), .B2(new_n826), .ZN(G1341gat));
  INV_X1    g626(.A(new_n815), .ZN(new_n828));
  OAI21_X1  g627(.A(G127gat), .B1(new_n828), .B2(new_n736), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n822), .A2(new_n259), .A3(new_n601), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(G1342gat));
  NOR2_X1   g630(.A1(new_n675), .A2(new_n697), .ZN(new_n832));
  NAND4_X1  g631(.A1(new_n814), .A2(new_n254), .A3(new_n551), .A4(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n828), .B2(new_n675), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1343gat));
  AOI211_X1 g635(.A(new_n506), .B(new_n383), .C1(new_n814), .C2(KEYINPUT121), .ZN(new_n837));
  OR2_X1    g636(.A1(new_n814), .A2(KEYINPUT121), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n837), .A2(new_n489), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n248), .A2(G141gat), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT58), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n383), .A2(new_n447), .A3(new_n697), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n506), .B1(new_n791), .B2(new_n813), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT57), .ZN(new_n848));
  AND3_X1   g647(.A1(new_n798), .A2(new_n644), .A3(new_n799), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n849), .B1(new_n246), .B2(new_n247), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n674), .B1(new_n850), .B2(new_n810), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n736), .B1(new_n851), .B2(new_n812), .ZN(new_n852));
  AOI211_X1 g651(.A(new_n848), .B(new_n506), .C1(new_n791), .C2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n843), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  OAI21_X1  g653(.A(G141gat), .B1(new_n854), .B2(new_n248), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n841), .A2(new_n842), .A3(new_n855), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n691), .B(new_n843), .C1(new_n847), .C2(new_n853), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n839), .A2(new_n840), .B1(new_n857), .B2(G141gat), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n842), .B2(new_n858), .ZN(G1344gat));
  NOR2_X1   g658(.A1(new_n388), .A2(KEYINPUT59), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n854), .B2(new_n647), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n506), .B(new_n845), .C1(new_n791), .C2(new_n813), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n674), .A2(new_n809), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n800), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n736), .B1(new_n851), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT123), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n819), .B2(new_n648), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n649), .A2(KEYINPUT123), .A3(new_n248), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT57), .B1(new_n869), .B2(new_n507), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n871), .A2(new_n647), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n388), .B1(new_n872), .B2(new_n843), .ZN(new_n873));
  XOR2_X1   g672(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n874));
  OAI21_X1  g673(.A(new_n861), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n839), .A2(new_n388), .A3(new_n671), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(G1345gat));
  OAI21_X1  g676(.A(G155gat), .B1(new_n854), .B2(new_n736), .ZN(new_n878));
  INV_X1    g677(.A(new_n839), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n736), .A2(G155gat), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n878), .B1(new_n879), .B2(new_n880), .ZN(G1346gat));
  OAI21_X1  g680(.A(G162gat), .B1(new_n854), .B2(new_n675), .ZN(new_n882));
  INV_X1    g681(.A(G162gat), .ZN(new_n883));
  NAND4_X1  g682(.A1(new_n837), .A2(new_n883), .A3(new_n832), .A4(new_n838), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(new_n884), .ZN(G1347gat));
  NAND2_X1  g684(.A1(new_n791), .A2(new_n813), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n670), .A2(new_n489), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n664), .A2(new_n507), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n890), .A2(new_n305), .A3(new_n248), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n886), .A2(new_n551), .A3(new_n887), .ZN(new_n892));
  AOI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n691), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n891), .A2(new_n893), .ZN(G1348gat));
  OAI21_X1  g693(.A(G176gat), .B1(new_n890), .B2(new_n647), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n892), .A2(new_n306), .A3(new_n671), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(KEYINPUT124), .ZN(G1349gat));
  OAI21_X1  g697(.A(new_n295), .B1(new_n890), .B2(new_n736), .ZN(new_n899));
  OAI211_X1 g698(.A(new_n892), .B(new_n601), .C1(new_n318), .C2(new_n319), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901));
  AOI22_X1  g700(.A1(new_n899), .A2(new_n900), .B1(KEYINPUT125), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(KEYINPUT125), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n902), .B(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n892), .A2(new_n312), .A3(new_n674), .ZN(new_n905));
  OAI21_X1  g704(.A(G190gat), .B1(new_n890), .B2(new_n675), .ZN(new_n906));
  AND2_X1   g705(.A1(new_n906), .A2(KEYINPUT61), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n906), .A2(KEYINPUT61), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n905), .B1(new_n907), .B2(new_n908), .ZN(G1351gat));
  NAND2_X1  g708(.A1(new_n887), .A2(new_n662), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n819), .B(new_n911), .C1(new_n862), .C2(new_n870), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(KEYINPUT126), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n868), .A2(new_n867), .ZN(new_n914));
  AOI22_X1  g713(.A1(new_n819), .A2(new_n849), .B1(new_n671), .B2(new_n809), .ZN(new_n915));
  OAI22_X1  g714(.A1(new_n915), .A2(new_n674), .B1(new_n800), .B2(new_n863), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n914), .B1(new_n916), .B2(new_n736), .ZN(new_n917));
  OAI21_X1  g716(.A(new_n848), .B1(new_n917), .B2(new_n506), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n844), .A2(new_n846), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n819), .A4(new_n911), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n913), .A2(G197gat), .A3(new_n922), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n844), .A2(new_n911), .ZN(new_n924));
  INV_X1    g723(.A(G197gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n691), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT127), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n923), .A2(KEYINPUT127), .A3(new_n926), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1352gat));
  INV_X1    g730(.A(G204gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n924), .A2(new_n932), .A3(new_n671), .ZN(new_n933));
  XNOR2_X1  g732(.A(new_n933), .B(KEYINPUT62), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n872), .B2(new_n911), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n934), .A2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n460), .A3(new_n601), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n871), .A2(new_n910), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(new_n601), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  NAND3_X1  g741(.A1(new_n924), .A2(new_n461), .A3(new_n674), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n871), .A2(new_n675), .A3(new_n910), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n944), .B2(new_n461), .ZN(G1355gat));
endmodule


