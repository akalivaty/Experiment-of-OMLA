//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:11 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n674, new_n675, new_n676, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n776, new_n777, new_n778,
    new_n779, new_n781, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n858, new_n859, new_n860, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  NAND2_X1  g002(.A1(G228gat), .A2(G233gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n204), .B(KEYINPUT77), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT72), .ZN(new_n207));
  XNOR2_X1  g006(.A(G141gat), .B(G148gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(G155gat), .B2(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n207), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(G155gat), .B(G162gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT2), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  INV_X1    g016(.A(G148gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G141gat), .A2(G148gat), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(new_n219), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n221), .A2(new_n207), .A3(new_n212), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n214), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT3), .ZN(new_n224));
  NAND2_X1  g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G197gat), .A2(G204gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(G197gat), .A2(G204gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(new_n225), .ZN(new_n232));
  NOR2_X1   g031(.A1(G211gat), .A2(G218gat), .ZN(new_n233));
  NOR3_X1   g032(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT69), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT69), .ZN(new_n235));
  INV_X1    g034(.A(G211gat), .ZN(new_n236));
  INV_X1    g035(.A(G218gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n235), .B1(new_n238), .B2(new_n225), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n231), .B1(new_n234), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT29), .ZN(new_n241));
  OR2_X1    g040(.A1(G197gat), .A2(G204gat), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n242), .A2(new_n228), .B1(new_n226), .B2(new_n225), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT69), .B1(new_n232), .B2(new_n233), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n238), .A2(new_n235), .A3(new_n225), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n223), .B1(new_n224), .B2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n240), .A2(new_n246), .ZN(new_n249));
  AOI21_X1  g048(.A(KEYINPUT3), .B1(new_n214), .B2(new_n222), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n249), .B1(new_n250), .B2(KEYINPUT29), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n248), .B1(new_n251), .B2(KEYINPUT78), .ZN(new_n252));
  AND3_X1   g051(.A1(new_n243), .A2(new_n244), .A3(new_n245), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n242), .A2(new_n228), .ZN(new_n254));
  AOI22_X1  g053(.A1(new_n244), .A2(new_n245), .B1(new_n254), .B2(new_n227), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n221), .A2(new_n207), .A3(new_n212), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n212), .B1(new_n221), .B2(new_n207), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n224), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n256), .B1(new_n259), .B2(new_n241), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT78), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n206), .B1(new_n252), .B2(new_n262), .ZN(new_n263));
  NOR3_X1   g062(.A1(new_n260), .A2(new_n248), .A3(new_n204), .ZN(new_n264));
  OAI21_X1  g063(.A(G22gat), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n224), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n257), .A2(new_n258), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n268), .B1(new_n260), .B2(new_n261), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n251), .A2(KEYINPUT78), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n205), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n264), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G78gat), .B(G106gat), .ZN(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n265), .A2(new_n274), .A3(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n276), .B1(new_n265), .B2(new_n274), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n203), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n263), .A2(G22gat), .A3(new_n264), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n272), .B1(new_n271), .B2(new_n273), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n275), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n274), .A3(new_n276), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(new_n202), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(new_n279), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G1gat), .B(G29gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n286), .B(KEYINPUT0), .ZN(new_n287));
  XNOR2_X1  g086(.A(G57gat), .B(G85gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n287), .B(new_n288), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  XOR2_X1   g091(.A(G127gat), .B(G134gat), .Z(new_n293));
  XNOR2_X1  g092(.A(G113gat), .B(G120gat), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n293), .B1(KEYINPUT1), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g094(.A(G113gat), .B(G120gat), .Z(new_n296));
  INV_X1    g095(.A(KEYINPUT1), .ZN(new_n297));
  XNOR2_X1  g096(.A(G127gat), .B(G134gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT73), .B1(new_n267), .B2(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n295), .A2(new_n299), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT73), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n223), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n301), .B(new_n304), .C1(new_n223), .C2(new_n302), .ZN(new_n305));
  NAND2_X1  g104(.A1(G225gat), .A2(G233gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT4), .ZN(new_n310));
  NOR3_X1   g109(.A1(new_n267), .A2(KEYINPUT73), .A3(new_n300), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n303), .B1(new_n223), .B2(new_n302), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT74), .ZN(new_n314));
  AOI21_X1  g113(.A(KEYINPUT4), .B1(new_n301), .B2(new_n304), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT4), .B1(new_n267), .B2(new_n300), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n214), .A2(KEYINPUT3), .A3(new_n222), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n259), .A2(new_n320), .A3(new_n300), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(new_n306), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n309), .B1(new_n319), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n301), .A2(KEYINPUT4), .A3(new_n304), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n267), .A2(new_n300), .ZN(new_n326));
  AOI21_X1  g125(.A(KEYINPUT75), .B1(new_n326), .B2(new_n310), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n322), .A2(KEYINPUT5), .ZN(new_n329));
  NAND4_X1  g128(.A1(new_n301), .A2(KEYINPUT75), .A3(new_n304), .A4(KEYINPUT4), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n290), .B(new_n292), .C1(new_n324), .C2(new_n331), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n318), .B1(new_n315), .B2(new_n316), .ZN(new_n333));
  AOI211_X1 g132(.A(KEYINPUT74), .B(KEYINPUT4), .C1(new_n301), .C2(new_n304), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n323), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n331), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n291), .B1(new_n337), .B2(new_n289), .ZN(new_n338));
  NOR3_X1   g137(.A1(new_n324), .A2(new_n290), .A3(new_n331), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT71), .ZN(new_n342));
  INV_X1    g141(.A(G183gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n343), .A2(KEYINPUT27), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT27), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G183gat), .ZN(new_n346));
  INV_X1    g145(.A(G190gat), .ZN(new_n347));
  NOR2_X1   g146(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n348));
  NAND4_X1  g147(.A1(new_n344), .A2(new_n346), .A3(new_n347), .A4(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT26), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT26), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n359));
  AND2_X1   g158(.A1(KEYINPUT66), .A2(KEYINPUT28), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n360), .A2(new_n348), .ZN(new_n361));
  AOI22_X1  g160(.A1(new_n357), .A2(new_n358), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT25), .ZN(new_n363));
  OAI211_X1 g162(.A(new_n363), .B(new_n358), .C1(new_n353), .C2(KEYINPUT23), .ZN(new_n364));
  INV_X1    g163(.A(G176gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT64), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT64), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(G176gat), .ZN(new_n368));
  AND2_X1   g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(G169gat), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n370), .A2(KEYINPUT23), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n364), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n350), .A2(KEYINPUT24), .ZN(new_n373));
  XOR2_X1   g172(.A(G183gat), .B(G190gat), .Z(new_n374));
  AOI21_X1  g173(.A(new_n373), .B1(new_n374), .B2(KEYINPUT24), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n352), .A2(new_n362), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n370), .A2(new_n365), .A3(KEYINPUT23), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n358), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(KEYINPUT65), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT23), .B1(new_n370), .B2(new_n365), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n347), .A2(G183gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n343), .A2(G190gat), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT24), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT65), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n377), .A2(new_n386), .A3(new_n358), .ZN(new_n387));
  INV_X1    g186(.A(new_n373), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT25), .B1(new_n382), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n376), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(G226gat), .A2(G233gat), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n256), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n385), .A2(new_n387), .A3(new_n388), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n380), .B1(new_n378), .B2(KEYINPUT65), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n363), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n358), .A2(new_n363), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n380), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n371), .A2(new_n366), .A3(new_n368), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n385), .A2(new_n400), .A3(new_n401), .A4(new_n388), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n359), .A2(new_n361), .ZN(new_n403));
  NOR3_X1   g202(.A1(new_n355), .A2(G169gat), .A3(G176gat), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT26), .B1(new_n370), .B2(new_n365), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n358), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n402), .B1(new_n407), .B2(new_n351), .ZN(new_n408));
  NOR3_X1   g207(.A1(new_n398), .A2(new_n408), .A3(KEYINPUT70), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT70), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n410), .B1(new_n376), .B2(new_n390), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n241), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n395), .B1(new_n412), .B2(new_n392), .ZN(new_n413));
  OAI21_X1  g212(.A(KEYINPUT70), .B1(new_n398), .B2(new_n408), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n376), .A2(new_n390), .A3(new_n410), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(new_n415), .A3(new_n393), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n241), .A3(new_n392), .ZN(new_n417));
  AND3_X1   g216(.A1(new_n416), .A2(new_n249), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n342), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n249), .B1(new_n391), .B2(new_n393), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT29), .B1(new_n414), .B2(new_n415), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n420), .B1(new_n421), .B2(new_n393), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n416), .A2(new_n249), .A3(new_n417), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n422), .A2(KEYINPUT71), .A3(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G8gat), .B(G36gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(G64gat), .B(G92gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n419), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n415), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n393), .B1(new_n430), .B2(new_n241), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n423), .B(new_n427), .C1(new_n431), .C2(new_n395), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n422), .A2(KEYINPUT30), .A3(new_n423), .A4(new_n427), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n285), .B1(new_n341), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT36), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n439));
  XOR2_X1   g238(.A(G71gat), .B(G99gat), .Z(new_n440));
  XNOR2_X1  g239(.A(G15gat), .B(G43gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  AND2_X1   g241(.A1(G227gat), .A2(G233gat), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n300), .B1(new_n398), .B2(new_n408), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n376), .A2(new_n390), .A3(new_n302), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n439), .B(new_n442), .C1(new_n447), .C2(KEYINPUT33), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT32), .ZN(new_n449));
  OR2_X1    g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n448), .A2(new_n450), .ZN(new_n451));
  OAI211_X1 g250(.A(KEYINPUT67), .B(new_n442), .C1(new_n447), .C2(KEYINPUT33), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n442), .A2(KEYINPUT33), .ZN(new_n453));
  NOR3_X1   g252(.A1(new_n447), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n445), .A2(new_n446), .A3(new_n444), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT68), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT34), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT34), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n460), .A2(new_n462), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n451), .B2(new_n455), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n438), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n456), .A2(new_n463), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n465), .A2(new_n451), .A3(new_n455), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n468), .A2(KEYINPUT36), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n279), .A2(new_n284), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n332), .A2(KEYINPUT81), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n335), .A2(new_n336), .ZN(new_n474));
  INV_X1    g273(.A(new_n331), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT81), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n290), .A4(new_n292), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n473), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n290), .B1(new_n324), .B2(new_n331), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n474), .A2(new_n289), .A3(new_n475), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n480), .A2(new_n481), .A3(new_n291), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT38), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n419), .A2(KEYINPUT37), .A3(new_n424), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT37), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n422), .A2(new_n486), .A3(new_n423), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n487), .A2(new_n428), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n484), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n394), .A2(new_n249), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n431), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n416), .A2(new_n256), .A3(new_n417), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT37), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n484), .B1(new_n491), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n487), .A2(new_n428), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n432), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n472), .B1(new_n483), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT40), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n328), .A2(new_n321), .A3(new_n330), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(new_n307), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n305), .A2(new_n307), .ZN(new_n502));
  AND3_X1   g301(.A1(new_n501), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT39), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n500), .A2(new_n504), .A3(new_n307), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n289), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n499), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT79), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT79), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n509), .B(new_n499), .C1(new_n503), .C2(new_n506), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n501), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(KEYINPUT40), .A3(new_n289), .A4(new_n505), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT80), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n508), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  OAI211_X1 g314(.A(new_n436), .B(new_n480), .C1(new_n512), .C2(new_n513), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g316(.A(new_n437), .B(new_n471), .C1(new_n498), .C2(new_n517), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n422), .A2(KEYINPUT71), .A3(new_n423), .ZN(new_n519));
  AOI21_X1  g318(.A(KEYINPUT71), .B1(new_n422), .B2(new_n423), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n519), .A2(new_n520), .A3(new_n427), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n434), .A2(new_n435), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n464), .A2(new_n466), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n472), .A2(new_n340), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n468), .A2(KEYINPUT82), .A3(new_n469), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT82), .B1(new_n468), .B2(new_n469), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT35), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n429), .A2(new_n530), .A3(new_n434), .A4(new_n435), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n531), .B1(new_n284), .B2(new_n279), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n483), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(G232gat), .A2(G233gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT41), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(G29gat), .A2(G36gat), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT14), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G29gat), .ZN(new_n542));
  INV_X1    g341(.A(G36gat), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G43gat), .B(G50gat), .ZN(new_n545));
  AND2_X1   g344(.A1(new_n545), .A2(KEYINPUT15), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT83), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n546), .B(KEYINPUT84), .ZN(new_n550));
  OAI22_X1  g349(.A1(new_n545), .A2(KEYINPUT15), .B1(new_n542), .B2(new_n543), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT85), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(new_n541), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n550), .B(new_n553), .C1(new_n552), .C2(new_n541), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n549), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT17), .ZN(new_n556));
  XOR2_X1   g355(.A(KEYINPUT90), .B(G85gat), .Z(new_n557));
  INV_X1    g356(.A(G92gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G85gat), .ZN(new_n560));
  OAI21_X1  g359(.A(KEYINPUT89), .B1(new_n560), .B2(new_n558), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT89), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n562), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n561), .A2(new_n563), .A3(KEYINPUT7), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT7), .ZN(new_n565));
  OAI211_X1 g364(.A(KEYINPUT89), .B(new_n565), .C1(new_n560), .C2(new_n558), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n567), .A2(KEYINPUT8), .ZN(new_n568));
  NAND4_X1  g367(.A1(new_n559), .A2(new_n564), .A3(new_n566), .A4(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT91), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n538), .B1(new_n556), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n555), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(new_n573), .ZN(new_n576));
  XOR2_X1   g375(.A(G190gat), .B(G218gat), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n536), .A2(new_n537), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT88), .Z(new_n580));
  XNOR2_X1  g379(.A(G134gat), .B(G162gat), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n580), .B(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(new_n578), .B(new_n582), .Z(new_n583));
  XOR2_X1   g382(.A(G57gat), .B(G64gat), .Z(new_n584));
  AND2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n584), .B1(KEYINPUT9), .B2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G71gat), .B(G78gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT21), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(G231gat), .A2(G233gat), .ZN(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G127gat), .B(G155gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(KEYINPUT20), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n592), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(G183gat), .B(G211gat), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(G15gat), .B(G22gat), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT16), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(G1gat), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n600), .B1(G1gat), .B2(new_n598), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G8gat), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n603), .B1(new_n589), .B2(new_n588), .ZN(new_n604));
  XOR2_X1   g403(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XOR2_X1   g405(.A(new_n597), .B(new_n606), .Z(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n583), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G120gat), .B(G148gat), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT94), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XOR2_X1   g411(.A(new_n611), .B(new_n612), .Z(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  OR2_X1    g413(.A1(new_n569), .A2(new_n570), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT92), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n588), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n571), .ZN(new_n618));
  NAND2_X1  g417(.A1(G230gat), .A2(G233gat), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT93), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n588), .A2(new_n625), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n626), .B1(new_n573), .B2(new_n627), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n619), .B(KEYINPUT95), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n614), .B1(new_n624), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n628), .A2(new_n619), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n622), .A2(new_n634), .A3(new_n623), .A4(new_n613), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT18), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n556), .A2(new_n603), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n555), .A2(new_n602), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G229gat), .A2(G233gat), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n638), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n639), .A2(KEYINPUT18), .A3(new_n642), .A4(new_n640), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT86), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n555), .B2(new_n602), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n640), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n642), .B(KEYINPUT13), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n644), .A2(new_n645), .A3(new_n650), .ZN(new_n651));
  XNOR2_X1  g450(.A(G113gat), .B(G141gat), .ZN(new_n652));
  INV_X1    g451(.A(G197gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(KEYINPUT11), .B(G169gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(new_n656), .B(KEYINPUT12), .Z(new_n657));
  NAND2_X1  g456(.A1(new_n651), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n657), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n659), .A3(new_n645), .A4(new_n650), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n535), .A2(new_n609), .A3(new_n637), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(KEYINPUT96), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n340), .ZN(new_n664));
  XOR2_X1   g463(.A(KEYINPUT97), .B(G1gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(G1324gat));
  INV_X1    g465(.A(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n436), .ZN(new_n668));
  AND2_X1   g467(.A1(new_n668), .A2(G8gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(KEYINPUT16), .B(G8gat), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(KEYINPUT42), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n672), .B1(KEYINPUT42), .B2(new_n671), .ZN(G1325gat));
  INV_X1    g472(.A(new_n529), .ZN(new_n674));
  OR3_X1    g473(.A1(new_n663), .A2(G15gat), .A3(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(G15gat), .B1(new_n663), .B2(new_n471), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n663), .A2(new_n472), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT98), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT43), .B(G22gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1327gat));
  NAND3_X1  g480(.A1(new_n608), .A2(new_n637), .A3(new_n661), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n535), .A2(new_n583), .A3(new_n683), .ZN(new_n684));
  NOR3_X1   g483(.A1(new_n684), .A2(G29gat), .A3(new_n340), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT99), .B(KEYINPUT45), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n526), .A2(KEYINPUT100), .A3(new_n533), .ZN(new_n689));
  AOI21_X1  g488(.A(KEYINPUT100), .B1(new_n526), .B2(new_n533), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n518), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n578), .B(new_n582), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n692), .A2(KEYINPUT44), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n436), .B1(new_n482), .B2(new_n332), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n471), .B1(new_n694), .B2(new_n472), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n292), .B1(new_n476), .B2(new_n290), .ZN(new_n696));
  AOI22_X1  g495(.A1(new_n473), .A2(new_n478), .B1(new_n696), .B2(new_n481), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n489), .A2(new_n496), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n285), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n507), .A2(KEYINPUT79), .B1(new_n512), .B2(new_n513), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n436), .A2(new_n480), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n512), .A2(new_n513), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .A4(new_n510), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n695), .B1(new_n699), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n468), .A2(KEYINPUT82), .A3(new_n469), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT82), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n706), .B1(new_n464), .B2(new_n466), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT35), .ZN(new_n708));
  AND4_X1   g507(.A1(new_n472), .A2(new_n705), .A3(new_n707), .A4(new_n708), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n709), .A2(new_n483), .B1(new_n525), .B2(KEYINPUT35), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n583), .B1(new_n704), .B2(new_n710), .ZN(new_n711));
  AOI22_X1  g510(.A1(new_n691), .A2(new_n693), .B1(new_n711), .B2(KEYINPUT44), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n688), .B1(new_n712), .B2(new_n682), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n583), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT100), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n534), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n526), .A2(new_n533), .A3(KEYINPUT100), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n715), .B1(new_n719), .B2(new_n518), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n714), .B1(new_n535), .B2(new_n583), .ZN(new_n721));
  OAI211_X1 g520(.A(KEYINPUT101), .B(new_n683), .C1(new_n720), .C2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n713), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(KEYINPUT102), .B1(new_n723), .B2(new_n340), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(G29gat), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n723), .A2(KEYINPUT102), .A3(new_n340), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n687), .B1(new_n725), .B2(new_n726), .ZN(G1328gat));
  OAI21_X1  g526(.A(G36gat), .B1(new_n723), .B2(new_n523), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n684), .A2(G36gat), .A3(new_n523), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT46), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1329gat));
  INV_X1    g530(.A(new_n712), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n683), .ZN(new_n733));
  OAI21_X1  g532(.A(G43gat), .B1(new_n733), .B2(new_n471), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n684), .A2(G43gat), .A3(new_n674), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n734), .A2(KEYINPUT47), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT103), .B(KEYINPUT47), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n471), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n713), .A2(new_n740), .A3(new_n722), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n735), .B1(new_n742), .B2(KEYINPUT104), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT104), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n744), .A3(G43gat), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT105), .B(new_n739), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT105), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n742), .A2(KEYINPUT104), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n745), .A3(new_n736), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n747), .B1(new_n749), .B2(new_n738), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n737), .B1(new_n746), .B2(new_n750), .ZN(G1330gat));
  NOR2_X1   g550(.A1(new_n472), .A2(G50gat), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT107), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT106), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n753), .B1(new_n684), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n755), .B1(new_n754), .B2(new_n684), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT48), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  OAI21_X1  g557(.A(G50gat), .B1(new_n733), .B2(new_n472), .ZN(new_n759));
  AND3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(KEYINPUT108), .ZN(new_n760));
  AOI21_X1  g559(.A(KEYINPUT108), .B1(new_n758), .B2(new_n759), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n713), .A2(new_n285), .A3(new_n722), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n756), .B1(new_n762), .B2(G50gat), .ZN(new_n763));
  OAI22_X1  g562(.A1(new_n760), .A2(new_n761), .B1(KEYINPUT48), .B2(new_n763), .ZN(G1331gat));
  INV_X1    g563(.A(new_n691), .ZN(new_n765));
  INV_X1    g564(.A(new_n661), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n609), .A2(new_n636), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n768), .A2(new_n341), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(G57gat), .ZN(G1332gat));
  NOR3_X1   g569(.A1(new_n765), .A2(new_n767), .A3(new_n523), .ZN(new_n771));
  NOR2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  AND2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n771), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n771), .B2(new_n772), .ZN(G1333gat));
  NAND3_X1  g574(.A1(new_n768), .A2(G71gat), .A3(new_n740), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n529), .B(KEYINPUT109), .ZN(new_n777));
  NOR3_X1   g576(.A1(new_n765), .A2(new_n767), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n776), .B1(new_n778), .B2(G71gat), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g579(.A1(new_n768), .A2(new_n285), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g581(.A1(new_n661), .A2(new_n607), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n691), .A2(new_n583), .A3(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT51), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(KEYINPUT51), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(KEYINPUT111), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n786), .A2(KEYINPUT111), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n636), .A2(new_n341), .A3(new_n557), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n783), .A2(new_n636), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT110), .Z(new_n792));
  NAND2_X1  g591(.A1(new_n732), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n793), .A2(new_n340), .ZN(new_n794));
  OAI22_X1  g593(.A1(new_n789), .A2(new_n790), .B1(new_n557), .B2(new_n794), .ZN(G1336gat));
  NOR3_X1   g594(.A1(new_n637), .A2(G92gat), .A3(new_n523), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n789), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n732), .A2(new_n436), .A3(new_n792), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(G92gat), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n786), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n803), .A2(new_n796), .B1(G92gat), .B2(new_n799), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n798), .A2(new_n802), .B1(new_n801), .B2(new_n804), .ZN(G1337gat));
  XNOR2_X1  g604(.A(KEYINPUT112), .B(G99gat), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n806), .B1(new_n793), .B2(new_n471), .ZN(new_n807));
  OR3_X1    g606(.A1(new_n637), .A2(new_n674), .A3(new_n806), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n789), .B2(new_n808), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n637), .A2(G106gat), .A3(new_n472), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n785), .B2(new_n786), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n813));
  AND2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(G106gat), .B1(new_n793), .B2(new_n472), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n815), .B1(new_n812), .B2(new_n813), .ZN(new_n816));
  OAI21_X1  g615(.A(KEYINPUT53), .B1(new_n814), .B2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n818), .B(new_n815), .C1(new_n789), .C2(new_n811), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(G1339gat));
  OR2_X1    g619(.A1(new_n648), .A2(new_n649), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n641), .A2(new_n643), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(new_n656), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT114), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT114), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n826), .A3(new_n656), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n825), .A2(new_n636), .A3(new_n660), .A4(new_n827), .ZN(new_n828));
  OR2_X1    g627(.A1(new_n631), .A2(KEYINPUT54), .ZN(new_n829));
  OAI211_X1 g628(.A(new_n626), .B(new_n629), .C1(new_n573), .C2(new_n627), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n634), .A2(KEYINPUT54), .A3(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n829), .A2(new_n831), .A3(new_n614), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT55), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n829), .A2(new_n831), .A3(KEYINPUT55), .A4(new_n614), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n635), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n828), .B1(new_n836), .B2(new_n766), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n692), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n825), .A2(new_n660), .A3(new_n827), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n692), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n836), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n607), .B1(new_n838), .B2(new_n842), .ZN(new_n843));
  NOR4_X1   g642(.A1(new_n583), .A2(new_n608), .A3(new_n636), .A4(new_n661), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n845), .A2(new_n340), .ZN(new_n846));
  AND4_X1   g645(.A1(new_n523), .A2(new_n846), .A3(new_n472), .A4(new_n524), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n661), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n341), .A2(new_n523), .ZN(new_n849));
  OR4_X1    g648(.A1(new_n285), .A2(new_n845), .A3(new_n674), .A4(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(G113gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(new_n766), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n848), .A2(new_n852), .ZN(G1340gat));
  AOI21_X1  g652(.A(G120gat), .B1(new_n847), .B2(new_n636), .ZN(new_n854));
  INV_X1    g653(.A(G120gat), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n850), .A2(new_n855), .A3(new_n637), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n854), .A2(new_n856), .ZN(G1341gat));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n847), .A2(new_n858), .A3(new_n607), .ZN(new_n859));
  OAI21_X1  g658(.A(G127gat), .B1(new_n850), .B2(new_n608), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n859), .A2(new_n860), .ZN(G1342gat));
  INV_X1    g660(.A(G134gat), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n862), .A3(new_n583), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n850), .B2(new_n692), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(KEYINPUT56), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G1343gat));
  NOR3_X1   g666(.A1(new_n740), .A2(new_n436), .A3(new_n472), .ZN(new_n868));
  AND2_X1   g667(.A1(new_n846), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n217), .A3(new_n661), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(new_n844), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n873));
  OR2_X1    g672(.A1(new_n828), .A2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n835), .A2(new_n635), .ZN(new_n875));
  INV_X1    g674(.A(new_n832), .ZN(new_n876));
  XOR2_X1   g675(.A(KEYINPUT116), .B(KEYINPUT55), .Z(new_n877));
  OAI211_X1 g676(.A(new_n875), .B(new_n661), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n828), .A2(new_n873), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n874), .A2(new_n878), .A3(new_n879), .ZN(new_n880));
  AOI22_X1  g679(.A1(new_n880), .A2(new_n692), .B1(new_n841), .B2(new_n840), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n872), .B1(new_n881), .B2(new_n607), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n871), .B1(new_n882), .B2(new_n285), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n692), .A2(new_n837), .B1(new_n840), .B2(new_n841), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n872), .B1(new_n884), .B2(new_n607), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n285), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n849), .A2(new_n740), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NOR4_X1   g688(.A1(new_n883), .A2(new_n887), .A3(new_n766), .A4(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n870), .B1(new_n890), .B2(new_n217), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT58), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n892), .B1(new_n870), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n870), .B1(new_n893), .B2(new_n892), .C1(new_n890), .C2(new_n217), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1344gat));
  NAND3_X1  g696(.A1(new_n869), .A2(new_n218), .A3(new_n636), .ZN(new_n898));
  NOR3_X1   g697(.A1(new_n883), .A2(new_n887), .A3(new_n889), .ZN(new_n899));
  AOI211_X1 g698(.A(KEYINPUT59), .B(new_n218), .C1(new_n899), .C2(new_n636), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT59), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT118), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n882), .A2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT118), .B(new_n872), .C1(new_n881), .C2(new_n607), .ZN(new_n904));
  NAND4_X1  g703(.A1(new_n903), .A2(new_n871), .A3(new_n285), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n886), .A2(KEYINPUT57), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n905), .A2(new_n636), .A3(new_n888), .A4(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n901), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n898), .B1(new_n900), .B2(new_n908), .ZN(G1345gat));
  AND3_X1   g708(.A1(new_n846), .A2(new_n607), .A3(new_n868), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n911));
  AOI21_X1  g710(.A(G155gat), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n912), .B1(new_n911), .B2(new_n910), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n899), .A2(G155gat), .A3(new_n607), .ZN(new_n914));
  AND2_X1   g713(.A1(new_n913), .A2(new_n914), .ZN(G1346gat));
  INV_X1    g714(.A(G162gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n869), .A2(new_n916), .A3(new_n583), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT120), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n917), .B(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n899), .A2(new_n583), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n916), .B2(new_n920), .ZN(G1347gat));
  AND3_X1   g720(.A1(new_n885), .A2(KEYINPUT121), .A3(new_n340), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT121), .B1(new_n885), .B2(new_n340), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n472), .A2(new_n436), .A3(new_n524), .ZN(new_n925));
  INV_X1    g724(.A(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n924), .A2(new_n661), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n340), .A2(new_n436), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n777), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n472), .B(new_n929), .C1(new_n843), .C2(new_n844), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT122), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n885), .A2(new_n932), .A3(new_n472), .A4(new_n929), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n766), .A2(new_n370), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n927), .A2(new_n370), .B1(new_n934), .B2(new_n935), .ZN(G1348gat));
  NOR2_X1   g735(.A1(new_n637), .A2(new_n369), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n931), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  OR2_X1    g737(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n636), .B(new_n926), .C1(new_n922), .C2(new_n923), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n940), .A2(new_n365), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n938), .A2(KEYINPUT123), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n939), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n939), .A2(new_n941), .A3(KEYINPUT124), .A4(new_n942), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(G1349gat));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n607), .A3(new_n933), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n931), .A2(KEYINPUT125), .A3(new_n933), .A4(new_n607), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n950), .A2(G183gat), .A3(new_n951), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n607), .A2(new_n344), .A3(new_n346), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n924), .A2(new_n926), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(KEYINPUT60), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT60), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n952), .A2(new_n957), .A3(new_n954), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1350gat));
  NOR2_X1   g758(.A1(new_n692), .A2(G190gat), .ZN(new_n960));
  OAI211_X1 g759(.A(new_n926), .B(new_n960), .C1(new_n922), .C2(new_n923), .ZN(new_n961));
  OR2_X1    g760(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(KEYINPUT126), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT61), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT127), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n931), .A2(new_n583), .A3(new_n933), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n965), .B1(new_n966), .B2(G190gat), .ZN(new_n967));
  AOI22_X1  g766(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n966), .A2(new_n965), .A3(G190gat), .ZN(new_n969));
  OR2_X1    g768(.A1(new_n967), .A2(new_n964), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n740), .A2(new_n472), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n436), .B(new_n972), .C1(new_n922), .C2(new_n923), .ZN(new_n973));
  INV_X1    g772(.A(new_n973), .ZN(new_n974));
  AOI21_X1  g773(.A(G197gat), .B1(new_n974), .B2(new_n661), .ZN(new_n975));
  AND2_X1   g774(.A1(new_n905), .A2(new_n906), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n740), .A2(new_n928), .ZN(new_n977));
  AND2_X1   g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n766), .A2(new_n653), .ZN(new_n979));
  AOI21_X1  g778(.A(new_n975), .B1(new_n978), .B2(new_n979), .ZN(G1352gat));
  NOR3_X1   g779(.A1(new_n973), .A2(G204gat), .A3(new_n637), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT62), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n905), .A2(new_n636), .A3(new_n906), .A4(new_n977), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n984), .A2(G204gat), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n981), .A2(new_n982), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n983), .A2(new_n985), .A3(new_n986), .ZN(G1353gat));
  NAND3_X1  g786(.A1(new_n974), .A2(new_n236), .A3(new_n607), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n905), .A2(new_n607), .A3(new_n906), .A4(new_n977), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(G1354gat));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n583), .A3(new_n977), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(G218gat), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n974), .A2(new_n237), .A3(new_n583), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1355gat));
endmodule


