//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n555, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT65), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n461), .A2(G137), .A3(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n464), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT66), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n465), .A2(new_n468), .A3(G101), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n471), .A2(new_n473), .A3(G125), .ZN(new_n474));
  NAND2_X1  g049(.A1(G113), .A2(G2104), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n462), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n470), .A2(new_n476), .ZN(G160));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n461), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n471), .A2(new_n473), .A3(new_n480), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(new_n462), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(G124), .ZN(new_n486));
  OAI21_X1  g061(.A(new_n479), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n483), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n487), .B1(G136), .B2(new_n488), .ZN(G162));
  NAND4_X1  g064(.A1(new_n471), .A2(new_n473), .A3(G138), .A4(new_n462), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n461), .A2(KEYINPUT69), .A3(G138), .A4(new_n462), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n490), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT68), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n462), .A2(G114), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g075(.A1(G102), .A2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n501), .A2(new_n503), .A3(KEYINPUT68), .A4(G2104), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n461), .A2(G126), .A3(G2105), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n494), .A2(new_n496), .A3(new_n505), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT6), .A2(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(new_n511), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n509), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT5), .A2(G543), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n513), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n525));
  OR3_X1    g100(.A1(new_n521), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n521), .B2(new_n524), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n526), .A2(new_n527), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT7), .ZN(new_n530));
  INV_X1    g105(.A(new_n512), .ZN(new_n531));
  INV_X1    g106(.A(G51), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(new_n516), .A2(new_n517), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n514), .A2(G89), .ZN(new_n535));
  NAND2_X1  g110(.A1(G63), .A2(G651), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n533), .A2(new_n537), .ZN(G168));
  NAND2_X1  g113(.A1(new_n512), .A2(G52), .ZN(new_n539));
  INV_X1    g114(.A(G90), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n539), .B1(new_n519), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n542), .A2(new_n523), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(G171));
  NAND2_X1  g119(.A1(new_n512), .A2(G43), .ZN(new_n545));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n519), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n523), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT71), .ZN(new_n551));
  OR3_X1    g126(.A1(new_n547), .A2(new_n549), .A3(KEYINPUT71), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n531), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n512), .A2(new_n562), .A3(G53), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n510), .A2(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(G91), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT72), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n534), .B2(new_n569), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n567), .B1(new_n570), .B2(G651), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n572));
  NOR3_X1   g147(.A1(new_n572), .A2(KEYINPUT72), .A3(new_n523), .ZN(new_n573));
  OAI211_X1 g148(.A(new_n564), .B(new_n566), .C1(new_n571), .C2(new_n573), .ZN(G299));
  INV_X1    g149(.A(G171), .ZN(G301));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n565), .A2(G87), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n512), .A2(G49), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  AOI22_X1  g156(.A1(new_n565), .A2(G86), .B1(new_n512), .B2(G48), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n516), .B2(new_n517), .ZN(new_n584));
  AND2_X1   g159(.A1(G73), .A2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(G651), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n565), .A2(G85), .B1(new_n512), .B2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n523), .B2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n592));
  AND3_X1   g167(.A1(new_n565), .A2(new_n592), .A3(G92), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n592), .B1(new_n565), .B2(G92), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT10), .ZN(new_n595));
  OR3_X1    g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n593), .B2(new_n594), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n534), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n600), .A2(G651), .B1(G54), .B2(new_n512), .ZN(new_n601));
  AND3_X1   g176(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G284));
  OAI21_X1  g178(.A(new_n591), .B1(new_n602), .B2(G868), .ZN(G321));
  NAND2_X1  g179(.A1(G286), .A2(G868), .ZN(new_n605));
  INV_X1    g180(.A(G299), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n605), .B1(new_n606), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n602), .B1(new_n609), .B2(G860), .ZN(G148));
  OAI21_X1  g185(.A(KEYINPUT74), .B1(new_n553), .B2(G868), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n612), .A2(G559), .ZN(new_n613));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  NOR2_X1   g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n611), .B(KEYINPUT74), .S(new_n615), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n461), .A2(new_n465), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(G2100), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n488), .A2(G135), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n484), .A2(G123), .ZN(new_n623));
  OR2_X1    g198(.A1(G99), .A2(G2105), .ZN(new_n624));
  OAI211_X1 g199(.A(new_n624), .B(G2104), .C1(G111), .C2(new_n462), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n622), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  OR2_X1    g201(.A1(new_n626), .A2(G2096), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n627), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(G14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n636), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G1341), .B(G1348), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n630), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n641), .A2(new_n642), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n644), .A2(KEYINPUT75), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(KEYINPUT75), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(KEYINPUT76), .B(KEYINPUT18), .Z(new_n649));
  XOR2_X1   g224(.A(G2084), .B(G2090), .Z(new_n650));
  XNOR2_X1  g225(.A(G2067), .B(G2678), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  INV_X1    g231(.A(new_n649), .ZN(new_n657));
  AOI21_X1  g232(.A(new_n656), .B1(new_n652), .B2(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT77), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n659), .B(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1971), .B(G1976), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT19), .ZN(new_n664));
  XOR2_X1   g239(.A(G1956), .B(G2474), .Z(new_n665));
  XOR2_X1   g240(.A(G1961), .B(G1966), .Z(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AND2_X1   g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n665), .A2(new_n666), .ZN(new_n669));
  NOR3_X1   g244(.A1(new_n664), .A2(new_n669), .A3(new_n667), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n669), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT78), .B(KEYINPUT20), .Z(new_n672));
  AOI211_X1 g247(.A(new_n668), .B(new_n670), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n673), .B1(new_n671), .B2(new_n672), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT79), .ZN(new_n675));
  XOR2_X1   g250(.A(G1981), .B(G1986), .Z(new_n676));
  XNOR2_X1  g251(.A(G1991), .B(G1996), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n675), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G23), .ZN(new_n683));
  INV_X1    g258(.A(G288), .ZN(new_n684));
  OAI21_X1  g259(.A(new_n683), .B1(new_n684), .B2(new_n682), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT33), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G1976), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n682), .A2(KEYINPUT81), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n682), .A2(KEYINPUT81), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(G22), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(G166), .B2(new_n690), .ZN(new_n692));
  INV_X1    g267(.A(G1971), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G6), .A2(G16), .ZN(new_n695));
  INV_X1    g270(.A(G305), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT32), .B(G1981), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n687), .A2(new_n694), .A3(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n488), .A2(G131), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n484), .A2(G119), .ZN(new_n705));
  OR2_X1    g280(.A1(G95), .A2(G2105), .ZN(new_n706));
  OAI211_X1 g281(.A(new_n706), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n704), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n703), .B1(new_n709), .B2(new_n702), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT80), .Z(new_n711));
  XOR2_X1   g286(.A(KEYINPUT35), .B(G1991), .Z(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n700), .A2(KEYINPUT34), .ZN(new_n714));
  INV_X1    g289(.A(new_n690), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n715), .A2(G24), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n716), .B(KEYINPUT82), .Z(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G290), .B2(new_n690), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1986), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT36), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n719), .B1(KEYINPUT83), .B2(new_n720), .ZN(new_n721));
  NOR4_X1   g296(.A1(new_n701), .A2(new_n713), .A3(new_n714), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(KEYINPUT83), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n702), .A2(G35), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(G162), .B2(new_n702), .ZN(new_n727));
  XNOR2_X1  g302(.A(KEYINPUT29), .B(G2090), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n727), .B(new_n728), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n612), .A2(G16), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n682), .A2(G4), .ZN(new_n732));
  AND2_X1   g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n682), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n682), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n736), .A2(G1961), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT87), .Z(new_n738));
  INV_X1    g313(.A(KEYINPUT24), .ZN(new_n739));
  INV_X1    g314(.A(G34), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G160), .B2(new_n702), .ZN(new_n743));
  OAI22_X1  g318(.A1(new_n626), .A2(new_n702), .B1(G2084), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G2084), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(new_n736), .B2(G1961), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR2_X1   g322(.A1(G168), .A2(new_n682), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n682), .B2(G21), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT84), .B(G1966), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g326(.A(KEYINPUT31), .B(G11), .ZN(new_n752));
  INV_X1    g327(.A(KEYINPUT30), .ZN(new_n753));
  AND3_X1   g328(.A1(new_n753), .A2(KEYINPUT86), .A3(G28), .ZN(new_n754));
  AOI21_X1  g329(.A(KEYINPUT86), .B1(new_n753), .B2(G28), .ZN(new_n755));
  OAI221_X1 g330(.A(new_n702), .B1(new_n753), .B2(G28), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NAND4_X1  g331(.A1(new_n747), .A2(new_n751), .A3(new_n752), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(G164), .A2(G29), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G27), .B2(G29), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT88), .B(G2078), .Z(new_n760));
  AOI211_X1 g335(.A(new_n738), .B(new_n757), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n690), .A2(G19), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n553), .B2(new_n690), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1341), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n702), .A2(G26), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT28), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n488), .A2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n484), .A2(G128), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n462), .A2(G116), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(G29), .ZN(new_n772));
  INV_X1    g347(.A(G2067), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n733), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(G1348), .B2(new_n775), .ZN(new_n776));
  NAND4_X1  g351(.A1(new_n734), .A2(new_n761), .A3(new_n764), .A4(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n749), .A2(new_n750), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(KEYINPUT85), .Z(new_n779));
  NAND2_X1  g354(.A1(new_n488), .A2(G139), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n781));
  INV_X1    g356(.A(KEYINPUT25), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  AOI22_X1  g358(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n784));
  OAI211_X1 g359(.A(new_n780), .B(new_n783), .C1(new_n462), .C2(new_n784), .ZN(new_n785));
  MUX2_X1   g360(.A(G33), .B(new_n785), .S(G29), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2072), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n759), .A2(new_n760), .ZN(new_n788));
  NOR3_X1   g363(.A1(new_n779), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  INV_X1    g364(.A(G1996), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n488), .A2(G141), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n484), .A2(G129), .ZN(new_n792));
  NAND3_X1  g367(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT26), .ZN(new_n794));
  OR2_X1    g369(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  AOI22_X1  g371(.A1(new_n795), .A2(new_n796), .B1(G105), .B2(new_n465), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n791), .A2(new_n792), .A3(new_n797), .ZN(new_n798));
  MUX2_X1   g373(.A(G32), .B(new_n798), .S(G29), .Z(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(KEYINPUT27), .Z(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n789), .B1(new_n790), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n800), .A2(G1996), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n715), .A2(G20), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(KEYINPUT89), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT23), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n682), .B2(new_n606), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G1956), .ZN(new_n808));
  NOR4_X1   g383(.A1(new_n777), .A2(new_n802), .A3(new_n803), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g384(.A1(new_n724), .A2(new_n725), .A3(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(new_n512), .A2(G55), .ZN(new_n812));
  INV_X1    g387(.A(G93), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n812), .B1(new_n519), .B2(new_n813), .ZN(new_n814));
  AOI22_X1  g389(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(new_n523), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(G860), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT37), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n817), .B1(new_n551), .B2(new_n552), .ZN(new_n821));
  INV_X1    g396(.A(new_n817), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n550), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n612), .A2(new_n609), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(KEYINPUT90), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n818), .B1(new_n828), .B2(KEYINPUT39), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n820), .B1(new_n830), .B2(new_n831), .ZN(G145));
  XNOR2_X1  g407(.A(new_n771), .B(new_n507), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n619), .B(KEYINPUT94), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n837));
  OR3_X1    g412(.A1(new_n462), .A2(KEYINPUT93), .A3(G118), .ZN(new_n838));
  OAI21_X1  g413(.A(KEYINPUT93), .B1(new_n462), .B2(G118), .ZN(new_n839));
  OR2_X1    g414(.A1(G106), .A2(G2105), .ZN(new_n840));
  NAND4_X1  g415(.A1(new_n838), .A2(G2104), .A3(new_n839), .A4(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n488), .A2(G142), .ZN(new_n843));
  OR2_X1    g418(.A1(new_n843), .A2(KEYINPUT91), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n843), .A2(KEYINPUT91), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n484), .A2(G130), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(KEYINPUT92), .Z(new_n848));
  AOI21_X1  g423(.A(new_n837), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n846), .A2(new_n848), .A3(new_n837), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n850), .A2(new_n708), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(new_n851), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n709), .B1(new_n853), .B2(new_n849), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n785), .B(new_n798), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n855), .B1(new_n852), .B2(new_n854), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n836), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n852), .A2(new_n854), .ZN(new_n860));
  INV_X1    g435(.A(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n862), .A2(new_n835), .A3(new_n856), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n859), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n626), .B(G160), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(G162), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n864), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(G37), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n859), .A2(new_n863), .A3(new_n866), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n868), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n613), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(KEYINPUT96), .B1(new_n612), .B2(G559), .ZN(new_n876));
  AND3_X1   g451(.A1(new_n875), .A2(new_n824), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n824), .B1(new_n876), .B2(new_n875), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT97), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n612), .B1(new_n880), .B2(new_n606), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n880), .B2(new_n606), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n612), .A2(KEYINPUT97), .A3(G299), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n873), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(KEYINPUT41), .A3(new_n883), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT41), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n879), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n884), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n890), .B(KEYINPUT98), .C1(new_n877), .C2(new_n878), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n885), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G166), .B(G288), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n696), .B(G290), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g471(.A1(G303), .A2(G288), .ZN(new_n897));
  NOR2_X1   g472(.A1(G166), .A2(new_n684), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT42), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(KEYINPUT42), .B1(new_n896), .B2(new_n899), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n892), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n904), .A2(new_n885), .A3(new_n889), .A4(new_n891), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(G868), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(KEYINPUT99), .B1(new_n822), .B2(new_n614), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT99), .A4(G868), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n910), .A2(KEYINPUT100), .A3(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(KEYINPUT100), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(G295));
  AND2_X1   g489(.A1(new_n910), .A2(new_n911), .ZN(G331));
  AND2_X1   g490(.A1(new_n888), .A2(new_n886), .ZN(new_n916));
  NAND2_X1  g491(.A1(G301), .A2(KEYINPUT101), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n918));
  NAND2_X1  g493(.A1(G171), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n917), .A2(G286), .A3(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(G171), .A2(new_n918), .A3(G168), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n922), .B1(new_n821), .B2(new_n823), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT102), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OR2_X1    g500(.A1(new_n821), .A2(new_n823), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(KEYINPUT102), .A3(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n824), .A2(new_n921), .A3(new_n920), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT103), .ZN(new_n930));
  OR3_X1    g505(.A1(new_n926), .A2(KEYINPUT103), .A3(new_n922), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT104), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n929), .A2(new_n923), .A3(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n926), .A2(KEYINPUT104), .A3(new_n922), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n916), .A2(new_n932), .B1(new_n890), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n900), .ZN(new_n938));
  AOI21_X1  g513(.A(G37), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n928), .A2(new_n890), .A3(new_n930), .A4(new_n931), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n888), .A2(new_n886), .A3(new_n934), .A4(new_n935), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n940), .B1(new_n943), .B2(new_n900), .ZN(new_n944));
  AOI211_X1 g519(.A(KEYINPUT105), .B(new_n938), .C1(new_n941), .C2(new_n942), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n939), .B(KEYINPUT43), .C1(new_n944), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n916), .A2(new_n932), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n936), .A2(new_n890), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n938), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n869), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n937), .A2(new_n938), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n946), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT44), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n939), .B(new_n947), .C1(new_n944), .C2(new_n945), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT43), .B1(new_n951), .B2(new_n952), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n955), .A2(new_n960), .ZN(G397));
  INV_X1    g536(.A(G1384), .ZN(new_n962));
  AND3_X1   g537(.A1(new_n492), .A2(new_n493), .A3(KEYINPUT4), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT45), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(G160), .A2(G40), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n771), .B(G2067), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n798), .B(new_n790), .ZN(new_n972));
  OR2_X1    g547(.A1(new_n709), .A2(new_n712), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n709), .A2(new_n712), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n971), .A2(new_n972), .A3(new_n973), .A4(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(G290), .B(G1986), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n969), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G40), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n470), .A2(new_n978), .A3(new_n476), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n507), .A2(new_n979), .A3(new_n962), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(G2067), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n496), .A2(new_n505), .A3(new_n506), .ZN(new_n983));
  AOI21_X1  g558(.A(G1384), .B1(new_n983), .B2(new_n494), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT50), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(new_n986));
  OAI211_X1 g561(.A(new_n985), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT106), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT106), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n984), .A2(new_n989), .A3(new_n985), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n986), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(KEYINPUT60), .B(new_n982), .C1(new_n991), .C2(G1348), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT118), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n968), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n989), .B1(new_n984), .B2(new_n985), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n987), .A2(KEYINPUT106), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n981), .B1(new_n997), .B2(new_n730), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT118), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT60), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n993), .A2(new_n602), .A3(new_n1000), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n992), .A2(KEYINPUT118), .A3(new_n612), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n998), .A2(KEYINPUT60), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI211_X1 g579(.A(KEYINPUT114), .B(new_n566), .C1(new_n571), .C2(new_n573), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT57), .ZN(new_n1006));
  NAND3_X1  g581(.A1(G299), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n570), .A2(new_n567), .A3(G651), .ZN(new_n1008));
  OAI21_X1  g583(.A(KEYINPUT72), .B1(new_n572), .B2(new_n523), .ZN(new_n1009));
  AOI22_X1  g584(.A1(new_n1008), .A2(new_n1009), .B1(G91), .B2(new_n565), .ZN(new_n1010));
  OAI211_X1 g585(.A(new_n1010), .B(new_n564), .C1(KEYINPUT114), .C2(KEYINPUT57), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(KEYINPUT113), .B(G1956), .Z(new_n1013));
  AOI21_X1  g588(.A(new_n1013), .B1(new_n994), .B2(new_n987), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n962), .ZN(new_n1015));
  XNOR2_X1  g590(.A(KEYINPUT56), .B(G2072), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT115), .ZN(new_n1017));
  AND4_X1   g592(.A1(new_n967), .A2(new_n979), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1012), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n967), .A2(new_n979), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n965), .A2(KEYINPUT50), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1022), .A2(new_n979), .A3(new_n987), .ZN(new_n1023));
  OAI211_X1 g598(.A(new_n1020), .B(new_n1021), .C1(new_n1023), .C2(new_n1013), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(KEYINPUT61), .A3(new_n1024), .ZN(new_n1025));
  XOR2_X1   g600(.A(KEYINPUT58), .B(G1341), .Z(new_n1026));
  NAND2_X1  g601(.A1(new_n980), .A2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(KEYINPUT116), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n967), .A2(new_n790), .A3(new_n1015), .A4(new_n979), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n980), .A2(new_n1030), .A3(new_n1026), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(new_n1029), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT59), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1032), .A2(new_n1033), .A3(new_n553), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(new_n1032), .B2(new_n553), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1025), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI211_X1 g611(.A(KEYINPUT117), .B(KEYINPUT61), .C1(new_n1019), .C2(new_n1024), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1019), .A2(new_n1024), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n1039), .B2(KEYINPUT61), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1004), .A2(new_n1038), .A3(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT119), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1019), .B1(new_n998), .B2(new_n612), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(new_n1024), .ZN(new_n1044));
  AND3_X1   g619(.A1(new_n1041), .A2(new_n1042), .A3(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1042), .B1(new_n1041), .B2(new_n1044), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n526), .A2(G8), .A3(new_n527), .ZN(new_n1047));
  XNOR2_X1  g622(.A(KEYINPUT108), .B(KEYINPUT55), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1047), .B(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT107), .B(G2090), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n994), .A2(new_n987), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT111), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1023), .A2(KEYINPUT111), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n967), .A2(new_n979), .A3(new_n1015), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1054), .A2(new_n1055), .B1(new_n693), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G8), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1049), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n684), .A2(G1976), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n980), .A2(G8), .A3(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(KEYINPUT52), .ZN(new_n1062));
  INV_X1    g637(.A(G1976), .ZN(new_n1063));
  AOI21_X1  g638(.A(KEYINPUT52), .B1(G288), .B2(new_n1063), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n980), .A2(G8), .A3(new_n1060), .A4(new_n1064), .ZN(new_n1065));
  XNOR2_X1  g640(.A(KEYINPUT109), .B(G1981), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n582), .A2(new_n586), .A3(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT110), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT110), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n582), .A2(new_n1069), .A3(new_n586), .A4(new_n1066), .ZN(new_n1070));
  AOI22_X1  g645(.A1(new_n1068), .A2(new_n1070), .B1(G1981), .B2(G305), .ZN(new_n1071));
  OAI211_X1 g646(.A(G8), .B(new_n980), .C1(new_n1071), .C2(KEYINPUT49), .ZN(new_n1072));
  AND2_X1   g647(.A1(new_n1071), .A2(KEYINPUT49), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1062), .B(new_n1065), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n994), .B(new_n1050), .C1(new_n995), .C2(new_n996), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1056), .A2(new_n693), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1058), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(new_n1049), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1074), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1059), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g655(.A(G2078), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n967), .A2(new_n1081), .A3(new_n1015), .A4(new_n979), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1084), .A2(KEYINPUT123), .ZN(new_n1085));
  INV_X1    g660(.A(G1961), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n997), .A2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1082), .A2(new_n1089), .A3(new_n1083), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1085), .A2(new_n1087), .A3(new_n1088), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n470), .A2(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n470), .A2(new_n1095), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1081), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1098));
  NOR4_X1   g673(.A1(new_n1096), .A2(new_n1097), .A3(new_n476), .A4(new_n1098), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(new_n967), .A3(new_n1015), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1085), .A2(new_n1087), .A3(new_n1090), .A4(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(G171), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1080), .B1(new_n1094), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT125), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(new_n1101), .B2(G171), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1091), .A2(G171), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1101), .A2(new_n1104), .A3(G171), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1093), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(G2084), .ZN(new_n1110));
  OAI211_X1 g685(.A(new_n1110), .B(new_n994), .C1(new_n995), .C2(new_n996), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1056), .A2(new_n750), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1058), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(G286), .A2(G8), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT120), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1115), .A2(KEYINPUT51), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NOR2_X1   g695(.A1(new_n1113), .A2(KEYINPUT121), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT122), .B(new_n1116), .C1(new_n1120), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1113), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT121), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(new_n1118), .A4(new_n1119), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1117), .A2(new_n1115), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1122), .A2(new_n1127), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1103), .A2(new_n1109), .A3(new_n1129), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1045), .A2(new_n1046), .A3(new_n1130), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1080), .A2(new_n1106), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1128), .ZN(new_n1133));
  AOI211_X1 g708(.A(new_n1124), .B(new_n1058), .C1(new_n1111), .C2(new_n1112), .ZN(new_n1134));
  INV_X1    g709(.A(new_n1119), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1121), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(new_n1126), .ZN(new_n1137));
  AOI21_X1  g712(.A(KEYINPUT62), .B1(new_n1137), .B2(new_n1122), .ZN(new_n1138));
  AND4_X1   g713(.A1(KEYINPUT62), .A2(new_n1122), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1132), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  OR2_X1    g715(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1141));
  NOR2_X1   g716(.A1(G288), .A2(G1976), .ZN(new_n1142));
  AOI22_X1  g717(.A1(new_n1141), .A2(new_n1142), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n980), .A2(G8), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1078), .A2(new_n1077), .ZN(new_n1145));
  OAI22_X1  g720(.A1(new_n1143), .A2(new_n1144), .B1(new_n1145), .B2(new_n1074), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1123), .A2(G286), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1059), .A2(new_n1079), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT112), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT63), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1059), .A2(new_n1079), .A3(new_n1147), .A4(KEYINPUT112), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  OR2_X1    g728(.A1(new_n1078), .A2(new_n1077), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1079), .A2(new_n1147), .A3(new_n1154), .A4(KEYINPUT63), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1146), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1140), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n977), .B1(new_n1131), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n969), .B1(new_n970), .B2(new_n798), .ZN(new_n1159));
  NOR3_X1   g734(.A1(new_n967), .A2(G1996), .A3(new_n968), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(KEYINPUT46), .ZN(new_n1161));
  OR2_X1    g736(.A1(new_n1160), .A2(KEYINPUT46), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1159), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  XOR2_X1   g738(.A(new_n1163), .B(KEYINPUT126), .Z(new_n1164));
  XNOR2_X1  g739(.A(new_n1164), .B(KEYINPUT47), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n971), .A2(new_n972), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n1166), .A2(new_n974), .B1(G2067), .B2(new_n771), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(new_n969), .ZN(new_n1168));
  AND2_X1   g743(.A1(new_n975), .A2(new_n969), .ZN(new_n1169));
  NOR2_X1   g744(.A1(G290), .A2(G1986), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n969), .A2(new_n1170), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n1171), .B(KEYINPUT48), .Z(new_n1172));
  OAI21_X1  g747(.A(new_n1168), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1165), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1158), .A2(new_n1174), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g750(.A1(G229), .A2(new_n459), .A3(G227), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n1177), .A2(new_n647), .ZN(new_n1178));
  NAND2_X1  g752(.A1(new_n1178), .A2(KEYINPUT127), .ZN(new_n1179));
  INV_X1    g753(.A(KEYINPUT127), .ZN(new_n1180));
  NAND3_X1  g754(.A1(new_n1177), .A2(new_n1180), .A3(new_n647), .ZN(new_n1181));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g756(.A1(new_n958), .A2(new_n1182), .A3(new_n871), .ZN(G225));
  INV_X1    g757(.A(G225), .ZN(G308));
endmodule


