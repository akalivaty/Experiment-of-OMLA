//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n969, new_n970, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT90), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n206), .B(G8gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n213), .B(KEYINPUT85), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT15), .ZN(new_n215));
  OR3_X1    g014(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT88), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(KEYINPUT87), .Z(new_n222));
  NOR2_X1   g021(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n215), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  OAI211_X1 g024(.A(KEYINPUT86), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(new_n218), .B2(KEYINPUT86), .ZN(new_n227));
  OAI211_X1 g026(.A(new_n214), .B(KEYINPUT15), .C1(new_n227), .C2(new_n222), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n209), .A2(new_n212), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G229gat), .A2(G233gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(KEYINPUT89), .A2(KEYINPUT17), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT89), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT17), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  AND3_X1   g034(.A1(new_n229), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n235), .B1(new_n229), .B2(new_n232), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n230), .B(new_n231), .C1(new_n238), .C2(new_n210), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n230), .ZN(new_n242));
  AND2_X1   g041(.A1(new_n225), .A2(new_n228), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n243), .A2(new_n233), .A3(new_n234), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n229), .A2(new_n232), .A3(new_n235), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n246), .B2(new_n208), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(KEYINPUT18), .A3(new_n231), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n209), .A2(new_n212), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(new_n243), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(new_n230), .ZN(new_n251));
  XOR2_X1   g050(.A(new_n231), .B(KEYINPUT91), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n252), .B(KEYINPUT13), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n241), .A2(new_n248), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G197gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(KEYINPUT11), .ZN(new_n258));
  INV_X1    g057(.A(G169gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n260), .B(KEYINPUT12), .Z(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(new_n261), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n263), .A2(new_n241), .A3(new_n254), .A4(new_n248), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT92), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT92), .B1(new_n262), .B2(new_n264), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G197gat), .B(G204gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT22), .ZN(new_n271));
  INV_X1    g070(.A(G211gat), .ZN(new_n272));
  INV_X1    g071(.A(G218gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G211gat), .B(G218gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n270), .A3(new_n274), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G183gat), .A2(G190gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(KEYINPUT24), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(KEYINPUT65), .A3(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n284), .B(new_n286), .C1(new_n291), .C2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR3_X1   g094(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n296));
  OAI21_X1  g095(.A(KEYINPUT23), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(G176gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n259), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT23), .ZN(new_n300));
  NOR2_X1   g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n299), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n293), .A2(new_n297), .A3(new_n303), .A4(KEYINPUT25), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n299), .B1(KEYINPUT23), .B2(new_n301), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n289), .A2(KEYINPUT24), .A3(new_n281), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n302), .A2(new_n300), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n281), .A2(KEYINPUT24), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n305), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n304), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n287), .A2(KEYINPUT27), .ZN(new_n313));
  AOI21_X1  g112(.A(G190gat), .B1(new_n313), .B2(KEYINPUT67), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT27), .ZN(new_n315));
  OR3_X1    g114(.A1(new_n315), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT28), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(G183gat), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n314), .A2(new_n316), .A3(new_n317), .A4(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(new_n318), .A3(new_n288), .ZN(new_n320));
  AOI21_X1  g119(.A(new_n282), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT26), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n323), .B1(new_n295), .B2(new_n296), .ZN(new_n324));
  INV_X1    g123(.A(new_n299), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT68), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n326), .B1(new_n301), .B2(new_n323), .ZN(new_n327));
  OAI211_X1 g126(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n322), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n312), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT76), .ZN(new_n332));
  NAND2_X1  g131(.A1(G226gat), .A2(G233gat), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n331), .A2(new_n332), .A3(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n304), .A2(new_n311), .B1(new_n322), .B2(new_n329), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT76), .B1(new_n336), .B2(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT69), .B1(new_n322), .B2(new_n329), .ZN(new_n341));
  AND4_X1   g140(.A1(KEYINPUT69), .A2(new_n329), .A3(new_n321), .A4(new_n319), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n312), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT69), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n321), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n327), .A2(new_n328), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT64), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(new_n259), .A3(new_n298), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT26), .B1(new_n350), .B2(new_n294), .ZN(new_n351));
  NOR3_X1   g150(.A1(new_n348), .A2(new_n351), .A3(new_n299), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n346), .B1(new_n347), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n329), .A2(KEYINPUT69), .A3(new_n321), .A4(new_n319), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n355), .A2(KEYINPUT74), .A3(new_n312), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n340), .B1(new_n345), .B2(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n280), .B(new_n339), .C1(new_n357), .C2(new_n334), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n345), .A2(new_n334), .A3(new_n356), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n278), .A2(new_n279), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT29), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n331), .A2(new_n361), .A3(new_n333), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G8gat), .B(G36gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT77), .ZN(new_n366));
  INV_X1    g165(.A(G64gat), .ZN(new_n367));
  XNOR2_X1  g166(.A(new_n366), .B(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(G92gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n358), .A2(new_n363), .A3(new_n370), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(KEYINPUT30), .A3(new_n373), .ZN(new_n374));
  AOI211_X1 g173(.A(KEYINPUT30), .B(new_n370), .C1(new_n358), .C2(new_n363), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT70), .ZN(new_n377));
  INV_X1    g176(.A(G120gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n378), .A2(G113gat), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G120gat), .ZN(new_n381));
  AOI21_X1  g180(.A(KEYINPUT1), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G127gat), .B(G134gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n377), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(G127gat), .A2(G134gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(G127gat), .A2(G134gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G113gat), .B(G120gat), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n387), .B(KEYINPUT70), .C1(new_n388), .C2(KEYINPUT1), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT71), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n380), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n391), .A2(new_n379), .A3(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n387), .A2(KEYINPUT1), .ZN(new_n394));
  AOI22_X1  g193(.A1(new_n384), .A2(new_n389), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  INV_X1    g195(.A(G141gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(G148gat), .ZN(new_n398));
  INV_X1    g197(.A(G148gat), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G141gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n398), .A2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(G155gat), .B(G162gat), .ZN(new_n402));
  NAND2_X1  g201(.A1(G155gat), .A2(G162gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT2), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n396), .A2(new_n401), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT78), .B1(new_n398), .B2(new_n400), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n402), .B1(new_n406), .B2(new_n404), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n395), .A2(KEYINPUT80), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT80), .B1(new_n395), .B2(new_n408), .ZN(new_n410));
  OAI22_X1  g209(.A1(new_n409), .A2(new_n410), .B1(new_n408), .B2(new_n395), .ZN(new_n411));
  NAND2_X1  g210(.A1(G225gat), .A2(G233gat), .ZN(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT79), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n415), .B1(new_n405), .B2(new_n407), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n399), .A2(G141gat), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n397), .A2(G148gat), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n396), .B(new_n404), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n402), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n402), .A3(new_n404), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(KEYINPUT79), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(KEYINPUT4), .A3(new_n395), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n409), .A2(new_n410), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n425), .B1(new_n426), .B2(KEYINPUT4), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n384), .A2(new_n389), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n394), .A2(new_n393), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT3), .B1(new_n405), .B2(new_n407), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT3), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n421), .A2(new_n432), .A3(new_n422), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n412), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT5), .B(new_n414), .C1(new_n427), .C2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT81), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(KEYINPUT4), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n424), .A2(new_n395), .ZN(new_n439));
  AOI22_X1  g238(.A1(new_n426), .A2(KEYINPUT4), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n413), .A2(KEYINPUT5), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n437), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n438), .A2(new_n439), .ZN(new_n443));
  INV_X1    g242(.A(new_n410), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n395), .A2(new_n408), .A3(KEYINPUT80), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT4), .A3(new_n445), .ZN(new_n446));
  AND4_X1   g245(.A1(new_n437), .A2(new_n443), .A3(new_n446), .A4(new_n441), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n436), .B1(new_n442), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(G1gat), .B(G29gat), .ZN(new_n449));
  XNOR2_X1  g248(.A(new_n449), .B(KEYINPUT0), .ZN(new_n450));
  XNOR2_X1  g249(.A(new_n450), .B(G57gat), .ZN(new_n451));
  XNOR2_X1  g250(.A(new_n451), .B(G85gat), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n440), .A2(new_n437), .A3(new_n441), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n443), .A2(new_n446), .A3(new_n441), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n452), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n458), .A2(new_n459), .A3(new_n436), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n453), .A2(new_n454), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n459), .B1(new_n458), .B2(new_n436), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT6), .ZN(new_n463));
  AOI22_X1  g262(.A1(new_n374), .A2(new_n376), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT31), .B(G50gat), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n465), .B(G106gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G22gat), .B(G78gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT82), .ZN(new_n470));
  INV_X1    g269(.A(new_n340), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n360), .B1(new_n433), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n421), .A2(KEYINPUT79), .A3(new_n422), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT79), .B1(new_n421), .B2(new_n422), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n432), .B1(new_n280), .B2(new_n340), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(G228gat), .ZN(new_n478));
  INV_X1    g277(.A(G233gat), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n470), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n340), .B1(new_n278), .B2(new_n279), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n416), .B(new_n423), .C1(KEYINPUT3), .C2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n433), .A2(new_n471), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n280), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n480), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(KEYINPUT82), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n481), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n360), .A2(new_n361), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n408), .B1(new_n490), .B2(new_n432), .ZN(new_n491));
  NOR3_X1   g290(.A1(new_n491), .A2(new_n487), .A3(new_n472), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n469), .B1(new_n489), .B2(new_n493), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n468), .B(new_n492), .C1(new_n481), .C2(new_n488), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n467), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g295(.A(KEYINPUT82), .B1(new_n486), .B2(new_n487), .ZN(new_n497));
  AOI211_X1 g296(.A(new_n470), .B(new_n480), .C1(new_n483), .C2(new_n485), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n493), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n468), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n489), .A2(new_n469), .A3(new_n493), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(new_n466), .A3(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n343), .A2(new_n395), .ZN(new_n504));
  NAND2_X1  g303(.A1(G227gat), .A2(G233gat), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n355), .A2(new_n430), .A3(new_n312), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT32), .ZN(new_n509));
  XOR2_X1   g308(.A(KEYINPUT72), .B(KEYINPUT33), .Z(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G15gat), .B(G43gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G71gat), .ZN(new_n514));
  INV_X1    g313(.A(G99gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n509), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n516), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n508), .B(KEYINPUT32), .C1(new_n511), .C2(new_n518), .ZN(new_n519));
  AND3_X1   g318(.A1(new_n355), .A2(new_n430), .A3(new_n312), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n430), .B1(new_n355), .B2(new_n312), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n505), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT34), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT73), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n523), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  OAI221_X1 g325(.A(new_n505), .B1(new_n524), .B2(new_n523), .C1(new_n520), .C2(new_n521), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  AND3_X1   g327(.A1(new_n517), .A2(new_n519), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n528), .B1(new_n517), .B2(new_n519), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n503), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT84), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT84), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n503), .B(new_n533), .C1(new_n529), .C2(new_n530), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n464), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT83), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n461), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n453), .A2(KEYINPUT83), .A3(new_n454), .A4(new_n460), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(new_n463), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n531), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT35), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n374), .A2(new_n376), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n540), .A2(new_n541), .A3(new_n542), .A4(new_n543), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n440), .A2(new_n412), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT39), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n452), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n411), .A2(new_n413), .ZN(new_n548));
  OAI211_X1 g347(.A(new_n548), .B(KEYINPUT39), .C1(new_n412), .C2(new_n440), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT40), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n550), .A2(new_n462), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(KEYINPUT40), .A3(new_n549), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n374), .A2(new_n376), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT37), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n364), .A2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT38), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n359), .A2(new_n362), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n280), .ZN(new_n558));
  INV_X1    g357(.A(new_n356), .ZN(new_n559));
  AOI21_X1  g358(.A(KEYINPUT74), .B1(new_n355), .B2(new_n312), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n471), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n338), .B1(new_n561), .B2(new_n333), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n558), .B(KEYINPUT37), .C1(new_n562), .C2(new_n280), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n555), .A2(new_n556), .A3(new_n563), .A4(new_n370), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n358), .A2(KEYINPUT37), .A3(new_n363), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT37), .B1(new_n358), .B2(new_n363), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n565), .A2(new_n566), .A3(new_n371), .ZN(new_n567));
  OAI211_X1 g366(.A(new_n372), .B(new_n564), .C1(new_n567), .C2(new_n556), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n553), .B(new_n503), .C1(new_n568), .C2(new_n540), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT36), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(new_n529), .B2(new_n530), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n517), .A2(new_n519), .ZN(new_n572));
  INV_X1    g371(.A(new_n528), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n517), .A2(new_n519), .A3(new_n528), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n574), .A2(KEYINPUT36), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n571), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n461), .A2(new_n463), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n373), .A2(KEYINPUT30), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n370), .B1(new_n358), .B2(new_n363), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n578), .B1(new_n581), .B2(new_n375), .ZN(new_n582));
  INV_X1    g381(.A(new_n503), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n577), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n536), .A2(new_n544), .B1(new_n569), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n367), .A2(G57gat), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n587));
  INV_X1    g386(.A(G57gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n588), .A2(G64gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n586), .A2(KEYINPUT94), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(G71gat), .A2(G78gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT9), .ZN(new_n593));
  NAND2_X1  g392(.A1(G71gat), .A2(G78gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(KEYINPUT93), .A2(KEYINPUT9), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n597), .B1(new_n589), .B2(new_n586), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n598), .A2(new_n592), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n594), .B(KEYINPUT93), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n602), .A2(KEYINPUT21), .ZN(new_n603));
  INV_X1    g402(.A(G127gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n601), .B(KEYINPUT95), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT21), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(new_n249), .ZN(new_n608));
  AND2_X1   g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n605), .A2(new_n608), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n612));
  XNOR2_X1  g411(.A(G155gat), .B(G183gat), .ZN(new_n613));
  XOR2_X1   g412(.A(new_n612), .B(new_n613), .Z(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n611), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G231gat), .A2(G233gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n272), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n614), .B1(new_n609), .B2(new_n610), .ZN(new_n619));
  AND3_X1   g418(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n618), .B1(new_n616), .B2(new_n619), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G85gat), .A2(G92gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT7), .ZN(new_n624));
  NAND2_X1  g423(.A1(G99gat), .A2(G106gat), .ZN(new_n625));
  INV_X1    g424(.A(G85gat), .ZN(new_n626));
  AOI22_X1  g425(.A1(KEYINPUT8), .A2(new_n625), .B1(new_n626), .B2(new_n369), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g427(.A(G99gat), .B(G106gat), .Z(new_n629));
  NOR2_X1   g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(KEYINPUT97), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n629), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT98), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n631), .A2(new_n602), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n632), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n636), .A2(new_n601), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT99), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n631), .A2(new_n633), .A3(new_n638), .A4(new_n602), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n635), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT100), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n635), .A2(new_n637), .A3(new_n645), .A4(new_n639), .ZN(new_n646));
  INV_X1    g445(.A(new_n636), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(KEYINPUT10), .A3(new_n606), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(new_n641), .ZN(new_n650));
  XNOR2_X1  g449(.A(G120gat), .B(G148gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(KEYINPUT101), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n298), .ZN(new_n653));
  INV_X1    g452(.A(G204gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n644), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n655), .ZN(new_n658));
  INV_X1    g457(.A(new_n643), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n642), .B1(new_n646), .B2(new_n648), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(KEYINPUT102), .B(new_n658), .C1(new_n659), .C2(new_n660), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n657), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n647), .B1(new_n244), .B2(new_n245), .ZN(new_n666));
  AND2_X1   g465(.A1(G232gat), .A2(G233gat), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT41), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n668), .B1(new_n636), .B2(new_n243), .ZN(new_n669));
  OAI21_X1  g468(.A(G190gat), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n669), .ZN(new_n671));
  OAI211_X1 g470(.A(new_n288), .B(new_n671), .C1(new_n238), .C2(new_n647), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(new_n273), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n670), .A2(new_n672), .A3(G218gat), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n667), .A2(KEYINPUT41), .ZN(new_n677));
  XNOR2_X1  g476(.A(G134gat), .B(G162gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n677), .B(new_n678), .Z(new_n679));
  NAND4_X1  g478(.A1(new_n674), .A2(new_n675), .A3(new_n676), .A4(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n681));
  INV_X1    g480(.A(new_n679), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g482(.A1(new_n622), .A2(new_n665), .A3(new_n680), .A4(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT103), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n620), .A2(new_n621), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n683), .A2(new_n680), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n689), .A3(new_n665), .ZN(new_n690));
  AOI211_X1 g489(.A(new_n269), .B(new_n585), .C1(new_n685), .C2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n578), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G1gat), .ZN(G1324gat));
  INV_X1    g493(.A(new_n543), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n697));
  AND2_X1   g496(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n207), .B1(new_n691), .B2(new_n695), .ZN(new_n700));
  OAI21_X1  g499(.A(KEYINPUT42), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n701), .B1(KEYINPUT42), .B2(new_n699), .ZN(G1325gat));
  NOR2_X1   g501(.A1(new_n529), .A2(new_n530), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g503(.A(G15gat), .B1(new_n691), .B2(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n577), .A2(G15gat), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n705), .B1(new_n691), .B2(new_n706), .ZN(G1326gat));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n583), .ZN(new_n708));
  XNOR2_X1  g507(.A(KEYINPUT43), .B(G22gat), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n708), .B(new_n709), .ZN(G1327gat));
  INV_X1    g509(.A(new_n657), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n663), .A2(new_n664), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n622), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n262), .A2(new_n264), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT44), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n536), .A2(new_n544), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n568), .A2(new_n540), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n553), .A2(new_n503), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n584), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n719), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n718), .B1(new_n723), .B2(new_n687), .ZN(new_n724));
  INV_X1    g523(.A(new_n687), .ZN(new_n725));
  AOI211_X1 g524(.A(KEYINPUT44), .B(new_n725), .C1(new_n719), .C2(new_n722), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n692), .B(new_n717), .C1(new_n724), .C2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(KEYINPUT105), .ZN(new_n728));
  OAI21_X1  g527(.A(KEYINPUT44), .B1(new_n585), .B2(new_n725), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n723), .A2(new_n718), .A3(new_n687), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT105), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n731), .A2(new_n732), .A3(new_n692), .A4(new_n717), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n728), .A2(G29gat), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g533(.A(new_n725), .B1(new_n719), .B2(new_n722), .ZN(new_n735));
  INV_X1    g534(.A(new_n269), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n578), .A2(G29gat), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n735), .A2(new_n736), .A3(new_n714), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(KEYINPUT104), .ZN(new_n739));
  AOI211_X1 g538(.A(new_n269), .B(new_n725), .C1(new_n719), .C2(new_n722), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT104), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n740), .A2(new_n741), .A3(new_n714), .A4(new_n737), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n739), .A2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT45), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n739), .A2(new_n742), .A3(KEYINPUT45), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT106), .B1(new_n734), .B2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n728), .A2(G29gat), .A3(new_n733), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT106), .ZN(new_n750));
  NAND4_X1  g549(.A1(new_n749), .A2(new_n750), .A3(new_n746), .A4(new_n745), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n748), .A2(new_n751), .ZN(G1328gat));
  AND2_X1   g551(.A1(new_n740), .A2(new_n714), .ZN(new_n753));
  INV_X1    g552(.A(G36gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n754), .A3(new_n695), .ZN(new_n755));
  XOR2_X1   g554(.A(new_n755), .B(KEYINPUT46), .Z(new_n756));
  AND3_X1   g555(.A1(new_n731), .A2(new_n695), .A3(new_n717), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(new_n754), .ZN(G1329gat));
  INV_X1    g557(.A(G43gat), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n753), .A2(KEYINPUT107), .A3(new_n759), .A4(new_n704), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT107), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n740), .A2(new_n759), .A3(new_n714), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(new_n703), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n731), .A2(new_n577), .A3(new_n717), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(G43gat), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT47), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n766), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1330gat));
  NAND3_X1  g570(.A1(new_n731), .A2(new_n583), .A3(new_n717), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n731), .A2(new_n774), .A3(new_n583), .A4(new_n717), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n773), .A2(G50gat), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(G50gat), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n753), .A2(new_n777), .A3(new_n583), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(KEYINPUT48), .A3(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n778), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n780), .B1(G50gat), .B2(new_n772), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(KEYINPUT48), .B2(new_n781), .ZN(G1331gat));
  NOR2_X1   g581(.A1(new_n665), .A2(new_n265), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n723), .A2(new_n688), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n784), .A2(new_n578), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(new_n588), .ZN(G1332gat));
  NOR2_X1   g585(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n543), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  AND2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(G1333gat));
  XOR2_X1   g593(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n795));
  XOR2_X1   g594(.A(new_n703), .B(KEYINPUT110), .Z(new_n796));
  OR3_X1    g595(.A1(new_n784), .A2(G71gat), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n577), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n798), .B1(new_n788), .B2(new_n789), .ZN(new_n799));
  INV_X1    g598(.A(G71gat), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n795), .B(new_n797), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n789), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n577), .B1(new_n803), .B2(new_n787), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G71gat), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n795), .B1(new_n805), .B2(new_n797), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n802), .A2(new_n806), .ZN(G1334gat));
  OAI21_X1  g606(.A(new_n583), .B1(new_n803), .B2(new_n787), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g608(.A1(new_n622), .A2(new_n265), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n735), .A2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n735), .A2(KEYINPUT51), .A3(new_n810), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n665), .A2(new_n578), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n815), .A2(new_n626), .A3(new_n816), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n731), .A2(new_n810), .A3(new_n816), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n817), .B1(new_n818), .B2(new_n626), .ZN(G1336gat));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n665), .A2(G92gat), .A3(new_n543), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g621(.A1(new_n731), .A2(new_n713), .A3(new_n810), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n823), .A2(new_n695), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n820), .B(new_n822), .C1(new_n824), .C2(new_n369), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n369), .B1(new_n823), .B2(new_n695), .ZN(new_n826));
  INV_X1    g625(.A(new_n822), .ZN(new_n827));
  OAI21_X1  g626(.A(KEYINPUT52), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n825), .A2(new_n828), .ZN(G1337gat));
  NAND2_X1  g628(.A1(new_n823), .A2(new_n577), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n823), .A2(KEYINPUT112), .A3(new_n577), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(G99gat), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n815), .A2(new_n515), .A3(new_n704), .A4(new_n713), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1338gat));
  INV_X1    g635(.A(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n823), .B2(new_n583), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n665), .A2(G106gat), .A3(new_n503), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n839), .B(KEYINPUT113), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n840), .B1(new_n813), .B2(new_n814), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT53), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g641(.A1(new_n815), .A2(new_n839), .ZN(new_n843));
  OR2_X1    g642(.A1(new_n843), .A2(KEYINPUT53), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n838), .B2(new_n844), .ZN(G1339gat));
  NOR2_X1   g644(.A1(new_n684), .A2(new_n265), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n646), .A2(new_n642), .A3(new_n648), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n650), .A2(KEYINPUT54), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT54), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n655), .B1(new_n660), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT55), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n848), .A2(new_n853), .A3(new_n850), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n657), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n255), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n230), .B1(new_n238), .B2(new_n210), .ZN(new_n857));
  NAND4_X1  g656(.A1(new_n857), .A2(KEYINPUT114), .A3(G229gat), .A4(G233gat), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT114), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n247), .B2(new_n231), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n858), .B(new_n860), .C1(new_n251), .C2(new_n253), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n263), .A2(new_n856), .B1(new_n861), .B2(new_n260), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n855), .A2(new_n687), .A3(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n855), .A2(new_n265), .B1(new_n713), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n863), .B1(new_n864), .B2(new_n687), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n846), .B1(new_n865), .B2(new_n686), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n532), .A2(new_n534), .ZN(new_n867));
  NOR4_X1   g666(.A1(new_n866), .A2(new_n578), .A3(new_n695), .A4(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n868), .A2(new_n380), .A3(new_n265), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n866), .A2(new_n578), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n695), .A2(new_n531), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n736), .A3(new_n871), .ZN(new_n872));
  AND3_X1   g671(.A1(new_n872), .A2(KEYINPUT115), .A3(G113gat), .ZN(new_n873));
  AOI21_X1  g672(.A(KEYINPUT115), .B1(new_n872), .B2(G113gat), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n869), .B1(new_n873), .B2(new_n874), .ZN(G1340gat));
  NAND2_X1  g674(.A1(new_n870), .A2(new_n871), .ZN(new_n876));
  OAI21_X1  g675(.A(G120gat), .B1(new_n876), .B2(new_n665), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n868), .A2(new_n378), .A3(new_n713), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(G1341gat));
  NOR3_X1   g678(.A1(new_n876), .A2(new_n604), .A3(new_n686), .ZN(new_n880));
  XNOR2_X1  g679(.A(new_n880), .B(KEYINPUT116), .ZN(new_n881));
  NAND4_X1  g680(.A1(new_n870), .A2(new_n543), .A3(new_n532), .A4(new_n534), .ZN(new_n882));
  NOR3_X1   g681(.A1(new_n882), .A2(KEYINPUT117), .A3(new_n686), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n868), .B2(new_n622), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n883), .A2(G127gat), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n881), .A2(new_n886), .ZN(G1342gat));
  NOR3_X1   g686(.A1(new_n882), .A2(G134gat), .A3(new_n725), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT56), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g690(.A(G134gat), .B1(new_n876), .B2(new_n725), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n890), .A2(new_n891), .A3(new_n892), .ZN(G1343gat));
  NOR3_X1   g692(.A1(new_n695), .A2(new_n577), .A3(new_n578), .ZN(new_n894));
  INV_X1    g693(.A(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n854), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n853), .B1(new_n848), .B2(new_n850), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n711), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n716), .A2(KEYINPUT92), .ZN(new_n899));
  INV_X1    g698(.A(new_n268), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n861), .A2(new_n260), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n264), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n665), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n725), .B1(new_n901), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n622), .B1(new_n905), .B2(new_n863), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n583), .B1(new_n906), .B2(new_n846), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n895), .B1(new_n907), .B2(KEYINPUT57), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT118), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n898), .A2(new_n716), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n725), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n622), .B1(new_n912), .B2(new_n863), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n910), .B(new_n583), .C1(new_n913), .C2(new_n846), .ZN(new_n914));
  NAND4_X1  g713(.A1(new_n908), .A2(new_n909), .A3(new_n736), .A4(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n855), .B1(new_n267), .B2(new_n268), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n713), .A2(new_n862), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n687), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n863), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n686), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(new_n846), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n503), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI211_X1 g721(.A(new_n914), .B(new_n894), .C1(new_n922), .C2(new_n910), .ZN(new_n923));
  OAI21_X1  g722(.A(KEYINPUT118), .B1(new_n923), .B2(new_n269), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n915), .A2(new_n924), .A3(G141gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n866), .A2(new_n503), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n894), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n927), .A2(G141gat), .A3(new_n269), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n928), .A2(KEYINPUT58), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(new_n923), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n397), .B1(new_n931), .B2(new_n265), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT58), .B1(new_n932), .B2(new_n928), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n930), .A2(new_n933), .ZN(G1344gat));
  NOR2_X1   g733(.A1(new_n399), .A2(KEYINPUT59), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n923), .B2(new_n665), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(KEYINPUT119), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n736), .B1(new_n690), .B2(new_n685), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n910), .B(new_n583), .C1(new_n906), .C2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(KEYINPUT57), .B1(new_n866), .B2(new_n503), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n939), .A2(new_n713), .A3(new_n940), .A4(new_n894), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G148gat), .ZN(new_n942));
  XOR2_X1   g741(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n943));
  NAND2_X1  g742(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT119), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n945), .B(new_n935), .C1(new_n923), .C2(new_n665), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n937), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(new_n927), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(new_n399), .A3(new_n713), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1345gat));
  AND3_X1   g749(.A1(new_n931), .A2(G155gat), .A3(new_n622), .ZN(new_n951));
  AOI21_X1  g750(.A(G155gat), .B1(new_n948), .B2(new_n622), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1346gat));
  OAI21_X1  g752(.A(G162gat), .B1(new_n923), .B2(new_n725), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n725), .A2(G162gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n927), .B2(new_n955), .ZN(G1347gat));
  NOR4_X1   g755(.A1(new_n866), .A2(new_n692), .A3(new_n543), .A4(new_n867), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT121), .Z(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n259), .A3(new_n265), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n855), .A2(new_n265), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n687), .B1(new_n960), .B2(new_n917), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n686), .B1(new_n961), .B2(new_n919), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(new_n921), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n695), .A2(new_n578), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n796), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n963), .A2(new_n503), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n269), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n959), .A2(new_n967), .ZN(G1348gat));
  NOR3_X1   g767(.A1(new_n966), .A2(new_n298), .A3(new_n665), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n958), .A2(new_n713), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n969), .B1(new_n970), .B2(new_n298), .ZN(G1349gat));
  NAND4_X1  g770(.A1(new_n957), .A2(new_n313), .A3(new_n318), .A4(new_n622), .ZN(new_n972));
  OAI21_X1  g771(.A(G183gat), .B1(new_n966), .B2(new_n686), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT60), .ZN(new_n975));
  NOR2_X1   g774(.A1(new_n975), .A2(KEYINPUT122), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n974), .B(new_n976), .ZN(G1350gat));
  NAND3_X1  g776(.A1(new_n958), .A2(new_n288), .A3(new_n687), .ZN(new_n978));
  OAI21_X1  g777(.A(G190gat), .B1(new_n966), .B2(new_n725), .ZN(new_n979));
  XNOR2_X1  g778(.A(new_n979), .B(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1351gat));
  AOI21_X1  g780(.A(new_n692), .B1(new_n962), .B2(new_n921), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n543), .A2(new_n503), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(new_n798), .A3(new_n983), .ZN(new_n984));
  NOR3_X1   g783(.A1(new_n984), .A2(G197gat), .A3(new_n716), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT123), .ZN(new_n986));
  NOR2_X1   g785(.A1(new_n964), .A2(new_n577), .ZN(new_n987));
  XOR2_X1   g786(.A(new_n987), .B(KEYINPUT124), .Z(new_n988));
  NAND3_X1  g787(.A1(new_n939), .A2(new_n940), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(G197gat), .B1(new_n989), .B2(new_n269), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n986), .A2(new_n990), .ZN(G1352gat));
  NAND4_X1  g790(.A1(new_n939), .A2(new_n713), .A3(new_n940), .A4(new_n988), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n992), .A2(G204gat), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n982), .A2(new_n798), .A3(new_n983), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT125), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n665), .A2(G204gat), .ZN(new_n997));
  NAND4_X1  g796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n982), .A2(new_n798), .A3(new_n983), .A4(new_n997), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n999), .A2(KEYINPUT62), .ZN(new_n1000));
  OAI21_X1  g799(.A(KEYINPUT125), .B1(new_n999), .B2(KEYINPUT62), .ZN(new_n1001));
  NAND4_X1  g800(.A1(new_n993), .A2(new_n998), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g803(.A1(new_n992), .A2(G204gat), .B1(KEYINPUT62), .B2(new_n999), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n1005), .A2(KEYINPUT126), .A3(new_n1001), .A4(new_n998), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1353gat));
  OAI21_X1  g806(.A(G211gat), .B1(new_n989), .B2(new_n686), .ZN(new_n1008));
  OR2_X1    g807(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n984), .A2(G211gat), .A3(new_n686), .ZN(new_n1010));
  XNOR2_X1  g809(.A(new_n1010), .B(KEYINPUT127), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1008), .A2(KEYINPUT63), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1009), .A2(new_n1011), .A3(new_n1012), .ZN(G1354gat));
  NOR3_X1   g812(.A1(new_n989), .A2(new_n273), .A3(new_n725), .ZN(new_n1014));
  AOI21_X1  g813(.A(G218gat), .B1(new_n994), .B2(new_n687), .ZN(new_n1015));
  NOR2_X1   g814(.A1(new_n1014), .A2(new_n1015), .ZN(G1355gat));
endmodule


