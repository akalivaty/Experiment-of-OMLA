//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 0 0 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n838, new_n839, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n848, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963, new_n964;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT80), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g004(.A1(KEYINPUT80), .A2(G155gat), .A3(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OR2_X1    g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(G141gat), .B(G148gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT81), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(G113gat), .B(G120gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G127gat), .B(G134gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G120gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G113gat), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G120gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G127gat), .A2(G134gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G127gat), .A2(G134gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT70), .ZN(new_n226));
  NOR3_X1   g025(.A1(new_n226), .A2(KEYINPUT71), .A3(KEYINPUT1), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n215), .B1(KEYINPUT71), .B2(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n217), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G141gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(G148gat), .ZN(new_n232));
  INV_X1    g031(.A(G148gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G141gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n232), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND4_X1  g036(.A1(new_n237), .A2(KEYINPUT81), .A3(new_n208), .A4(new_n207), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n208), .A2(new_n203), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n239), .A2(new_n235), .A3(new_n236), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n213), .A2(new_n230), .A3(new_n238), .A4(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT83), .B(KEYINPUT4), .Z(new_n243));
  NOR2_X1   g042(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n202), .B1(new_n242), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(KEYINPUT4), .ZN(new_n246));
  OAI211_X1 g045(.A(new_n246), .B(KEYINPUT85), .C1(new_n241), .C2(new_n243), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n213), .A2(new_n238), .A3(new_n240), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(KEYINPUT3), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT3), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n213), .A2(new_n238), .A3(new_n251), .A4(new_n240), .ZN(new_n252));
  INV_X1    g051(.A(new_n230), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(KEYINPUT82), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT82), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n250), .A2(new_n256), .A3(new_n252), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n248), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(G225gat), .A2(G233gat), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(KEYINPUT84), .B(KEYINPUT5), .Z(new_n262));
  NOR3_X1   g061(.A1(new_n259), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n249), .B(new_n230), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n262), .B1(new_n264), .B2(new_n260), .ZN(new_n265));
  INV_X1    g064(.A(new_n241), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(new_n243), .ZN(new_n267));
  AOI211_X1 g066(.A(new_n261), .B(new_n267), .C1(KEYINPUT4), .C2(new_n266), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(new_n258), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n263), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT0), .B(G57gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n271), .B(G85gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(G1gat), .B(G29gat), .ZN(new_n273));
  XOR2_X1   g072(.A(new_n272), .B(new_n273), .Z(new_n274));
  AOI21_X1  g073(.A(KEYINPUT6), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n276), .B1(new_n263), .B2(new_n269), .ZN(new_n277));
  OR2_X1    g076(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n275), .A2(new_n277), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G183gat), .ZN(new_n281));
  INV_X1    g080(.A(G190gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G183gat), .A2(G190gat), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT24), .A3(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n285), .B1(KEYINPUT24), .B2(new_n284), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT23), .ZN(new_n287));
  INV_X1    g086(.A(G169gat), .ZN(new_n288));
  INV_X1    g087(.A(G176gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT67), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT67), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n291), .B1(G169gat), .B2(G176gat), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n287), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n296), .A2(G169gat), .A3(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT68), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n286), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  OAI21_X1  g100(.A(KEYINPUT68), .B1(new_n293), .B2(new_n298), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n287), .B1(G169gat), .B2(G176gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n302), .A4(new_n303), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(KEYINPUT23), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n305), .A2(new_n303), .A3(new_n294), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT64), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n284), .A2(KEYINPUT24), .ZN(new_n308));
  AND2_X1   g107(.A1(G183gat), .A2(G190gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n308), .B1(new_n311), .B2(KEYINPUT24), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT64), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n305), .A2(new_n303), .A3(new_n313), .A4(new_n294), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n307), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT65), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n315), .A2(new_n319), .A3(new_n316), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n290), .A2(new_n292), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(new_n322), .B(new_n294), .C1(new_n324), .C2(KEYINPUT26), .ZN(new_n325));
  XOR2_X1   g124(.A(KEYINPUT27), .B(G183gat), .Z(new_n326));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OR2_X1    g127(.A1(new_n281), .A2(KEYINPUT27), .ZN(new_n329));
  AOI21_X1  g128(.A(G190gat), .B1(new_n329), .B2(KEYINPUT69), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT28), .B1(new_n328), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT28), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n326), .A2(new_n332), .A3(G190gat), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n325), .B(new_n284), .C1(new_n331), .C2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n321), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(G226gat), .A2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT78), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT78), .ZN(new_n339));
  AOI211_X1 g138(.A(new_n339), .B(new_n336), .C1(new_n321), .C2(new_n334), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  XNOR2_X1  g140(.A(G211gat), .B(G218gat), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n342), .B(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G197gat), .B(G204gat), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n346));
  OR2_X1    g145(.A1(new_n346), .A2(KEYINPUT22), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(KEYINPUT22), .ZN(new_n348));
  INV_X1    g147(.A(G211gat), .ZN(new_n349));
  INV_X1    g148(.A(G218gat), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n347), .B(new_n348), .C1(new_n349), .C2(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(new_n345), .A3(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(new_n342), .B(KEYINPUT76), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n351), .A2(new_n345), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT77), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n335), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n334), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT29), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n341), .B(new_n357), .C1(new_n361), .C2(new_n337), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT29), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n335), .A2(new_n363), .A3(new_n336), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n359), .A2(new_n360), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n356), .B(new_n364), .C1(new_n365), .C2(new_n336), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G64gat), .B(G92gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n368), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n369), .B(KEYINPUT79), .ZN(new_n370));
  INV_X1    g169(.A(G8gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n372), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n362), .A2(new_n366), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n373), .A2(KEYINPUT30), .A3(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT30), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n367), .A2(new_n377), .A3(new_n372), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n280), .A2(new_n379), .ZN(new_n380));
  XNOR2_X1  g179(.A(G78gat), .B(G106gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n381), .B(G22gat), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT86), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n352), .A2(new_n384), .A3(new_n355), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n353), .A2(new_n354), .A3(KEYINPUT86), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(new_n363), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT87), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g188(.A1(new_n385), .A2(KEYINPUT87), .A3(new_n363), .A4(new_n386), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(new_n251), .A3(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(new_n249), .ZN(new_n392));
  INV_X1    g191(.A(G228gat), .ZN(new_n393));
  INV_X1    g192(.A(G233gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n252), .A2(new_n363), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n357), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n392), .A2(new_n396), .A3(new_n398), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT31), .B(G50gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n251), .B1(new_n357), .B2(KEYINPUT29), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n402), .A2(new_n249), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(new_n398), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n395), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n399), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n399), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n383), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n399), .A2(new_n405), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n400), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n399), .A2(new_n401), .A3(new_n405), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(new_n382), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n408), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n335), .A2(new_n253), .ZN(new_n414));
  INV_X1    g213(.A(G227gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n415), .A2(new_n394), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n321), .A2(new_n230), .A3(new_n334), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT73), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT34), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT74), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT74), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n421), .A2(new_n425), .A3(new_n422), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n414), .A2(new_n418), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n416), .ZN(new_n429));
  XNOR2_X1  g228(.A(G15gat), .B(G43gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(G71gat), .ZN(new_n431));
  XNOR2_X1  g230(.A(new_n431), .B(G99gat), .ZN(new_n432));
  OR2_X1    g231(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n432), .A2(KEYINPUT72), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(KEYINPUT33), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n429), .A2(KEYINPUT32), .A3(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT32), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n428), .A2(new_n416), .B1(new_n437), .B2(KEYINPUT33), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n438), .B2(new_n432), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n419), .A2(new_n420), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OAI221_X1 g240(.A(new_n436), .B1(new_n420), .B2(new_n419), .C1(new_n432), .C2(new_n438), .ZN(new_n442));
  AND3_X1   g241(.A1(new_n427), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI22_X1  g242(.A1(new_n441), .A2(new_n442), .B1(new_n424), .B2(new_n426), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n413), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT35), .B1(new_n380), .B2(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n408), .A2(new_n412), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n442), .ZN(new_n448));
  INV_X1    g247(.A(new_n427), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n427), .A2(new_n441), .A3(new_n442), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n447), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT35), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n452), .A2(new_n453), .A3(new_n280), .A4(new_n379), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n380), .A2(new_n413), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT39), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n245), .A2(new_n247), .B1(new_n255), .B2(new_n257), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n458), .A2(KEYINPUT88), .A3(new_n260), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT88), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n460), .B1(new_n259), .B2(new_n261), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n457), .B1(new_n459), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n462), .A2(KEYINPUT89), .A3(new_n274), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT88), .B1(new_n458), .B2(new_n260), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n259), .A2(new_n460), .A3(new_n261), .ZN(new_n466));
  AOI21_X1  g265(.A(KEYINPUT39), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n464), .B1(new_n467), .B2(new_n276), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n459), .A2(new_n461), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n457), .B1(new_n264), .B2(new_n260), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n463), .A2(new_n468), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n379), .B1(new_n471), .B2(KEYINPUT40), .ZN(new_n472));
  OR2_X1    g271(.A1(new_n471), .A2(KEYINPUT40), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT90), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n472), .A2(new_n473), .A3(new_n474), .A4(new_n277), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n469), .A2(new_n470), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT89), .B1(new_n462), .B2(new_n274), .ZN(new_n477));
  NOR3_X1   g276(.A1(new_n467), .A2(new_n464), .A3(new_n276), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT40), .B(new_n476), .C1(new_n477), .C2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n479), .A2(new_n277), .A3(new_n378), .A4(new_n376), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n471), .A2(KEYINPUT40), .ZN(new_n481));
  OAI21_X1  g280(.A(KEYINPUT90), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(new_n280), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT37), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n372), .B1(new_n367), .B2(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n485), .B1(new_n484), .B2(new_n367), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT38), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n341), .B1(new_n361), .B2(new_n337), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(new_n356), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n364), .B1(new_n365), .B2(new_n336), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n484), .B1(new_n490), .B2(new_n357), .ZN(new_n491));
  AOI21_X1  g290(.A(KEYINPUT38), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n485), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g292(.A1(new_n483), .A2(new_n373), .A3(new_n487), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n475), .A2(new_n482), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n456), .B1(new_n495), .B2(new_n413), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n450), .A2(new_n451), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(KEYINPUT36), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT36), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n497), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n455), .B1(new_n496), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(G230gat), .A2(G233gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G99gat), .A2(G106gat), .ZN(new_n506));
  INV_X1    g305(.A(G85gat), .ZN(new_n507));
  INV_X1    g306(.A(G92gat), .ZN(new_n508));
  AOI22_X1  g307(.A1(KEYINPUT8), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT7), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n507), .B2(new_n508), .ZN(new_n511));
  NAND3_X1  g310(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  XNOR2_X1  g312(.A(G99gat), .B(G106gat), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT93), .ZN(new_n517));
  INV_X1    g316(.A(G64gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G57gat), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT92), .B(G57gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n520), .B1(new_n521), .B2(G64gat), .ZN(new_n522));
  NOR2_X1   g321(.A1(G71gat), .A2(G78gat), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n523), .A2(KEYINPUT9), .ZN(new_n524));
  NAND2_X1  g323(.A1(G71gat), .A2(G78gat), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n517), .B1(new_n522), .B2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(KEYINPUT92), .A2(G57gat), .ZN(new_n529));
  OAI21_X1  g328(.A(G64gat), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n519), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(new_n525), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n531), .A2(KEYINPUT93), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n527), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n523), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n525), .ZN(new_n536));
  XOR2_X1   g335(.A(G57gat), .B(G64gat), .Z(new_n537));
  AOI21_X1  g336(.A(new_n536), .B1(new_n537), .B2(KEYINPUT9), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(KEYINPUT94), .B1(new_n534), .B2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT94), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n541), .B(new_n538), .C1(new_n527), .C2(new_n533), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n516), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AOI221_X4 g342(.A(new_n517), .B1(new_n524), .B2(new_n525), .C1(new_n530), .C2(new_n519), .ZN(new_n544));
  AOI21_X1  g343(.A(KEYINPUT93), .B1(new_n531), .B2(new_n532), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n539), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n515), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT10), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT10), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n546), .A2(new_n541), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT94), .A3(new_n539), .ZN(new_n551));
  AOI211_X1 g350(.A(new_n549), .B(new_n516), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(KEYINPUT100), .B1(new_n548), .B2(new_n552), .ZN(new_n553));
  AOI21_X1  g352(.A(new_n515), .B1(new_n550), .B2(new_n551), .ZN(new_n554));
  INV_X1    g353(.A(new_n547), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n549), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT100), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n550), .A2(new_n551), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT10), .A3(new_n515), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n556), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n505), .B1(new_n553), .B2(new_n560), .ZN(new_n561));
  NOR3_X1   g360(.A1(new_n554), .A2(new_n504), .A3(new_n555), .ZN(new_n562));
  XNOR2_X1  g361(.A(G120gat), .B(G148gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(new_n289), .ZN(new_n564));
  INV_X1    g363(.A(G204gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NOR3_X1   g365(.A1(new_n561), .A2(new_n562), .A3(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n504), .B(KEYINPUT101), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n556), .B2(new_n559), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n570), .A2(new_n562), .ZN(new_n571));
  INV_X1    g370(.A(new_n566), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n567), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n503), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT14), .ZN(new_n579));
  INV_X1    g378(.A(G29gat), .ZN(new_n580));
  INV_X1    g379(.A(G36gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT91), .ZN(new_n583));
  OAI21_X1  g382(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT91), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(new_n579), .A3(new_n580), .A4(new_n581), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n580), .A2(new_n581), .ZN(new_n588));
  INV_X1    g387(.A(G50gat), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(G43gat), .ZN(new_n590));
  INV_X1    g389(.A(G43gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n591), .A2(G50gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT15), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n588), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n590), .A2(new_n592), .A3(KEYINPUT15), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n587), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n596), .ZN(new_n598));
  AND2_X1   g397(.A1(new_n582), .A2(new_n584), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n588), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(KEYINPUT17), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT17), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n597), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n578), .B1(new_n605), .B2(new_n516), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n515), .A2(new_n601), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n282), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n597), .A2(new_n603), .A3(new_n600), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n603), .B1(new_n597), .B2(new_n600), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n516), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n611), .A2(new_n282), .A3(new_n577), .A4(new_n607), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n350), .B1(new_n608), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n611), .A2(new_n577), .A3(new_n607), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G190gat), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n616), .A2(G218gat), .A3(new_n612), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(KEYINPUT99), .A3(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(KEYINPUT98), .A3(new_n617), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(G134gat), .B(G162gat), .ZN(new_n622));
  XOR2_X1   g421(.A(new_n622), .B(KEYINPUT97), .Z(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n620), .ZN(new_n625));
  NAND4_X1  g424(.A1(new_n614), .A2(KEYINPUT98), .A3(new_n625), .A4(new_n617), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n621), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n624), .B1(new_n621), .B2(new_n626), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n618), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n621), .A2(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n623), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n621), .A2(new_n624), .A3(new_n626), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n631), .A2(KEYINPUT99), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G15gat), .B(G22gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n636), .A2(G1gat), .ZN(new_n637));
  INV_X1    g436(.A(G1gat), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT16), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n637), .B1(new_n639), .B2(new_n636), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(new_n371), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n641), .B1(new_n558), .B2(KEYINPUT21), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(KEYINPUT21), .B2(new_n558), .ZN(new_n643));
  XNOR2_X1  g442(.A(G183gat), .B(G211gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n641), .ZN(new_n645));
  OR3_X1    g444(.A1(new_n558), .A2(new_n645), .A3(KEYINPUT21), .ZN(new_n646));
  AND3_X1   g445(.A1(new_n643), .A2(new_n644), .A3(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n644), .B1(new_n643), .B2(new_n646), .ZN(new_n648));
  XOR2_X1   g447(.A(G127gat), .B(G155gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT20), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n647), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(G231gat), .A2(G233gat), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(KEYINPUT19), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT95), .B(KEYINPUT96), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n650), .B1(new_n647), .B2(new_n648), .ZN(new_n656));
  AND3_X1   g455(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n655), .B1(new_n651), .B2(new_n656), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n635), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n605), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n641), .A2(new_n601), .ZN(new_n662));
  NAND2_X1  g461(.A1(G229gat), .A2(G233gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT18), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n641), .B(new_n601), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n663), .B(KEYINPUT13), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n661), .A2(KEYINPUT18), .A3(new_n662), .A4(new_n663), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT11), .B(G169gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G197gat), .ZN(new_n673));
  XOR2_X1   g472(.A(G113gat), .B(G141gat), .Z(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT12), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n671), .B(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n660), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n576), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n679), .A2(new_n280), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(new_n638), .ZN(G1324gat));
  NOR2_X1   g480(.A1(new_n679), .A2(new_n379), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n682), .A2(new_n371), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT103), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n685));
  AOI21_X1  g484(.A(KEYINPUT42), .B1(new_n682), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n679), .A2(new_n379), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AND2_X1   g488(.A1(new_n686), .A2(new_n688), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n684), .B1(new_n689), .B2(new_n690), .ZN(G1325gat));
  NOR3_X1   g490(.A1(new_n679), .A2(G15gat), .A3(new_n498), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n502), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n499), .A2(KEYINPUT104), .A3(new_n501), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n576), .A2(new_n678), .A3(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n692), .B1(G15gat), .B2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT105), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n679), .A2(new_n413), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  NOR3_X1   g501(.A1(new_n659), .A2(new_n574), .A3(new_n677), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n503), .A2(new_n634), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n580), .A3(new_n483), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n503), .A2(new_n634), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT106), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n446), .A2(new_n709), .A3(new_n454), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n446), .B2(new_n454), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n712), .B1(new_n496), .B2(new_n696), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT44), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n634), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n708), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n716), .A2(new_n703), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n280), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n706), .A2(new_n718), .ZN(G1328gat));
  INV_X1    g518(.A(new_n379), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n581), .A3(new_n720), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT46), .Z(new_n722));
  NAND3_X1  g521(.A1(new_n716), .A2(new_n720), .A3(new_n703), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(new_n581), .ZN(G1329gat));
  NAND3_X1  g524(.A1(new_n716), .A2(new_n696), .A3(new_n703), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n498), .A2(G43gat), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n726), .A2(G43gat), .B1(new_n704), .B2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT48), .ZN(new_n731));
  OAI21_X1  g530(.A(G50gat), .B1(new_n717), .B2(new_n413), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n704), .A2(new_n589), .A3(new_n447), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n730), .B(new_n731), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(KEYINPUT107), .A2(KEYINPUT48), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n730), .A2(new_n731), .ZN(new_n736));
  AND4_X1   g535(.A1(new_n735), .A2(new_n732), .A3(new_n736), .A4(new_n733), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n734), .A2(new_n737), .ZN(G1331gat));
  AND4_X1   g537(.A1(new_n659), .A2(new_n713), .A3(new_n635), .A4(new_n677), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(new_n574), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n280), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(new_n521), .ZN(G1332gat));
  NOR2_X1   g541(.A1(new_n740), .A2(new_n379), .ZN(new_n743));
  NOR2_X1   g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  AND2_X1   g543(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n743), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n746), .B1(new_n743), .B2(new_n744), .ZN(G1333gat));
  AND2_X1   g546(.A1(new_n739), .A2(new_n574), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n696), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n740), .A2(G71gat), .ZN(new_n750));
  AOI22_X1  g549(.A1(new_n749), .A2(G71gat), .B1(new_n750), .B2(new_n497), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g551(.A1(new_n748), .A2(new_n447), .ZN(new_n753));
  XNOR2_X1  g552(.A(new_n753), .B(G78gat), .ZN(G1335gat));
  INV_X1    g553(.A(new_n677), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n659), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n713), .A2(new_n634), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(KEYINPUT51), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT51), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n713), .A2(new_n759), .A3(new_n634), .A4(new_n756), .ZN(new_n760));
  AND2_X1   g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n761), .A2(new_n574), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(new_n507), .A3(new_n483), .ZN(new_n763));
  INV_X1    g562(.A(new_n756), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n764), .B1(new_n708), .B2(new_n715), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n765), .A2(new_n483), .A3(new_n574), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT108), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n763), .B1(new_n767), .B2(new_n507), .ZN(G1336gat));
  NAND4_X1  g567(.A1(new_n765), .A2(G92gat), .A3(new_n574), .A4(new_n720), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n758), .A2(new_n574), .A3(new_n720), .A4(new_n760), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n508), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n769), .B(new_n771), .C1(KEYINPUT109), .C2(KEYINPUT52), .ZN(new_n772));
  NAND2_X1  g571(.A1(KEYINPUT109), .A2(KEYINPUT52), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1337gat));
  INV_X1    g573(.A(G99gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n762), .A2(new_n775), .A3(new_n497), .ZN(new_n776));
  AND3_X1   g575(.A1(new_n713), .A2(new_n714), .A3(new_n634), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n714), .B1(new_n503), .B2(new_n634), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n574), .B(new_n756), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n694), .A2(new_n695), .ZN(new_n780));
  OAI21_X1  g579(.A(G99gat), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n776), .A2(new_n781), .ZN(G1338gat));
  OAI21_X1  g581(.A(G106gat), .B1(new_n779), .B2(new_n413), .ZN(new_n783));
  AOI21_X1  g582(.A(KEYINPUT53), .B1(new_n783), .B2(KEYINPUT110), .ZN(new_n784));
  INV_X1    g583(.A(G106gat), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n761), .A2(new_n785), .A3(new_n574), .A4(new_n447), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n783), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n786), .B(new_n783), .C1(KEYINPUT110), .C2(KEYINPUT53), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n788), .A2(new_n789), .ZN(G1339gat));
  INV_X1    g589(.A(new_n659), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT54), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n572), .B1(new_n570), .B2(new_n792), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n556), .A2(new_n559), .ZN(new_n794));
  OAI21_X1  g593(.A(KEYINPUT54), .B1(new_n794), .B2(new_n568), .ZN(new_n795));
  OAI211_X1 g594(.A(KEYINPUT55), .B(new_n793), .C1(new_n561), .C2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n548), .A2(KEYINPUT100), .A3(new_n552), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n557), .B1(new_n556), .B2(new_n559), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n504), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n548), .A2(new_n552), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n792), .B1(new_n801), .B2(new_n569), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT111), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT55), .A4(new_n793), .ZN(new_n805));
  INV_X1    g604(.A(new_n567), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n797), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(KEYINPUT112), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT112), .ZN(new_n809));
  NAND4_X1  g608(.A1(new_n797), .A2(new_n805), .A3(new_n809), .A4(new_n806), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n793), .B1(new_n561), .B2(new_n795), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT55), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n808), .A2(new_n755), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n666), .A2(new_n669), .A3(new_n676), .A4(new_n670), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n667), .A2(new_n668), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n663), .B1(new_n661), .B2(new_n662), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n675), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n574), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n634), .B1(new_n814), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n813), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n823), .B1(new_n807), .B2(KEYINPUT112), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n634), .A3(new_n820), .A4(new_n810), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n791), .B1(new_n822), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n635), .A2(new_n575), .A3(new_n659), .A4(new_n677), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n280), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n829), .A2(new_n452), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n830), .A2(new_n379), .ZN(new_n831));
  OAI21_X1  g630(.A(G113gat), .B1(new_n831), .B2(new_n677), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n755), .A2(new_n220), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT113), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n832), .B1(new_n831), .B2(new_n834), .ZN(G1340gat));
  NOR2_X1   g634(.A1(new_n831), .A2(new_n575), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(new_n218), .ZN(G1341gat));
  INV_X1    g636(.A(G127gat), .ZN(new_n838));
  AOI21_X1  g637(.A(KEYINPUT114), .B1(new_n838), .B2(KEYINPUT115), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n839), .B1(KEYINPUT114), .B2(new_n838), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n831), .A2(new_n791), .ZN(new_n841));
  MUX2_X1   g640(.A(new_n839), .B(new_n840), .S(new_n841), .Z(G1342gat));
  NAND2_X1  g641(.A1(new_n634), .A2(new_n379), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT116), .Z(new_n844));
  NOR2_X1   g643(.A1(new_n844), .A2(G134gat), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n845), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n846), .B(KEYINPUT56), .Z(new_n847));
  OAI21_X1  g646(.A(G134gat), .B1(new_n831), .B2(new_n635), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n847), .A2(new_n848), .ZN(G1343gat));
  NAND3_X1  g648(.A1(new_n829), .A2(new_n447), .A3(new_n780), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n720), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n755), .A2(new_n231), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n853), .A2(new_n854), .ZN(new_n857));
  OR3_X1    g656(.A1(new_n852), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT58), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n696), .A2(new_n280), .A3(new_n720), .ZN(new_n860));
  AND3_X1   g659(.A1(new_n808), .A2(new_n810), .A3(new_n813), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n819), .B1(new_n629), .B2(new_n633), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n755), .A2(new_n813), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n821), .B1(new_n807), .B2(new_n863), .ZN(new_n864));
  AOI22_X1  g663(.A1(new_n861), .A2(new_n862), .B1(new_n635), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n828), .B1(new_n865), .B2(new_n659), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT57), .A4(new_n447), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n633), .A3(new_n629), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n659), .B1(new_n825), .B2(new_n869), .ZN(new_n870));
  NOR4_X1   g669(.A1(new_n791), .A2(new_n634), .A3(new_n574), .A4(new_n755), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT57), .B(new_n447), .C1(new_n870), .C2(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT117), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n827), .A2(new_n828), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n875), .B2(new_n447), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n860), .B1(new_n874), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g676(.A(G141gat), .B1(new_n877), .B2(new_n677), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n858), .A2(new_n859), .A3(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n852), .A2(new_n856), .A3(new_n857), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n413), .B1(new_n827), .B2(new_n828), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n868), .B(new_n873), .C1(KEYINPUT57), .C2(new_n881), .ZN(new_n882));
  AND3_X1   g681(.A1(new_n882), .A2(KEYINPUT118), .A3(new_n860), .ZN(new_n883));
  AOI21_X1  g682(.A(KEYINPUT118), .B1(new_n882), .B2(new_n860), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n755), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n880), .B1(new_n885), .B2(G141gat), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n886), .A2(KEYINPUT120), .A3(new_n859), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT120), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n877), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n882), .A2(KEYINPUT118), .A3(new_n860), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n677), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n858), .B1(new_n892), .B2(new_n231), .ZN(new_n893));
  AOI21_X1  g692(.A(new_n888), .B1(new_n893), .B2(KEYINPUT58), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n879), .B1(new_n887), .B2(new_n894), .ZN(G1344gat));
  NOR2_X1   g694(.A1(new_n883), .A2(new_n884), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n575), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  INV_X1    g697(.A(new_n866), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n898), .B1(new_n899), .B2(new_n413), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n881), .A2(KEYINPUT57), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(new_n574), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n860), .A2(KEYINPUT59), .ZN(new_n904));
  OAI22_X1  g703(.A1(new_n897), .A2(KEYINPUT59), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(G148gat), .B1(new_n851), .B2(new_n574), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n905), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n906), .ZN(G1345gat));
  AOI21_X1  g706(.A(G155gat), .B1(new_n851), .B2(new_n659), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n896), .A2(new_n791), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n909), .B2(G155gat), .ZN(G1346gat));
  OAI21_X1  g709(.A(G162gat), .B1(new_n896), .B2(new_n635), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n850), .A2(G162gat), .A3(new_n844), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT121), .Z(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1347gat));
  AOI21_X1  g713(.A(new_n445), .B1(new_n827), .B2(new_n828), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n483), .A2(new_n379), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n677), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(new_n288), .ZN(G1348gat));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n575), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(new_n289), .ZN(G1349gat));
  NOR2_X1   g720(.A1(new_n917), .A2(new_n791), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(new_n326), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n923), .B1(G183gat), .B2(new_n922), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT122), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(KEYINPUT60), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n924), .B(new_n926), .ZN(G1350gat));
  NAND3_X1  g726(.A1(new_n915), .A2(new_n634), .A3(new_n916), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT123), .B1(new_n928), .B2(G190gat), .ZN(new_n929));
  INV_X1    g728(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n928), .A2(KEYINPUT123), .A3(G190gat), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n930), .A2(KEYINPUT124), .A3(new_n931), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(KEYINPUT61), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT61), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n932), .A2(new_n933), .A3(new_n937), .ZN(new_n938));
  OAI211_X1 g737(.A(new_n936), .B(new_n938), .C1(G190gat), .C2(new_n928), .ZN(G1351gat));
  NAND2_X1  g738(.A1(new_n780), .A2(new_n916), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n940), .B1(new_n900), .B2(new_n901), .ZN(new_n941));
  INV_X1    g740(.A(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n677), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n881), .A2(new_n780), .A3(new_n916), .ZN(new_n944));
  INV_X1    g743(.A(new_n944), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n945), .A2(G197gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n943), .B1(new_n677), .B2(new_n946), .ZN(G1352gat));
  NAND3_X1  g746(.A1(new_n944), .A2(new_n565), .A3(new_n574), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT62), .Z(new_n949));
  OAI21_X1  g748(.A(G204gat), .B1(new_n903), .B2(new_n940), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n949), .A2(new_n950), .ZN(G1353gat));
  AOI21_X1  g750(.A(new_n349), .B1(new_n941), .B2(new_n659), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n952), .A2(KEYINPUT63), .ZN(new_n953));
  OR2_X1    g752(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n955));
  OR3_X1    g754(.A1(new_n952), .A2(new_n955), .A3(KEYINPUT63), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n953), .A2(KEYINPUT125), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n955), .B1(new_n952), .B2(KEYINPUT63), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n954), .A2(new_n956), .A3(new_n957), .A4(new_n958), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n944), .A2(new_n349), .A3(new_n659), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n944), .B2(new_n634), .ZN(new_n962));
  XOR2_X1   g761(.A(new_n962), .B(KEYINPUT127), .Z(new_n963));
  NOR3_X1   g762(.A1(new_n942), .A2(new_n350), .A3(new_n635), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n963), .A2(new_n964), .ZN(G1355gat));
endmodule


