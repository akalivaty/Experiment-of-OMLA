

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U555 ( .A(n706), .B(n705), .ZN(n712) );
  NOR2_X1 U556 ( .A1(G2104), .A2(n532), .ZN(n893) );
  NOR2_X2 U557 ( .A1(n717), .A2(n716), .ZN(n718) );
  INV_X1 U558 ( .A(G2105), .ZN(n532) );
  NOR2_X2 U559 ( .A1(n755), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U560 ( .A1(G2104), .A2(G2105), .ZN(n531) );
  OR2_X1 U561 ( .A1(n618), .A2(n617), .ZN(n619) );
  INV_X1 U562 ( .A(KEYINPUT23), .ZN(n527) );
  XOR2_X1 U563 ( .A(KEYINPUT71), .B(n613), .Z(n521) );
  AND2_X1 U564 ( .A1(G1976), .A2(G288), .ZN(n522) );
  AND2_X1 U565 ( .A1(n937), .A2(n815), .ZN(n523) );
  AND2_X1 U566 ( .A1(n768), .A2(n767), .ZN(n524) );
  OR2_X1 U567 ( .A1(n765), .A2(n757), .ZN(n525) );
  AND2_X1 U568 ( .A1(n758), .A2(n525), .ZN(n526) );
  INV_X1 U569 ( .A(KEYINPUT27), .ZN(n701) );
  INV_X1 U570 ( .A(KEYINPUT90), .ZN(n713) );
  XNOR2_X1 U571 ( .A(n713), .B(KEYINPUT28), .ZN(n714) );
  XNOR2_X1 U572 ( .A(n715), .B(n714), .ZN(n716) );
  NAND2_X1 U573 ( .A1(n689), .A2(n772), .ZN(n723) );
  NAND2_X1 U574 ( .A1(G8), .A2(n723), .ZN(n765) );
  NOR2_X1 U575 ( .A1(n802), .A2(n523), .ZN(n803) );
  NOR2_X1 U576 ( .A1(G651), .A2(n642), .ZN(n654) );
  AND2_X2 U577 ( .A1(n532), .A2(G2104), .ZN(n886) );
  XNOR2_X1 U578 ( .A(n528), .B(n527), .ZN(n530) );
  NAND2_X1 U579 ( .A1(G101), .A2(n886), .ZN(n528) );
  AND2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n892) );
  NAND2_X1 U581 ( .A1(n892), .A2(G113), .ZN(n529) );
  NAND2_X1 U582 ( .A1(n530), .A2(n529), .ZN(n536) );
  XOR2_X2 U583 ( .A(KEYINPUT17), .B(n531), .Z(n888) );
  NAND2_X1 U584 ( .A1(G137), .A2(n888), .ZN(n534) );
  NAND2_X1 U585 ( .A1(G125), .A2(n893), .ZN(n533) );
  NAND2_X1 U586 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U587 ( .A1(n536), .A2(n535), .ZN(G160) );
  XNOR2_X1 U588 ( .A(KEYINPUT74), .B(KEYINPUT6), .ZN(n541) );
  INV_X1 U589 ( .A(G651), .ZN(n543) );
  NOR2_X1 U590 ( .A1(G543), .A2(n543), .ZN(n537) );
  XOR2_X2 U591 ( .A(KEYINPUT1), .B(n537), .Z(n653) );
  NAND2_X1 U592 ( .A1(G63), .A2(n653), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT0), .B(G543), .Z(n642) );
  NAND2_X1 U594 ( .A1(G51), .A2(n654), .ZN(n538) );
  NAND2_X1 U595 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U596 ( .A(n541), .B(n540), .ZN(n549) );
  NOR2_X1 U597 ( .A1(G651), .A2(G543), .ZN(n658) );
  NAND2_X1 U598 ( .A1(n658), .A2(G89), .ZN(n542) );
  XNOR2_X1 U599 ( .A(n542), .B(KEYINPUT4), .ZN(n545) );
  NOR2_X1 U600 ( .A1(n642), .A2(n543), .ZN(n657) );
  NAND2_X1 U601 ( .A1(G76), .A2(n657), .ZN(n544) );
  NAND2_X1 U602 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U603 ( .A(KEYINPUT5), .B(n546), .ZN(n547) );
  XNOR2_X1 U604 ( .A(KEYINPUT73), .B(n547), .ZN(n548) );
  NOR2_X1 U605 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U606 ( .A(KEYINPUT7), .B(n550), .Z(G168) );
  XOR2_X1 U607 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U608 ( .A1(G138), .A2(n888), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G102), .A2(n886), .ZN(n551) );
  NAND2_X1 U610 ( .A1(n552), .A2(n551), .ZN(n556) );
  NAND2_X1 U611 ( .A1(G114), .A2(n892), .ZN(n554) );
  NAND2_X1 U612 ( .A1(G126), .A2(n893), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U614 ( .A1(n556), .A2(n555), .ZN(G164) );
  NAND2_X1 U615 ( .A1(G72), .A2(n657), .ZN(n558) );
  NAND2_X1 U616 ( .A1(G85), .A2(n658), .ZN(n557) );
  NAND2_X1 U617 ( .A1(n558), .A2(n557), .ZN(n562) );
  NAND2_X1 U618 ( .A1(G60), .A2(n653), .ZN(n560) );
  NAND2_X1 U619 ( .A1(G47), .A2(n654), .ZN(n559) );
  NAND2_X1 U620 ( .A1(n560), .A2(n559), .ZN(n561) );
  OR2_X1 U621 ( .A1(n562), .A2(n561), .ZN(G290) );
  XNOR2_X1 U622 ( .A(G2427), .B(KEYINPUT97), .ZN(n572) );
  XOR2_X1 U623 ( .A(G2443), .B(G2438), .Z(n564) );
  XNOR2_X1 U624 ( .A(G2430), .B(G2454), .ZN(n563) );
  XNOR2_X1 U625 ( .A(n564), .B(n563), .ZN(n568) );
  XOR2_X1 U626 ( .A(KEYINPUT96), .B(G2435), .Z(n566) );
  XNOR2_X1 U627 ( .A(G1348), .B(G1341), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n566), .B(n565), .ZN(n567) );
  XOR2_X1 U629 ( .A(n568), .B(n567), .Z(n570) );
  XNOR2_X1 U630 ( .A(G2451), .B(G2446), .ZN(n569) );
  XNOR2_X1 U631 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U632 ( .A(n572), .B(n571), .ZN(n573) );
  AND2_X1 U633 ( .A1(n573), .A2(G14), .ZN(G401) );
  NAND2_X1 U634 ( .A1(G64), .A2(n653), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G52), .A2(n654), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U637 ( .A(KEYINPUT64), .B(n576), .ZN(n581) );
  NAND2_X1 U638 ( .A1(G77), .A2(n657), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G90), .A2(n658), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n579) );
  XOR2_X1 U641 ( .A(KEYINPUT9), .B(n579), .Z(n580) );
  NOR2_X1 U642 ( .A1(n581), .A2(n580), .ZN(G171) );
  INV_X1 U643 ( .A(G57), .ZN(G237) );
  NAND2_X1 U644 ( .A1(G75), .A2(n657), .ZN(n582) );
  XOR2_X1 U645 ( .A(KEYINPUT80), .B(n582), .Z(n589) );
  NAND2_X1 U646 ( .A1(G62), .A2(n653), .ZN(n584) );
  NAND2_X1 U647 ( .A1(G50), .A2(n654), .ZN(n583) );
  NAND2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U649 ( .A(n585), .B(KEYINPUT79), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G88), .A2(n658), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U652 ( .A1(n589), .A2(n588), .ZN(G166) );
  NAND2_X1 U653 ( .A1(n654), .A2(G53), .ZN(n596) );
  NAND2_X1 U654 ( .A1(G78), .A2(n657), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G65), .A2(n653), .ZN(n590) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n594) );
  NAND2_X1 U657 ( .A1(n658), .A2(G91), .ZN(n592) );
  XOR2_X1 U658 ( .A(KEYINPUT66), .B(n592), .Z(n593) );
  NOR2_X1 U659 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U660 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(KEYINPUT67), .B(n597), .Z(G299) );
  NAND2_X1 U662 ( .A1(G94), .A2(G452), .ZN(n598) );
  XNOR2_X1 U663 ( .A(n598), .B(KEYINPUT65), .ZN(G173) );
  NAND2_X1 U664 ( .A1(G7), .A2(G661), .ZN(n599) );
  XNOR2_X1 U665 ( .A(n599), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U666 ( .A(KEYINPUT68), .B(KEYINPUT11), .Z(n601) );
  INV_X1 U667 ( .A(G223), .ZN(n820) );
  NAND2_X1 U668 ( .A1(G567), .A2(n820), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n601), .B(n600), .ZN(G234) );
  NAND2_X1 U670 ( .A1(n653), .A2(G56), .ZN(n602) );
  XOR2_X1 U671 ( .A(KEYINPUT14), .B(n602), .Z(n609) );
  NAND2_X1 U672 ( .A1(n657), .A2(G68), .ZN(n603) );
  XNOR2_X1 U673 ( .A(KEYINPUT69), .B(n603), .ZN(n606) );
  NAND2_X1 U674 ( .A1(n658), .A2(G81), .ZN(n604) );
  XOR2_X1 U675 ( .A(KEYINPUT12), .B(n604), .Z(n605) );
  NOR2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT13), .ZN(n608) );
  NOR2_X1 U678 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U679 ( .A(n610), .B(KEYINPUT70), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G43), .A2(n654), .ZN(n611) );
  NAND2_X1 U681 ( .A1(n612), .A2(n611), .ZN(n955) );
  INV_X1 U682 ( .A(G860), .ZN(n826) );
  OR2_X1 U683 ( .A1(n955), .A2(n826), .ZN(G153) );
  INV_X1 U684 ( .A(G171), .ZN(G301) );
  NAND2_X1 U685 ( .A1(G92), .A2(n658), .ZN(n613) );
  NAND2_X1 U686 ( .A1(G54), .A2(n654), .ZN(n614) );
  NAND2_X1 U687 ( .A1(n521), .A2(n614), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G79), .A2(n657), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G66), .A2(n653), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U691 ( .A(n619), .B(KEYINPUT15), .ZN(n620) );
  XOR2_X2 U692 ( .A(KEYINPUT72), .B(n620), .Z(n935) );
  NOR2_X1 U693 ( .A1(n935), .A2(G868), .ZN(n622) );
  INV_X1 U694 ( .A(G868), .ZN(n673) );
  NOR2_X1 U695 ( .A1(n673), .A2(G301), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n622), .A2(n621), .ZN(G284) );
  NAND2_X1 U697 ( .A1(G286), .A2(G868), .ZN(n624) );
  NAND2_X1 U698 ( .A1(G299), .A2(n673), .ZN(n623) );
  NAND2_X1 U699 ( .A1(n624), .A2(n623), .ZN(G297) );
  NAND2_X1 U700 ( .A1(n826), .A2(G559), .ZN(n625) );
  INV_X1 U701 ( .A(n935), .ZN(n670) );
  NAND2_X1 U702 ( .A1(n625), .A2(n670), .ZN(n626) );
  XNOR2_X1 U703 ( .A(n626), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U704 ( .A1(G868), .A2(n955), .ZN(n629) );
  NAND2_X1 U705 ( .A1(n670), .A2(G868), .ZN(n627) );
  NOR2_X1 U706 ( .A1(G559), .A2(n627), .ZN(n628) );
  NOR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(G282) );
  NAND2_X1 U708 ( .A1(G135), .A2(n888), .ZN(n631) );
  NAND2_X1 U709 ( .A1(G111), .A2(n892), .ZN(n630) );
  NAND2_X1 U710 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U711 ( .A1(n893), .A2(G123), .ZN(n632) );
  XOR2_X1 U712 ( .A(KEYINPUT18), .B(n632), .Z(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n636) );
  NAND2_X1 U714 ( .A1(n886), .A2(G99), .ZN(n635) );
  NAND2_X1 U715 ( .A1(n636), .A2(n635), .ZN(n970) );
  XOR2_X1 U716 ( .A(n970), .B(G2096), .Z(n638) );
  XNOR2_X1 U717 ( .A(G2100), .B(KEYINPUT75), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(G156) );
  NAND2_X1 U719 ( .A1(G49), .A2(n654), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G74), .A2(G651), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U722 ( .A1(n653), .A2(n641), .ZN(n644) );
  NAND2_X1 U723 ( .A1(n642), .A2(G87), .ZN(n643) );
  NAND2_X1 U724 ( .A1(n644), .A2(n643), .ZN(G288) );
  NAND2_X1 U725 ( .A1(G48), .A2(n654), .ZN(n645) );
  XNOR2_X1 U726 ( .A(n645), .B(KEYINPUT78), .ZN(n652) );
  NAND2_X1 U727 ( .A1(G86), .A2(n658), .ZN(n647) );
  NAND2_X1 U728 ( .A1(G61), .A2(n653), .ZN(n646) );
  NAND2_X1 U729 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n657), .A2(G73), .ZN(n648) );
  XOR2_X1 U731 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U733 ( .A1(n652), .A2(n651), .ZN(G305) );
  XNOR2_X1 U734 ( .A(G166), .B(G299), .ZN(n664) );
  NAND2_X1 U735 ( .A1(G67), .A2(n653), .ZN(n656) );
  NAND2_X1 U736 ( .A1(G55), .A2(n654), .ZN(n655) );
  NAND2_X1 U737 ( .A1(n656), .A2(n655), .ZN(n662) );
  NAND2_X1 U738 ( .A1(G80), .A2(n657), .ZN(n660) );
  NAND2_X1 U739 ( .A1(G93), .A2(n658), .ZN(n659) );
  NAND2_X1 U740 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U741 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U742 ( .A(n663), .B(KEYINPUT76), .Z(n825) );
  XOR2_X1 U743 ( .A(n664), .B(n825), .Z(n665) );
  XNOR2_X1 U744 ( .A(KEYINPUT19), .B(n665), .ZN(n667) );
  XNOR2_X1 U745 ( .A(G288), .B(KEYINPUT81), .ZN(n666) );
  XNOR2_X1 U746 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U747 ( .A(n668), .B(G290), .ZN(n669) );
  XNOR2_X1 U748 ( .A(n669), .B(G305), .ZN(n832) );
  NAND2_X1 U749 ( .A1(n670), .A2(G559), .ZN(n671) );
  XOR2_X1 U750 ( .A(n955), .B(n671), .Z(n827) );
  XOR2_X1 U751 ( .A(n832), .B(n827), .Z(n672) );
  NOR2_X1 U752 ( .A1(n673), .A2(n672), .ZN(n675) );
  NOR2_X1 U753 ( .A1(n825), .A2(G868), .ZN(n674) );
  NOR2_X1 U754 ( .A1(n675), .A2(n674), .ZN(G295) );
  NAND2_X1 U755 ( .A1(G2078), .A2(G2084), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT20), .B(n676), .Z(n677) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n677), .ZN(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U761 ( .A1(G132), .A2(G82), .ZN(n680) );
  XNOR2_X1 U762 ( .A(n680), .B(KEYINPUT82), .ZN(n681) );
  XNOR2_X1 U763 ( .A(n681), .B(KEYINPUT22), .ZN(n682) );
  NOR2_X1 U764 ( .A1(G218), .A2(n682), .ZN(n683) );
  NAND2_X1 U765 ( .A1(G96), .A2(n683), .ZN(n830) );
  NAND2_X1 U766 ( .A1(n830), .A2(G2106), .ZN(n687) );
  NAND2_X1 U767 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U768 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U769 ( .A1(G108), .A2(n685), .ZN(n831) );
  NAND2_X1 U770 ( .A1(n831), .A2(G567), .ZN(n686) );
  NAND2_X1 U771 ( .A1(n687), .A2(n686), .ZN(n912) );
  NAND2_X1 U772 ( .A1(G661), .A2(G483), .ZN(n688) );
  NOR2_X1 U773 ( .A1(n912), .A2(n688), .ZN(n824) );
  NAND2_X1 U774 ( .A1(n824), .A2(G36), .ZN(G176) );
  INV_X1 U775 ( .A(G166), .ZN(G303) );
  NAND2_X1 U776 ( .A1(G40), .A2(G160), .ZN(n770) );
  XNOR2_X1 U777 ( .A(n770), .B(KEYINPUT83), .ZN(n689) );
  NOR2_X1 U778 ( .A1(G164), .A2(G1384), .ZN(n772) );
  BUF_X2 U779 ( .A(n723), .Z(n735) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n735), .ZN(n691) );
  INV_X1 U781 ( .A(n735), .ZN(n695) );
  NAND2_X1 U782 ( .A1(G2067), .A2(n695), .ZN(n690) );
  NAND2_X1 U783 ( .A1(n691), .A2(n690), .ZN(n699) );
  NAND2_X1 U784 ( .A1(n935), .A2(n699), .ZN(n693) );
  NAND2_X1 U785 ( .A1(G1341), .A2(n735), .ZN(n692) );
  NAND2_X1 U786 ( .A1(n693), .A2(n692), .ZN(n694) );
  NOR2_X1 U787 ( .A1(n955), .A2(n694), .ZN(n698) );
  NAND2_X1 U788 ( .A1(n695), .A2(G1996), .ZN(n696) );
  XNOR2_X1 U789 ( .A(n696), .B(KEYINPUT26), .ZN(n697) );
  NAND2_X1 U790 ( .A1(n698), .A2(n697), .ZN(n710) );
  NOR2_X1 U791 ( .A1(n935), .A2(n699), .ZN(n708) );
  INV_X1 U792 ( .A(n723), .ZN(n700) );
  NAND2_X1 U793 ( .A1(n700), .A2(G2072), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n702), .B(n701), .ZN(n704) );
  NAND2_X1 U795 ( .A1(G1956), .A2(n735), .ZN(n703) );
  NAND2_X1 U796 ( .A1(n704), .A2(n703), .ZN(n706) );
  INV_X1 U797 ( .A(KEYINPUT89), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n712), .A2(G299), .ZN(n707) );
  NOR2_X1 U799 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U800 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U801 ( .A(KEYINPUT91), .B(n711), .ZN(n717) );
  NAND2_X1 U802 ( .A1(G299), .A2(n712), .ZN(n715) );
  XNOR2_X1 U803 ( .A(n718), .B(KEYINPUT29), .ZN(n722) );
  XNOR2_X1 U804 ( .A(KEYINPUT25), .B(G2078), .ZN(n914) );
  NOR2_X1 U805 ( .A1(n735), .A2(n914), .ZN(n720) );
  AND2_X1 U806 ( .A1(n735), .A2(G1961), .ZN(n719) );
  NOR2_X1 U807 ( .A1(n720), .A2(n719), .ZN(n728) );
  NAND2_X1 U808 ( .A1(G171), .A2(n728), .ZN(n721) );
  NAND2_X1 U809 ( .A1(n722), .A2(n721), .ZN(n734) );
  NOR2_X1 U810 ( .A1(G1966), .A2(n765), .ZN(n747) );
  NOR2_X1 U811 ( .A1(G2084), .A2(n735), .ZN(n744) );
  NOR2_X1 U812 ( .A1(n747), .A2(n744), .ZN(n724) );
  XNOR2_X1 U813 ( .A(n724), .B(KEYINPUT92), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n725), .A2(G8), .ZN(n726) );
  XNOR2_X1 U815 ( .A(n726), .B(KEYINPUT30), .ZN(n727) );
  NOR2_X1 U816 ( .A1(G168), .A2(n727), .ZN(n730) );
  NOR2_X1 U817 ( .A1(G171), .A2(n728), .ZN(n729) );
  NOR2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U819 ( .A(KEYINPUT93), .B(n731), .ZN(n732) );
  XNOR2_X1 U820 ( .A(n732), .B(KEYINPUT31), .ZN(n733) );
  NAND2_X1 U821 ( .A1(n734), .A2(n733), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n745), .A2(G286), .ZN(n740) );
  NOR2_X1 U823 ( .A1(G1971), .A2(n765), .ZN(n737) );
  NOR2_X1 U824 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U825 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U826 ( .A1(n738), .A2(G303), .ZN(n739) );
  NAND2_X1 U827 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U828 ( .A(n741), .B(KEYINPUT94), .ZN(n742) );
  NAND2_X1 U829 ( .A1(n742), .A2(G8), .ZN(n743) );
  XNOR2_X1 U830 ( .A(n743), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U831 ( .A1(G8), .A2(n744), .ZN(n749) );
  INV_X1 U832 ( .A(n745), .ZN(n746) );
  NOR2_X1 U833 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U834 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U835 ( .A1(n751), .A2(n750), .ZN(n759) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n952) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n950) );
  NOR2_X1 U838 ( .A1(n952), .A2(n950), .ZN(n752) );
  NAND2_X1 U839 ( .A1(n759), .A2(n752), .ZN(n754) );
  NOR2_X1 U840 ( .A1(n765), .A2(n522), .ZN(n753) );
  AND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  XNOR2_X1 U842 ( .A(n756), .B(KEYINPUT95), .ZN(n758) );
  NAND2_X1 U843 ( .A1(KEYINPUT33), .A2(n950), .ZN(n757) );
  XOR2_X1 U844 ( .A(G1981), .B(G305), .Z(n944) );
  NAND2_X1 U845 ( .A1(n526), .A2(n944), .ZN(n769) );
  NOR2_X1 U846 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U847 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U848 ( .A1(n759), .A2(n761), .ZN(n762) );
  NAND2_X1 U849 ( .A1(n762), .A2(n765), .ZN(n768) );
  NOR2_X1 U850 ( .A1(G1981), .A2(G305), .ZN(n763) );
  XOR2_X1 U851 ( .A(n763), .B(KEYINPUT24), .Z(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n766) );
  XOR2_X1 U853 ( .A(n766), .B(KEYINPUT88), .Z(n767) );
  NAND2_X1 U854 ( .A1(n769), .A2(n524), .ZN(n804) );
  XOR2_X1 U855 ( .A(KEYINPUT83), .B(n770), .Z(n771) );
  NOR2_X1 U856 ( .A1(n772), .A2(n771), .ZN(n815) );
  NAND2_X1 U857 ( .A1(G140), .A2(n888), .ZN(n774) );
  NAND2_X1 U858 ( .A1(G104), .A2(n886), .ZN(n773) );
  NAND2_X1 U859 ( .A1(n774), .A2(n773), .ZN(n775) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n775), .ZN(n780) );
  NAND2_X1 U861 ( .A1(G116), .A2(n892), .ZN(n777) );
  NAND2_X1 U862 ( .A1(G128), .A2(n893), .ZN(n776) );
  NAND2_X1 U863 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U864 ( .A(n778), .B(KEYINPUT35), .Z(n779) );
  NOR2_X1 U865 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U866 ( .A(KEYINPUT36), .B(n781), .Z(n782) );
  XNOR2_X1 U867 ( .A(KEYINPUT84), .B(n782), .ZN(n871) );
  XOR2_X1 U868 ( .A(G2067), .B(KEYINPUT37), .Z(n813) );
  NAND2_X1 U869 ( .A1(n871), .A2(n813), .ZN(n783) );
  XNOR2_X1 U870 ( .A(n783), .B(KEYINPUT85), .ZN(n976) );
  NAND2_X1 U871 ( .A1(n815), .A2(n976), .ZN(n811) );
  NAND2_X1 U872 ( .A1(G95), .A2(n886), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G119), .A2(n893), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n888), .A2(G131), .ZN(n786) );
  XOR2_X1 U876 ( .A(KEYINPUT86), .B(n786), .Z(n787) );
  NOR2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U878 ( .A1(n892), .A2(G107), .ZN(n789) );
  NAND2_X1 U879 ( .A1(n790), .A2(n789), .ZN(n899) );
  AND2_X1 U880 ( .A1(n899), .A2(G1991), .ZN(n799) );
  NAND2_X1 U881 ( .A1(G141), .A2(n888), .ZN(n792) );
  NAND2_X1 U882 ( .A1(G117), .A2(n892), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n795) );
  NAND2_X1 U884 ( .A1(n886), .A2(G105), .ZN(n793) );
  XOR2_X1 U885 ( .A(KEYINPUT38), .B(n793), .Z(n794) );
  NOR2_X1 U886 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U887 ( .A1(n893), .A2(G129), .ZN(n796) );
  NAND2_X1 U888 ( .A1(n797), .A2(n796), .ZN(n883) );
  AND2_X1 U889 ( .A1(n883), .A2(G1996), .ZN(n798) );
  NOR2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n984) );
  INV_X1 U891 ( .A(n984), .ZN(n800) );
  NAND2_X1 U892 ( .A1(n800), .A2(n815), .ZN(n805) );
  NAND2_X1 U893 ( .A1(n811), .A2(n805), .ZN(n801) );
  XOR2_X1 U894 ( .A(KEYINPUT87), .B(n801), .Z(n802) );
  XNOR2_X1 U895 ( .A(G1986), .B(G290), .ZN(n937) );
  NAND2_X1 U896 ( .A1(n804), .A2(n803), .ZN(n818) );
  NOR2_X1 U897 ( .A1(G1996), .A2(n883), .ZN(n979) );
  INV_X1 U898 ( .A(n805), .ZN(n808) );
  NOR2_X1 U899 ( .A1(G1986), .A2(G290), .ZN(n806) );
  NOR2_X1 U900 ( .A1(G1991), .A2(n899), .ZN(n973) );
  NOR2_X1 U901 ( .A1(n806), .A2(n973), .ZN(n807) );
  NOR2_X1 U902 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U903 ( .A1(n979), .A2(n809), .ZN(n810) );
  XNOR2_X1 U904 ( .A(KEYINPUT39), .B(n810), .ZN(n812) );
  NAND2_X1 U905 ( .A1(n812), .A2(n811), .ZN(n814) );
  OR2_X1 U906 ( .A1(n871), .A2(n813), .ZN(n983) );
  NAND2_X1 U907 ( .A1(n814), .A2(n983), .ZN(n816) );
  NAND2_X1 U908 ( .A1(n816), .A2(n815), .ZN(n817) );
  NAND2_X1 U909 ( .A1(n818), .A2(n817), .ZN(n819) );
  XNOR2_X1 U910 ( .A(KEYINPUT40), .B(n819), .ZN(G329) );
  NAND2_X1 U911 ( .A1(n820), .A2(G2106), .ZN(n821) );
  XNOR2_X1 U912 ( .A(n821), .B(KEYINPUT98), .ZN(G217) );
  AND2_X1 U913 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U914 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U915 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(G188) );
  XOR2_X1 U918 ( .A(n825), .B(KEYINPUT77), .Z(n829) );
  NAND2_X1 U919 ( .A1(n827), .A2(n826), .ZN(n828) );
  XNOR2_X1 U920 ( .A(n829), .B(n828), .ZN(G145) );
  INV_X1 U921 ( .A(G132), .ZN(G219) );
  INV_X1 U922 ( .A(G120), .ZN(G236) );
  INV_X1 U923 ( .A(G82), .ZN(G220) );
  INV_X1 U924 ( .A(G69), .ZN(G235) );
  NOR2_X1 U925 ( .A1(n831), .A2(n830), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(n832), .B(G286), .Z(n834) );
  XNOR2_X1 U928 ( .A(G171), .B(n935), .ZN(n833) );
  XNOR2_X1 U929 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U930 ( .A(n835), .B(n955), .Z(n836) );
  NOR2_X1 U931 ( .A1(G37), .A2(n836), .ZN(G397) );
  XOR2_X1 U932 ( .A(G2096), .B(G2090), .Z(n838) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2072), .ZN(n837) );
  XNOR2_X1 U934 ( .A(n838), .B(n837), .ZN(n848) );
  XOR2_X1 U935 ( .A(KEYINPUT100), .B(G2678), .Z(n840) );
  XNOR2_X1 U936 ( .A(KEYINPUT99), .B(KEYINPUT102), .ZN(n839) );
  XNOR2_X1 U937 ( .A(n840), .B(n839), .ZN(n844) );
  XOR2_X1 U938 ( .A(G2100), .B(KEYINPUT101), .Z(n842) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n841) );
  XNOR2_X1 U940 ( .A(n842), .B(n841), .ZN(n843) );
  XOR2_X1 U941 ( .A(n844), .B(n843), .Z(n846) );
  XNOR2_X1 U942 ( .A(G2078), .B(G2084), .ZN(n845) );
  XNOR2_X1 U943 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U944 ( .A(n848), .B(n847), .Z(G227) );
  XOR2_X1 U945 ( .A(G1956), .B(G1966), .Z(n850) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1976), .ZN(n849) );
  XNOR2_X1 U947 ( .A(n850), .B(n849), .ZN(n854) );
  XOR2_X1 U948 ( .A(G1961), .B(G1981), .Z(n852) );
  XNOR2_X1 U949 ( .A(G1996), .B(G1991), .ZN(n851) );
  XNOR2_X1 U950 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U951 ( .A(n854), .B(n853), .Z(n856) );
  XNOR2_X1 U952 ( .A(G2474), .B(KEYINPUT41), .ZN(n855) );
  XNOR2_X1 U953 ( .A(n856), .B(n855), .ZN(n858) );
  XOR2_X1 U954 ( .A(G1971), .B(KEYINPUT103), .Z(n857) );
  XNOR2_X1 U955 ( .A(n858), .B(n857), .ZN(G229) );
  NAND2_X1 U956 ( .A1(G124), .A2(n893), .ZN(n859) );
  XNOR2_X1 U957 ( .A(n859), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G100), .A2(n886), .ZN(n860) );
  XOR2_X1 U959 ( .A(KEYINPUT105), .B(n860), .Z(n861) );
  NAND2_X1 U960 ( .A1(n862), .A2(n861), .ZN(n867) );
  NAND2_X1 U961 ( .A1(n888), .A2(G136), .ZN(n863) );
  XNOR2_X1 U962 ( .A(n863), .B(KEYINPUT104), .ZN(n865) );
  NAND2_X1 U963 ( .A1(G112), .A2(n892), .ZN(n864) );
  NAND2_X1 U964 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U965 ( .A1(n867), .A2(n866), .ZN(G162) );
  XOR2_X1 U966 ( .A(KEYINPUT110), .B(KEYINPUT109), .Z(n869) );
  XNOR2_X1 U967 ( .A(KEYINPUT48), .B(KEYINPUT46), .ZN(n868) );
  XNOR2_X1 U968 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(n870), .B(G162), .Z(n873) );
  XOR2_X1 U970 ( .A(G164), .B(n871), .Z(n872) );
  XNOR2_X1 U971 ( .A(n873), .B(n872), .ZN(n874) );
  XNOR2_X1 U972 ( .A(n970), .B(n874), .ZN(n885) );
  NAND2_X1 U973 ( .A1(G139), .A2(n888), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G103), .A2(n886), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n882) );
  NAND2_X1 U976 ( .A1(n893), .A2(G127), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT108), .ZN(n879) );
  NAND2_X1 U978 ( .A1(G115), .A2(n892), .ZN(n878) );
  NAND2_X1 U979 ( .A1(n879), .A2(n878), .ZN(n880) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n880), .Z(n881) );
  NOR2_X1 U981 ( .A1(n882), .A2(n881), .ZN(n965) );
  XOR2_X1 U982 ( .A(n883), .B(n965), .Z(n884) );
  XNOR2_X1 U983 ( .A(n885), .B(n884), .ZN(n903) );
  NAND2_X1 U984 ( .A1(n886), .A2(G106), .ZN(n887) );
  XOR2_X1 U985 ( .A(KEYINPUT107), .B(n887), .Z(n890) );
  NAND2_X1 U986 ( .A1(n888), .A2(G142), .ZN(n889) );
  NAND2_X1 U987 ( .A1(n890), .A2(n889), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n891), .B(KEYINPUT45), .ZN(n898) );
  NAND2_X1 U989 ( .A1(G118), .A2(n892), .ZN(n895) );
  NAND2_X1 U990 ( .A1(G130), .A2(n893), .ZN(n894) );
  NAND2_X1 U991 ( .A1(n895), .A2(n894), .ZN(n896) );
  XOR2_X1 U992 ( .A(KEYINPUT106), .B(n896), .Z(n897) );
  NAND2_X1 U993 ( .A1(n898), .A2(n897), .ZN(n900) );
  XOR2_X1 U994 ( .A(n900), .B(n899), .Z(n901) );
  XOR2_X1 U995 ( .A(G160), .B(n901), .Z(n902) );
  XNOR2_X1 U996 ( .A(n903), .B(n902), .ZN(n904) );
  NOR2_X1 U997 ( .A1(G37), .A2(n904), .ZN(n905) );
  XOR2_X1 U998 ( .A(KEYINPUT111), .B(n905), .Z(G395) );
  NOR2_X1 U999 ( .A1(G227), .A2(G229), .ZN(n906) );
  XNOR2_X1 U1000 ( .A(KEYINPUT49), .B(n906), .ZN(n907) );
  NOR2_X1 U1001 ( .A1(G397), .A2(n907), .ZN(n911) );
  NOR2_X1 U1002 ( .A1(n912), .A2(G401), .ZN(n908) );
  XOR2_X1 U1003 ( .A(KEYINPUT112), .B(n908), .Z(n909) );
  NOR2_X1 U1004 ( .A1(G395), .A2(n909), .ZN(n910) );
  NAND2_X1 U1005 ( .A1(n911), .A2(n910), .ZN(G225) );
  INV_X1 U1006 ( .A(G225), .ZN(G308) );
  INV_X1 U1007 ( .A(n912), .ZN(G319) );
  INV_X1 U1008 ( .A(G96), .ZN(G221) );
  INV_X1 U1009 ( .A(G108), .ZN(G238) );
  INV_X1 U1010 ( .A(KEYINPUT55), .ZN(n991) );
  XOR2_X1 U1011 ( .A(G25), .B(G1991), .Z(n913) );
  NAND2_X1 U1012 ( .A1(n913), .A2(G28), .ZN(n923) );
  XNOR2_X1 U1013 ( .A(G27), .B(n914), .ZN(n921) );
  XNOR2_X1 U1014 ( .A(G1996), .B(G32), .ZN(n919) );
  XNOR2_X1 U1015 ( .A(G2067), .B(G26), .ZN(n916) );
  XNOR2_X1 U1016 ( .A(G2072), .B(G33), .ZN(n915) );
  NOR2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(KEYINPUT117), .B(n917), .ZN(n918) );
  NOR2_X1 U1019 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1021 ( .A1(n923), .A2(n922), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n924) );
  XNOR2_X1 U1023 ( .A(n925), .B(n924), .ZN(n927) );
  XNOR2_X1 U1024 ( .A(G35), .B(G2090), .ZN(n926) );
  NOR2_X1 U1025 ( .A1(n927), .A2(n926), .ZN(n930) );
  XOR2_X1 U1026 ( .A(G2084), .B(G34), .Z(n928) );
  XNOR2_X1 U1027 ( .A(KEYINPUT54), .B(n928), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  XNOR2_X1 U1029 ( .A(n991), .B(n931), .ZN(n933) );
  INV_X1 U1030 ( .A(G29), .ZN(n932) );
  NAND2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(G11), .A2(n934), .ZN(n964) );
  XNOR2_X1 U1033 ( .A(KEYINPUT56), .B(G16), .ZN(n961) );
  XNOR2_X1 U1034 ( .A(G1348), .B(n935), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n936), .B(KEYINPUT119), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n522), .A2(n937), .ZN(n938) );
  NAND2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n941) );
  XNOR2_X1 U1038 ( .A(G1956), .B(G299), .ZN(n940) );
  NOR2_X1 U1039 ( .A1(n941), .A2(n940), .ZN(n943) );
  NAND2_X1 U1040 ( .A1(G1971), .A2(G303), .ZN(n942) );
  NAND2_X1 U1041 ( .A1(n943), .A2(n942), .ZN(n948) );
  XNOR2_X1 U1042 ( .A(G1966), .B(G168), .ZN(n945) );
  NAND2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1044 ( .A(KEYINPUT57), .B(n946), .Z(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n959) );
  XNOR2_X1 U1046 ( .A(G1961), .B(G171), .ZN(n949) );
  XNOR2_X1 U1047 ( .A(n949), .B(KEYINPUT120), .ZN(n954) );
  XOR2_X1 U1048 ( .A(n950), .B(KEYINPUT121), .Z(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1055 ( .A(KEYINPUT122), .B(n962), .Z(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n995) );
  XOR2_X1 U1057 ( .A(G164), .B(G2078), .Z(n968) );
  XOR2_X1 U1058 ( .A(n965), .B(KEYINPUT116), .Z(n966) );
  XNOR2_X1 U1059 ( .A(G2072), .B(n966), .ZN(n967) );
  NOR2_X1 U1060 ( .A1(n968), .A2(n967), .ZN(n969) );
  XOR2_X1 U1061 ( .A(KEYINPUT50), .B(n969), .Z(n989) );
  XNOR2_X1 U1062 ( .A(G160), .B(G2084), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  NOR2_X1 U1064 ( .A1(n973), .A2(n972), .ZN(n974) );
  XNOR2_X1 U1065 ( .A(n974), .B(KEYINPUT113), .ZN(n975) );
  NOR2_X1 U1066 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1067 ( .A(KEYINPUT114), .B(n977), .ZN(n982) );
  XOR2_X1 U1068 ( .A(G2090), .B(G162), .Z(n978) );
  NOR2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1070 ( .A(KEYINPUT51), .B(n980), .Z(n981) );
  NAND2_X1 U1071 ( .A1(n982), .A2(n981), .ZN(n986) );
  NAND2_X1 U1072 ( .A1(n984), .A2(n983), .ZN(n985) );
  NOR2_X1 U1073 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1074 ( .A(KEYINPUT115), .B(n987), .ZN(n988) );
  NOR2_X1 U1075 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1076 ( .A(KEYINPUT52), .B(n990), .ZN(n992) );
  NAND2_X1 U1077 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1078 ( .A1(n993), .A2(G29), .ZN(n994) );
  NAND2_X1 U1079 ( .A1(n995), .A2(n994), .ZN(n1023) );
  XNOR2_X1 U1080 ( .A(G1348), .B(KEYINPUT59), .ZN(n996) );
  XNOR2_X1 U1081 ( .A(n996), .B(G4), .ZN(n1004) );
  XOR2_X1 U1082 ( .A(G1956), .B(G20), .Z(n997) );
  XNOR2_X1 U1083 ( .A(KEYINPUT123), .B(n997), .ZN(n1002) );
  XNOR2_X1 U1084 ( .A(G1981), .B(G6), .ZN(n999) );
  XNOR2_X1 U1085 ( .A(G19), .B(G1341), .ZN(n998) );
  NOR2_X1 U1086 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1087 ( .A(KEYINPUT124), .B(n1000), .Z(n1001) );
  NOR2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1006) );
  XNOR2_X1 U1090 ( .A(KEYINPUT125), .B(KEYINPUT60), .ZN(n1005) );
  XNOR2_X1 U1091 ( .A(n1006), .B(n1005), .ZN(n1017) );
  XNOR2_X1 U1092 ( .A(G1986), .B(G24), .ZN(n1012) );
  XNOR2_X1 U1093 ( .A(G1971), .B(G22), .ZN(n1007) );
  XNOR2_X1 U1094 ( .A(n1007), .B(KEYINPUT126), .ZN(n1009) );
  XNOR2_X1 U1095 ( .A(G23), .B(G1976), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1097 ( .A(KEYINPUT127), .B(n1010), .ZN(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1099 ( .A(KEYINPUT58), .B(n1013), .Z(n1015) );
  XNOR2_X1 U1100 ( .A(G1966), .B(G21), .ZN(n1014) );
  NOR2_X1 U1101 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NAND2_X1 U1102 ( .A1(n1017), .A2(n1016), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(G5), .B(G1961), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1020), .Z(n1021) );
  NOR2_X1 U1106 ( .A1(G16), .A2(n1021), .ZN(n1022) );
  NOR2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(n1024), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

