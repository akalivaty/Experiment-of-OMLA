//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 0 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n552, new_n553, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n576,
    new_n577, new_n578, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n607, new_n608, new_n611,
    new_n613, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT67), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT68), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n459), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n465));
  NOR3_X1   g040(.A1(new_n464), .A2(G2105), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G137), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n459), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G125), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n468), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G2105), .ZN(new_n474));
  XNOR2_X1  g049(.A(KEYINPUT68), .B(G2104), .ZN(new_n475));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(G101), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n467), .A2(new_n474), .A3(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(G160));
  OAI211_X1 g054(.A(G2105), .B(new_n469), .C1(new_n475), .C2(new_n459), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n466), .A2(G136), .ZN(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n476), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n488), .A2(new_n476), .A3(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n471), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n462), .A2(G2104), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n460), .A2(KEYINPUT68), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT3), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n493), .A2(G138), .A3(new_n476), .A4(new_n469), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n490), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  NOR2_X1   g071(.A1(new_n476), .A2(G114), .ZN(new_n497));
  OAI21_X1  g072(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n480), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n495), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(G651), .ZN(new_n503));
  OAI21_X1  g078(.A(KEYINPUT6), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT69), .A3(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G50), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n501), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n517), .A2(new_n503), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n509), .A2(KEYINPUT70), .A3(G50), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n513), .A2(new_n515), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n507), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G88), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n512), .A2(new_n518), .A3(new_n519), .A4(new_n522), .ZN(G303));
  INV_X1    g098(.A(G303), .ZN(G166));
  AND2_X1   g099(.A1(new_n509), .A2(G51), .ZN(new_n525));
  AND2_X1   g100(.A1(G63), .A2(G651), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n516), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(new_n527), .B2(new_n528), .ZN(new_n530));
  AND2_X1   g105(.A1(new_n521), .A2(G89), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n525), .A2(new_n530), .A3(new_n531), .ZN(G168));
  NAND2_X1  g107(.A1(new_n521), .A2(G90), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n509), .A2(G52), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n535));
  OAI211_X1 g110(.A(new_n533), .B(new_n534), .C1(new_n503), .C2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n537));
  OR2_X1    g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n537), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n520), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT72), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n543), .A2(new_n544), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n545), .A2(G651), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g122(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n547), .A2(KEYINPUT73), .ZN(new_n549));
  AOI22_X1  g124(.A1(G43), .A2(new_n509), .B1(new_n521), .B2(G81), .ZN(new_n550));
  NAND4_X1  g125(.A1(new_n548), .A2(G860), .A3(new_n549), .A4(new_n550), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT74), .Z(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  NAND2_X1  g132(.A1(new_n509), .A2(G53), .ZN(new_n558));
  AND2_X1   g133(.A1(KEYINPUT75), .A2(KEYINPUT9), .ZN(new_n559));
  XOR2_X1   g134(.A(new_n558), .B(new_n559), .Z(new_n560));
  INV_X1    g135(.A(KEYINPUT76), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(new_n521), .ZN(new_n563));
  INV_X1    g138(.A(G91), .ZN(new_n564));
  OR3_X1    g139(.A1(new_n563), .A2(KEYINPUT77), .A3(new_n564), .ZN(new_n565));
  OAI21_X1  g140(.A(KEYINPUT77), .B1(new_n563), .B2(new_n564), .ZN(new_n566));
  NAND2_X1  g141(.A1(G78), .A2(G543), .ZN(new_n567));
  INV_X1    g142(.A(G65), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n520), .B2(new_n568), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n565), .A2(new_n566), .B1(G651), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n558), .B(new_n559), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(KEYINPUT76), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n562), .A2(new_n570), .A3(new_n572), .ZN(G299));
  INV_X1    g148(.A(G171), .ZN(G301));
  INV_X1    g149(.A(G168), .ZN(G286));
  OAI21_X1  g150(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n516), .A2(G87), .A3(new_n504), .A4(new_n506), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n504), .A2(G49), .A3(G543), .A4(new_n506), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(G288));
  NAND2_X1  g154(.A1(new_n509), .A2(G48), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n521), .A2(G86), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n520), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n584), .A2(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n580), .A2(new_n581), .A3(new_n585), .ZN(G305));
  NAND2_X1  g161(.A1(new_n521), .A2(G85), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n588));
  XNOR2_X1  g163(.A(KEYINPUT78), .B(G47), .ZN(new_n589));
  OAI221_X1 g164(.A(new_n587), .B1(new_n588), .B2(new_n503), .C1(new_n510), .C2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  AND2_X1   g166(.A1(new_n521), .A2(G92), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT10), .ZN(new_n593));
  INV_X1    g168(.A(G54), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT79), .ZN(new_n595));
  AOI21_X1  g170(.A(new_n594), .B1(new_n510), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n509), .A2(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(G79), .A2(G543), .ZN(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n520), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n596), .A2(new_n597), .B1(G651), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT80), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n602), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n591), .B1(new_n604), .B2(G868), .ZN(G284));
  OAI21_X1  g180(.A(new_n591), .B1(new_n604), .B2(G868), .ZN(G321));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G299), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G297));
  OAI21_X1  g184(.A(new_n608), .B1(new_n607), .B2(G168), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n604), .B1(new_n611), .B2(G860), .ZN(G148));
  NAND3_X1  g187(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(new_n607), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n604), .A2(new_n611), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT81), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n614), .B1(new_n616), .B2(new_n607), .ZN(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g193(.A1(new_n475), .A2(new_n476), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(new_n471), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(KEYINPUT12), .Z(new_n621));
  XOR2_X1   g196(.A(KEYINPUT82), .B(G2100), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n621), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n481), .A2(G123), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n466), .A2(G135), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  INV_X1    g202(.A(KEYINPUT83), .ZN(new_n628));
  INV_X1    g203(.A(G111), .ZN(new_n629));
  AOI22_X1  g204(.A1(new_n627), .A2(new_n628), .B1(new_n629), .B2(G2105), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(new_n628), .B2(new_n627), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n625), .A2(new_n626), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(G2096), .Z(new_n633));
  NAND2_X1  g208(.A1(new_n624), .A2(new_n633), .ZN(G156));
  XNOR2_X1  g209(.A(G2427), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT84), .ZN(new_n636));
  INV_X1    g211(.A(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT15), .B(G2435), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(G2438), .ZN(new_n639));
  OR2_X1    g214(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n639), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n640), .A2(new_n641), .A3(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(G2443), .B(G2446), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT16), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n646), .A2(new_n650), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(new_n653), .ZN(G401));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  OR2_X1    g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n658), .B(KEYINPUT88), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n661), .A2(new_n659), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n660), .A2(KEYINPUT17), .ZN(new_n663));
  OAI221_X1 g238(.A(new_n657), .B1(new_n658), .B2(new_n659), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n655), .A2(new_n658), .A3(new_n656), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT18), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(G227));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT19), .ZN(new_n672));
  XOR2_X1   g247(.A(G1956), .B(G2474), .Z(new_n673));
  XOR2_X1   g248(.A(G1961), .B(G1966), .Z(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OR2_X1    g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n673), .A2(new_n674), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n672), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  OR2_X1    g253(.A1(new_n672), .A2(new_n677), .ZN(new_n679));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n676), .B(new_n678), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n680), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(G1991), .ZN(new_n683));
  INV_X1    g258(.A(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(G1981), .B(G1986), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G229));
  NOR2_X1   g264(.A1(G16), .A2(G23), .ZN(new_n690));
  NAND2_X1  g265(.A1(G288), .A2(KEYINPUT93), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT93), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n576), .A2(new_n577), .A3(new_n692), .A4(new_n578), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n690), .B1(new_n694), .B2(G16), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT33), .B(G1976), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n695), .A2(new_n696), .ZN(new_n698));
  MUX2_X1   g273(.A(G6), .B(G305), .S(G16), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT32), .B(G1981), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT91), .B(KEYINPUT92), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  AOI211_X1 g278(.A(new_n697), .B(new_n698), .C1(new_n701), .C2(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT90), .B(G16), .ZN(new_n705));
  MUX2_X1   g280(.A(G22), .B(G303), .S(new_n705), .Z(new_n706));
  INV_X1    g281(.A(G1971), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n704), .B(new_n708), .C1(new_n703), .C2(new_n701), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT94), .B(KEYINPUT34), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G24), .B(G290), .S(new_n705), .Z(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(G1986), .Z(new_n713));
  NOR2_X1   g288(.A1(G25), .A2(G29), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n481), .A2(G119), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n466), .A2(G131), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n476), .A2(G107), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT89), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n714), .B1(new_n720), .B2(G29), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT35), .B(G1991), .Z(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n711), .A2(new_n713), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT36), .ZN(new_n725));
  INV_X1    g300(.A(G20), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n705), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT23), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(G299), .B2(G16), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(G1956), .ZN(new_n730));
  INV_X1    g305(.A(new_n604), .ZN(new_n731));
  MUX2_X1   g306(.A(G4), .B(new_n731), .S(G16), .Z(new_n732));
  OAI21_X1  g307(.A(new_n730), .B1(new_n732), .B2(G1348), .ZN(new_n733));
  MUX2_X1   g308(.A(G21), .B(G286), .S(G16), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT100), .Z(new_n735));
  NAND2_X1  g310(.A1(new_n735), .A2(G1966), .ZN(new_n736));
  MUX2_X1   g311(.A(G5), .B(G301), .S(G16), .Z(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(G1961), .ZN(new_n738));
  INV_X1    g313(.A(G29), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(G35), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n740), .B1(G162), .B2(new_n739), .ZN(new_n741));
  XOR2_X1   g316(.A(KEYINPUT29), .B(G2090), .Z(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n737), .A2(G1961), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n736), .A2(new_n738), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  AOI211_X1 g320(.A(new_n733), .B(new_n745), .C1(G1348), .C2(new_n732), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n739), .A2(G26), .ZN(new_n747));
  OR2_X1    g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G116), .C2(new_n476), .ZN(new_n749));
  INV_X1    g324(.A(new_n466), .ZN(new_n750));
  INV_X1    g325(.A(G140), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G128), .B2(new_n481), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n747), .B1(new_n754), .B2(G29), .ZN(new_n755));
  MUX2_X1   g330(.A(new_n747), .B(new_n755), .S(KEYINPUT28), .Z(new_n756));
  INV_X1    g331(.A(G2067), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n739), .A2(G33), .ZN(new_n758));
  XOR2_X1   g333(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n759));
  NAND3_X1  g334(.A1(new_n476), .A2(G103), .A3(G2104), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G139), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  NAND3_X1  g339(.A1(new_n469), .A2(new_n470), .A3(G127), .ZN(new_n765));
  NAND2_X1  g340(.A1(G115), .A2(G2104), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n476), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n758), .B1(new_n768), .B2(new_n739), .ZN(new_n769));
  AOI22_X1  g344(.A1(new_n756), .A2(new_n757), .B1(G2072), .B2(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G2072), .B2(new_n769), .ZN(new_n771));
  INV_X1    g346(.A(G28), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT30), .ZN(new_n773));
  AOI21_X1  g348(.A(G29), .B1(new_n772), .B2(KEYINPUT30), .ZN(new_n774));
  OR2_X1    g349(.A1(KEYINPUT31), .A2(G11), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT31), .A2(G11), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n773), .A2(new_n774), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g352(.A1(KEYINPUT24), .A2(G34), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n739), .B1(KEYINPUT24), .B2(G34), .ZN(new_n779));
  OAI22_X1  g354(.A1(G160), .A2(new_n739), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n777), .B1(new_n739), .B2(new_n632), .C1(new_n780), .C2(G2084), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(G2084), .B2(new_n780), .ZN(new_n782));
  INV_X1    g357(.A(G19), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n705), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n613), .B2(new_n705), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT95), .B(G1341), .Z(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n782), .B(new_n787), .C1(new_n735), .C2(G1966), .ZN(new_n788));
  OAI22_X1  g363(.A1(new_n756), .A2(new_n757), .B1(new_n786), .B2(new_n785), .ZN(new_n789));
  NOR3_X1   g364(.A1(new_n771), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NOR2_X1   g365(.A1(G29), .A2(G32), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n481), .A2(G129), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT98), .ZN(new_n793));
  NAND3_X1  g368(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(KEYINPUT26), .Z(new_n795));
  INV_X1    g370(.A(G105), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n619), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(new_n466), .B2(G141), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT99), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n791), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XOR2_X1   g376(.A(KEYINPUT27), .B(G1996), .Z(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n739), .A2(G27), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G164), .B2(new_n739), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT102), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT101), .B(G2078), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n803), .A2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n725), .A2(new_n746), .A3(new_n790), .A4(new_n809), .ZN(G150));
  INV_X1    g385(.A(G150), .ZN(G311));
  NAND2_X1  g386(.A1(new_n604), .A2(G559), .ZN(new_n812));
  XOR2_X1   g387(.A(KEYINPUT38), .B(KEYINPUT39), .Z(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n509), .A2(G55), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT103), .B(G93), .ZN(new_n817));
  OAI221_X1 g392(.A(new_n815), .B1(new_n816), .B2(new_n503), .C1(new_n563), .C2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n613), .B(new_n818), .ZN(new_n819));
  AOI21_X1  g394(.A(G860), .B1(new_n814), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n820), .B1(new_n819), .B2(new_n814), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT104), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n818), .A2(G860), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT37), .Z(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(G145));
  MUX2_X1   g400(.A(new_n799), .B(new_n800), .S(new_n768), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(new_n719), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n753), .B(KEYINPUT105), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n828), .B(G162), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n632), .B(new_n478), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n827), .B(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n466), .A2(G142), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n476), .A2(G118), .ZN(new_n834));
  OAI21_X1  g409(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G130), .B2(new_n481), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(G164), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n621), .Z(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  AND2_X1   g415(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(G37), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n832), .B2(new_n840), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT40), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(G395));
  INV_X1    g421(.A(KEYINPUT81), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n615), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n848), .B(new_n819), .ZN(new_n849));
  INV_X1    g424(.A(new_n602), .ZN(new_n850));
  OR3_X1    g425(.A1(G299), .A2(KEYINPUT107), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(KEYINPUT107), .B1(G299), .B2(new_n850), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(G299), .A2(new_n850), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT106), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n849), .A2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT109), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n859), .A2(KEYINPUT42), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT41), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n854), .B(KEYINPUT106), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n851), .A2(new_n852), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n853), .A2(new_n856), .A3(KEYINPUT41), .ZN(new_n866));
  AND2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI211_X1 g442(.A(new_n858), .B(new_n861), .C1(new_n849), .C2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n819), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n848), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n616), .A2(new_n819), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AND3_X1   g447(.A1(new_n870), .A2(new_n871), .A3(new_n857), .ZN(new_n873));
  OAI21_X1  g448(.A(new_n860), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(G305), .B(KEYINPUT108), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n694), .ZN(new_n876));
  XNOR2_X1  g451(.A(G303), .B(G290), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n876), .B(new_n877), .ZN(new_n878));
  AOI21_X1  g453(.A(new_n878), .B1(new_n859), .B2(KEYINPUT42), .ZN(new_n879));
  AND3_X1   g454(.A1(new_n868), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n879), .B1(new_n868), .B2(new_n874), .ZN(new_n881));
  OAI21_X1  g456(.A(G868), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n818), .A2(new_n607), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(G295));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n883), .ZN(G331));
  NOR2_X1   g460(.A1(KEYINPUT111), .A2(KEYINPUT44), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT111), .ZN(new_n887));
  INV_X1    g462(.A(KEYINPUT44), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n878), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n538), .A2(G168), .A3(new_n539), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G168), .B1(new_n538), .B2(new_n539), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT110), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT110), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n895), .A2(new_n896), .A3(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n898), .A2(new_n869), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n819), .A2(new_n894), .A3(new_n897), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n901), .B1(new_n865), .B2(new_n866), .ZN(new_n902));
  AOI22_X1  g477(.A1(new_n856), .A2(new_n853), .B1(new_n899), .B2(new_n900), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n890), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(new_n842), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n865), .A2(new_n866), .ZN(new_n906));
  INV_X1    g481(.A(new_n901), .ZN(new_n907));
  AOI211_X1 g482(.A(new_n890), .B(new_n903), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OAI21_X1  g483(.A(KEYINPUT43), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n910), .A2(new_n878), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT43), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n911), .A2(new_n912), .A3(new_n842), .A4(new_n904), .ZN(new_n913));
  AOI211_X1 g488(.A(new_n886), .B(new_n889), .C1(new_n909), .C2(new_n913), .ZN(new_n914));
  AND4_X1   g489(.A1(new_n887), .A2(new_n909), .A3(new_n913), .A4(new_n888), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(G397));
  NAND4_X1  g491(.A1(new_n467), .A2(G40), .A3(new_n474), .A4(new_n477), .ZN(new_n917));
  INV_X1    g492(.A(G138), .ZN(new_n918));
  NOR4_X1   g493(.A1(new_n464), .A2(new_n918), .A3(G2105), .A4(new_n465), .ZN(new_n919));
  OAI22_X1  g494(.A1(new_n919), .A2(new_n488), .B1(new_n471), .B2(new_n489), .ZN(new_n920));
  INV_X1    g495(.A(new_n499), .ZN(new_n921));
  AOI21_X1  g496(.A(G1384), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(KEYINPUT112), .B(KEYINPUT45), .Z(new_n923));
  AOI21_X1  g498(.A(new_n917), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G1384), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n495), .B2(new_n499), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(G1966), .B1(new_n924), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G2084), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n926), .A2(KEYINPUT50), .ZN(new_n931));
  INV_X1    g506(.A(new_n917), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT50), .ZN(new_n933));
  OAI211_X1 g508(.A(new_n933), .B(new_n925), .C1(new_n495), .C2(new_n499), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT117), .B1(new_n929), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1966), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n922), .A2(KEYINPUT45), .ZN(new_n938));
  INV_X1    g513(.A(new_n923), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n932), .B1(new_n926), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n937), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT117), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n931), .A2(new_n930), .A3(new_n932), .A4(new_n934), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(G286), .A2(G8), .ZN(new_n945));
  INV_X1    g520(.A(new_n945), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n936), .A2(new_n944), .A3(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n936), .A2(G8), .A3(new_n944), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT118), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT118), .ZN(new_n951));
  NAND4_X1  g526(.A1(new_n936), .A2(new_n944), .A3(new_n951), .A4(G8), .ZN(new_n952));
  XOR2_X1   g527(.A(new_n945), .B(KEYINPUT119), .Z(new_n953));
  NAND3_X1  g528(.A1(new_n950), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT51), .ZN(new_n955));
  INV_X1    g530(.A(G8), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n956), .B1(new_n941), .B2(new_n943), .ZN(new_n957));
  NOR3_X1   g532(.A1(new_n957), .A2(KEYINPUT51), .A3(new_n946), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n948), .B1(new_n955), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n926), .A2(new_n939), .ZN(new_n961));
  INV_X1    g536(.A(G2078), .ZN(new_n962));
  OAI211_X1 g537(.A(KEYINPUT45), .B(new_n925), .C1(new_n495), .C2(new_n499), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n932), .A4(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT53), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n924), .A2(KEYINPUT53), .A3(new_n962), .A4(new_n928), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n968));
  XOR2_X1   g543(.A(KEYINPUT120), .B(G1961), .Z(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n966), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(G171), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT121), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n966), .A2(new_n970), .ZN(new_n974));
  OR2_X1    g549(.A1(new_n964), .A2(new_n965), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(G301), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT121), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n971), .A2(new_n977), .A3(G171), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n973), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT54), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(new_n975), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(G171), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n974), .A2(G301), .A3(new_n967), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n983), .A2(KEYINPUT54), .A3(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n986), .B1(new_n694), .B2(G1976), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n956), .B1(new_n922), .B2(new_n932), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n694), .A2(new_n986), .A3(G1976), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n988), .A2(new_n989), .A3(new_n990), .A4(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(G305), .A2(G1981), .ZN(new_n994));
  INV_X1    g569(.A(G1981), .ZN(new_n995));
  NAND4_X1  g570(.A1(new_n580), .A2(new_n581), .A3(new_n995), .A4(new_n585), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT49), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g574(.A1(new_n994), .A2(KEYINPUT49), .A3(new_n996), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n989), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(G8), .B1(new_n926), .B2(new_n917), .ZN(new_n1002));
  AOI211_X1 g577(.A(KEYINPUT114), .B(new_n991), .C1(new_n691), .C2(new_n693), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1002), .A2(new_n987), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT52), .ZN(new_n1005));
  OAI211_X1 g580(.A(new_n993), .B(new_n1001), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n968), .A2(G2090), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n917), .B1(new_n926), .B2(new_n939), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n963), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n707), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n956), .B1(new_n1007), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(KEYINPUT113), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT55), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(G166), .B2(new_n956), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1013), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1006), .B1(new_n1011), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1017), .ZN(new_n1019));
  OR2_X1    g594(.A1(new_n968), .A2(KEYINPUT115), .ZN(new_n1020));
  AOI21_X1  g595(.A(G2090), .B1(new_n968), .B2(KEYINPUT115), .ZN(new_n1021));
  AOI22_X1  g596(.A1(new_n1020), .A2(new_n1021), .B1(new_n707), .B2(new_n1009), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1019), .B1(new_n1022), .B2(new_n956), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n1018), .A2(new_n1023), .A3(KEYINPUT122), .ZN(new_n1024));
  AOI21_X1  g599(.A(KEYINPUT122), .B1(new_n1018), .B2(new_n1023), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n981), .B(new_n985), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(KEYINPUT123), .B1(new_n960), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(new_n985), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1018), .A2(new_n1023), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT122), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1018), .A2(new_n1023), .A3(KEYINPUT122), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1028), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n1034));
  INV_X1    g609(.A(new_n953), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n949), .B2(KEYINPUT118), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1034), .B1(new_n1036), .B2(new_n952), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n947), .B1(new_n1037), .B2(new_n958), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1033), .A2(new_n1038), .A3(new_n1039), .A4(new_n981), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1009), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  INV_X1    g617(.A(G1956), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1041), .A2(new_n1042), .B1(new_n1043), .B2(new_n968), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n560), .A2(KEYINPUT57), .ZN(new_n1045));
  AOI22_X1  g620(.A1(G299), .A2(KEYINPUT57), .B1(new_n570), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n968), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n922), .A2(new_n932), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1048), .A2(G1348), .B1(G2067), .B2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1051), .A2(new_n731), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1047), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n731), .B1(new_n1051), .B2(KEYINPUT60), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  OR2_X1    g631(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT60), .ZN(new_n1058));
  NOR3_X1   g633(.A1(new_n1050), .A2(new_n604), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1059), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1057), .A2(new_n1060), .B1(new_n1058), .B2(new_n1050), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1041), .A2(new_n684), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND2_X1  g638(.A1(new_n1049), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n613), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  XOR2_X1   g640(.A(new_n1065), .B(KEYINPUT59), .Z(new_n1066));
  INV_X1    g641(.A(new_n1047), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT61), .ZN(new_n1068));
  OR3_X1    g643(.A1(new_n1067), .A2(new_n1068), .A3(new_n1053), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1068), .B1(new_n1067), .B2(new_n1053), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1066), .A2(new_n1069), .A3(new_n1070), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1054), .B1(new_n1061), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1027), .A2(new_n1040), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n958), .B1(new_n954), .B2(KEYINPUT51), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT62), .B1(new_n1074), .B2(new_n948), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT62), .ZN(new_n1076));
  OAI211_X1 g651(.A(new_n1076), .B(new_n947), .C1(new_n1037), .C2(new_n958), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1031), .A2(new_n1032), .B1(new_n978), .B2(new_n973), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1075), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(KEYINPUT124), .ZN(new_n1080));
  INV_X1    g655(.A(new_n1001), .ZN(new_n1081));
  NOR3_X1   g656(.A1(new_n1081), .A2(G1976), .A3(G288), .ZN(new_n1082));
  INV_X1    g657(.A(new_n996), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n989), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1011), .A2(new_n1017), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1084), .B1(new_n1085), .B2(new_n1006), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n957), .A2(G168), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT63), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1090), .B(new_n1018), .C1(new_n1017), .C2(new_n1011), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1089), .B1(new_n1029), .B2(new_n1088), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1086), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT124), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1075), .A2(new_n1094), .A3(new_n1077), .A4(new_n1078), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1073), .A2(new_n1080), .A3(new_n1093), .A4(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n961), .A2(new_n917), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n753), .B(new_n757), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n684), .B1(new_n793), .B2(new_n798), .ZN(new_n1099));
  AOI211_X1 g674(.A(new_n1098), .B(new_n1099), .C1(new_n800), .C2(new_n684), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n719), .B(new_n722), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(G290), .B(G1986), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1097), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1096), .A2(new_n1104), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1097), .B1(new_n1098), .B2(new_n799), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1097), .A2(KEYINPUT46), .A3(new_n684), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT46), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1097), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(G1996), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1106), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  XNOR2_X1  g686(.A(new_n1111), .B(KEYINPUT47), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1109), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n1109), .A2(G1986), .A3(G290), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT48), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n720), .A2(new_n722), .ZN(new_n1116));
  XOR2_X1   g691(.A(new_n1116), .B(KEYINPUT125), .Z(new_n1117));
  AOI22_X1  g692(.A1(new_n1100), .A2(new_n1117), .B1(new_n757), .B2(new_n753), .ZN(new_n1118));
  OAI221_X1 g693(.A(new_n1112), .B1(new_n1113), .B2(new_n1115), .C1(new_n1109), .C2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(new_n1119), .B(KEYINPUT126), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1105), .A2(new_n1120), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g696(.A(G319), .ZN(new_n1123));
  OR3_X1    g697(.A1(G401), .A2(new_n1123), .A3(G227), .ZN(new_n1124));
  NOR2_X1   g698(.A1(G229), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g699(.A(new_n1125), .B1(new_n841), .B2(new_n843), .ZN(new_n1126));
  AND2_X1   g700(.A1(new_n909), .A2(new_n913), .ZN(new_n1127));
  NOR2_X1   g701(.A1(new_n1126), .A2(new_n1127), .ZN(G308));
  INV_X1    g702(.A(G308), .ZN(G225));
endmodule


