//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 1 1 1 1 0 0 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945;
  INV_X1    g000(.A(G472), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT64), .B(G146), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G143), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n193));
  NAND4_X1  g007(.A1(new_n192), .A2(KEYINPUT68), .A3(new_n193), .A4(G128), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(G143), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n190), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n197), .A2(new_n193), .A3(G128), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT68), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n194), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n203));
  XNOR2_X1  g017(.A(KEYINPUT69), .B(G128), .ZN(new_n204));
  INV_X1    g018(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT64), .A2(G146), .ZN(new_n207));
  INV_X1    g021(.A(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT64), .A2(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n189), .A2(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n206), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n202), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  INV_X1    g029(.A(G134), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G137), .ZN(new_n217));
  INV_X1    g031(.A(G137), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G134), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n215), .B1(new_n217), .B2(new_n219), .ZN(new_n220));
  OR2_X1    g034(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT65), .B1(new_n216), .B2(G137), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT11), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n219), .A2(KEYINPUT65), .A3(new_n224), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n223), .A2(new_n225), .A3(new_n215), .A4(new_n217), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n220), .A2(KEYINPUT67), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n221), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT71), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n221), .A2(new_n226), .A3(KEYINPUT71), .A4(new_n227), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n214), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  XNOR2_X1  g046(.A(KEYINPUT2), .B(G113), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OR2_X1    g052(.A1(new_n234), .A2(new_n235), .ZN(new_n239));
  XNOR2_X1  g053(.A(new_n238), .B(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n223), .A2(new_n217), .A3(new_n225), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n215), .A2(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n243), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n223), .A2(new_n225), .A3(new_n245), .A4(new_n217), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT0), .ZN(new_n248));
  INV_X1    g062(.A(G128), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(new_n210), .B2(new_n211), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n248), .A2(new_n249), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n251), .A2(new_n252), .B1(new_n192), .B2(new_n250), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n232), .A2(new_n241), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT28), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AOI22_X1  g071(.A1(new_n194), .A2(new_n201), .B1(new_n212), .B2(new_n206), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n254), .B1(new_n258), .B2(new_n228), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n240), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n232), .A2(new_n241), .A3(KEYINPUT28), .A4(new_n254), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n257), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G237), .ZN(new_n263));
  INV_X1    g077(.A(G953), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n263), .A2(new_n264), .A3(G210), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT74), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT26), .B(G101), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT76), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n262), .A2(KEYINPUT76), .A3(new_n270), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT30), .ZN(new_n275));
  AOI21_X1  g089(.A(KEYINPUT72), .B1(new_n259), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n232), .A2(KEYINPUT30), .A3(new_n254), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND4_X1  g092(.A1(new_n232), .A2(KEYINPUT72), .A3(KEYINPUT30), .A4(new_n254), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n241), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n255), .ZN(new_n281));
  NOR3_X1   g095(.A1(new_n280), .A2(new_n281), .A3(new_n270), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT31), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n273), .B(new_n274), .C1(new_n282), .C2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(KEYINPUT75), .A2(KEYINPUT31), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n279), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n281), .B1(new_n286), .B2(new_n240), .ZN(new_n287));
  INV_X1    g101(.A(new_n270), .ZN(new_n288));
  OR2_X1    g102(.A1(KEYINPUT75), .A2(KEYINPUT31), .ZN(new_n289));
  AND4_X1   g103(.A1(new_n285), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n187), .B(new_n188), .C1(new_n284), .C2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n288), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(KEYINPUT31), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n282), .A2(new_n285), .A3(new_n289), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n273), .A4(new_n274), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n297), .A2(KEYINPUT32), .A3(new_n187), .A4(new_n188), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n287), .A2(new_n270), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n262), .A2(new_n288), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT29), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n232), .A2(new_n254), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n240), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n303), .A2(new_n304), .A3(new_n255), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n302), .A2(KEYINPUT77), .A3(new_n240), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(KEYINPUT28), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n257), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n188), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G472), .B1(new_n301), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n298), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G217), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n313), .B1(G234), .B2(new_n188), .ZN(new_n314));
  INV_X1    g128(.A(G119), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G128), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n317), .B1(new_n315), .B2(G128), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n204), .A2(G119), .ZN(new_n319));
  OAI211_X1 g133(.A(new_n316), .B(new_n318), .C1(new_n319), .C2(new_n317), .ZN(new_n320));
  OR3_X1    g134(.A1(new_n320), .A2(KEYINPUT79), .A3(G110), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n316), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT24), .B(G110), .Z(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT79), .B1(new_n320), .B2(G110), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n191), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n329), .B(KEYINPUT80), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT16), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n331), .A2(new_n332), .A3(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT78), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n335));
  NAND4_X1  g149(.A1(new_n335), .A2(new_n331), .A3(new_n332), .A4(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n332), .A2(G125), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  OAI211_X1 g154(.A(new_n334), .B(new_n336), .C1(new_n340), .C2(new_n331), .ZN(new_n341));
  OR2_X1    g155(.A1(new_n341), .A2(new_n189), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n327), .A2(new_n330), .A3(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n341), .B(G146), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n320), .A2(G110), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n346), .B1(new_n322), .B2(new_n324), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n343), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n264), .A2(G221), .A3(G234), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n348), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n343), .A2(new_n347), .A3(new_n351), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n188), .A3(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT25), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n355), .A2(new_n356), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n314), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n353), .A2(new_n354), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n314), .A2(G902), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n312), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(G214), .B1(G237), .B2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G104), .ZN(new_n369));
  INV_X1    g183(.A(G104), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G107), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G101), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n370), .B2(G107), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(new_n368), .A3(G104), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n374), .A2(new_n376), .A3(new_n371), .ZN(new_n377));
  AND2_X1   g191(.A1(KEYINPUT84), .A2(G101), .ZN(new_n378));
  NOR2_X1   g192(.A1(KEYINPUT84), .A2(G101), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(KEYINPUT85), .B1(new_n377), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n374), .A2(new_n376), .A3(new_n371), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n378), .A2(new_n379), .ZN(new_n384));
  NOR3_X1   g198(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n373), .B1(new_n381), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT86), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n373), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n368), .A2(G104), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n390), .B1(KEYINPUT3), .B2(new_n369), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n391), .A2(KEYINPUT85), .A3(new_n380), .A4(new_n376), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n383), .B1(new_n382), .B2(new_n384), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n389), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT86), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT5), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n315), .A3(G116), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT89), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n315), .A3(KEYINPUT89), .A4(G116), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(G113), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(KEYINPUT5), .B2(new_n235), .ZN(new_n402));
  INV_X1    g216(.A(new_n236), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n388), .A2(new_n395), .A3(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n392), .A2(new_n393), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n382), .A2(G101), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n409), .ZN(new_n410));
  OR2_X1    g224(.A1(new_n409), .A2(KEYINPUT4), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n240), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  NAND4_X1  g226(.A1(new_n388), .A2(KEYINPUT90), .A3(new_n395), .A4(new_n404), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n407), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n415));
  XOR2_X1   g229(.A(G110), .B(G122), .Z(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT91), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n414), .A2(KEYINPUT91), .A3(new_n415), .A4(new_n416), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n258), .A2(new_n338), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n338), .B2(new_n253), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n264), .A2(G224), .ZN(new_n424));
  XNOR2_X1  g238(.A(new_n424), .B(KEYINPUT92), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n414), .A2(new_n416), .ZN(new_n427));
  INV_X1    g241(.A(new_n416), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n407), .A2(new_n428), .A3(new_n412), .A4(new_n413), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n427), .A2(KEYINPUT6), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n421), .A2(new_n426), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n424), .A2(KEYINPUT7), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n423), .B(new_n432), .ZN(new_n433));
  XOR2_X1   g247(.A(new_n401), .B(KEYINPUT94), .Z(new_n434));
  NAND2_X1  g248(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n403), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n436), .A2(new_n388), .A3(new_n395), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n437), .B1(new_n394), .B2(new_n404), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT93), .B(KEYINPUT8), .Z(new_n439));
  XNOR2_X1  g253(.A(new_n416), .B(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n433), .B1(new_n438), .B2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(G902), .B1(new_n441), .B2(new_n429), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n431), .A2(new_n442), .ZN(new_n443));
  OAI21_X1  g257(.A(G210), .B1(G237), .B2(G902), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n431), .A2(new_n444), .A3(new_n442), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n367), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  XOR2_X1   g262(.A(KEYINPUT9), .B(G234), .Z(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(G221), .B1(new_n450), .B2(G902), .ZN(new_n451));
  XNOR2_X1  g265(.A(new_n451), .B(KEYINPUT81), .ZN(new_n452));
  INV_X1    g266(.A(G469), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n188), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n388), .A2(new_n214), .A3(new_n395), .A4(KEYINPUT10), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT10), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n249), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n192), .A2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n194), .B2(new_n201), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n456), .B1(new_n459), .B2(new_n386), .ZN(new_n460));
  INV_X1    g274(.A(new_n247), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n410), .A2(new_n253), .A3(new_n411), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n455), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n264), .A2(G227), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT82), .ZN(new_n465));
  XNOR2_X1  g279(.A(G110), .B(G140), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n465), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT88), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n455), .A2(new_n460), .A3(new_n462), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n469), .B1(new_n470), .B2(new_n247), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n470), .A2(new_n469), .A3(new_n247), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT86), .B1(new_n408), .B2(new_n373), .ZN(new_n475));
  AOI211_X1 g289(.A(new_n387), .B(new_n389), .C1(new_n392), .C2(new_n393), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n258), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT87), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n459), .A2(new_n386), .ZN(new_n480));
  OAI211_X1 g294(.A(KEYINPUT87), .B(new_n258), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n482), .A2(KEYINPUT12), .A3(new_n247), .ZN(new_n483));
  AOI21_X1  g297(.A(KEYINPUT12), .B1(new_n482), .B2(new_n247), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n463), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n467), .B(KEYINPUT83), .Z(new_n486));
  INV_X1    g300(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n474), .B1(new_n485), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n454), .B1(new_n488), .B2(G469), .ZN(new_n489));
  INV_X1    g303(.A(new_n468), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n490), .B1(new_n483), .B2(new_n484), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n472), .A2(new_n473), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n467), .B1(new_n493), .B2(new_n463), .ZN(new_n494));
  OAI211_X1 g308(.A(new_n453), .B(new_n188), .C1(new_n492), .C2(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n452), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT100), .ZN(new_n497));
  AND2_X1   g311(.A1(new_n264), .A2(G952), .ZN(new_n498));
  INV_X1    g312(.A(G234), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n498), .B1(new_n499), .B2(new_n263), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g315(.A(G902), .B(G953), .C1(new_n499), .C2(new_n263), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n502), .B(KEYINPUT99), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(KEYINPUT21), .B(G898), .Z(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n501), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n370), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n330), .B1(new_n189), .B2(new_n328), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n263), .A2(new_n264), .A3(G214), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(new_n208), .ZN(new_n513));
  NAND2_X1  g327(.A1(KEYINPUT18), .A2(G131), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n513), .B(G131), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n344), .B1(new_n517), .B2(KEYINPUT17), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n513), .A2(KEYINPUT17), .A3(G131), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n519), .B(KEYINPUT96), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n510), .B(new_n516), .C1(new_n518), .C2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  XNOR2_X1  g336(.A(new_n328), .B(KEYINPUT19), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n191), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n342), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT95), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT95), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n342), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n517), .A3(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n510), .B1(new_n529), .B2(new_n516), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT20), .ZN(new_n532));
  INV_X1    g346(.A(G475), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n531), .A2(new_n532), .A3(new_n533), .A4(new_n188), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n533), .B(new_n188), .C1(new_n522), .C2(new_n530), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT20), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT97), .B(G475), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n516), .B1(new_n518), .B2(new_n520), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n510), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n538), .B1(new_n540), .B2(G902), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n204), .A2(G143), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n249), .B2(G143), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(G134), .ZN(new_n544));
  INV_X1    g358(.A(G116), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT14), .A3(G122), .ZN(new_n546));
  XNOR2_X1  g360(.A(G116), .B(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(G107), .B(new_n546), .C1(new_n548), .C2(KEYINPUT14), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n547), .A2(new_n368), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n544), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT13), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n216), .B1(new_n542), .B2(new_n552), .ZN(new_n553));
  OR2_X1    g367(.A1(new_n553), .A2(new_n543), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n547), .B(new_n368), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n543), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n554), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n450), .A2(new_n313), .A3(G953), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n551), .B2(new_n557), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT98), .B(new_n188), .C1(new_n559), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(G478), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(KEYINPUT15), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n551), .A2(new_n557), .ZN(new_n565));
  INV_X1    g379(.A(new_n558), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n551), .A2(new_n557), .A3(new_n558), .ZN(new_n568));
  AOI21_X1  g382(.A(G902), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n569), .A2(KEYINPUT98), .B1(KEYINPUT15), .B2(new_n562), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n564), .B1(new_n570), .B2(new_n561), .ZN(new_n571));
  AND4_X1   g385(.A1(new_n508), .A2(new_n537), .A3(new_n541), .A4(new_n571), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n448), .A2(new_n496), .A3(new_n497), .A4(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n431), .A2(new_n444), .A3(new_n442), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n444), .B1(new_n431), .B2(new_n442), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n572), .B(new_n366), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n452), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n493), .A2(new_n490), .ZN(new_n578));
  INV_X1    g392(.A(new_n463), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n482), .A2(new_n247), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT12), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n482), .A2(KEYINPUT12), .A3(new_n247), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n579), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  OAI211_X1 g398(.A(G469), .B(new_n578), .C1(new_n584), .C2(new_n486), .ZN(new_n585));
  INV_X1    g399(.A(new_n454), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(new_n473), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n463), .B1(new_n588), .B2(new_n471), .ZN(new_n589));
  INV_X1    g403(.A(new_n467), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI211_X1 g405(.A(G469), .B(G902), .C1(new_n591), .C2(new_n491), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n577), .B1(new_n587), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT100), .B1(new_n576), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n365), .A2(new_n573), .A3(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(new_n384), .ZN(G3));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n508), .B(new_n366), .C1(new_n574), .C2(new_n575), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n537), .A2(new_n541), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n569), .A2(new_n562), .ZN(new_n601));
  NAND2_X1  g415(.A1(G478), .A2(G902), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n603), .B1(new_n567), .B2(KEYINPUT101), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n559), .B2(new_n560), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n567), .B(new_n568), .C1(KEYINPUT101), .C2(new_n603), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g421(.A(new_n601), .B(new_n602), .C1(new_n607), .C2(new_n562), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n600), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n597), .B1(new_n598), .B2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n448), .A2(KEYINPUT102), .A3(new_n508), .A4(new_n609), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n188), .B1(new_n284), .B2(new_n290), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G472), .ZN(new_n615));
  AND2_X1   g429(.A1(new_n615), .A2(new_n291), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n593), .A2(new_n363), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n613), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XOR2_X1   g432(.A(KEYINPUT34), .B(G104), .Z(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G6));
  OR2_X1    g434(.A1(new_n599), .A2(new_n571), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n598), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n616), .A3(new_n617), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(new_n368), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G9));
  NOR2_X1   g440(.A1(new_n352), .A2(KEYINPUT36), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n348), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n361), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n359), .A2(new_n629), .ZN(new_n630));
  NAND4_X1  g444(.A1(new_n594), .A2(new_n573), .A3(new_n616), .A4(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT37), .B(G110), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G12));
  AND3_X1   g447(.A1(new_n312), .A2(new_n496), .A3(new_n630), .ZN(new_n634));
  INV_X1    g448(.A(G900), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n501), .B1(new_n504), .B2(new_n635), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n599), .A2(new_n571), .A3(new_n636), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n637), .B(new_n366), .C1(new_n575), .C2(new_n574), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT104), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n448), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n634), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G128), .ZN(G30));
  NOR2_X1   g458(.A1(new_n574), .A2(new_n575), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT38), .Z(new_n646));
  NOR3_X1   g460(.A1(new_n600), .A2(new_n571), .A3(new_n367), .ZN(new_n647));
  AND2_X1   g461(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n636), .B(KEYINPUT39), .Z(new_n649));
  NAND2_X1  g463(.A1(new_n496), .A2(new_n649), .ZN(new_n650));
  OR2_X1    g464(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n305), .A2(new_n306), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n188), .B1(new_n652), .B2(new_n288), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n287), .A2(new_n270), .ZN(new_n654));
  OAI21_X1  g468(.A(G472), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n293), .A2(new_n298), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n630), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n648), .A2(new_n651), .A3(new_n658), .A4(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT105), .B(G143), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G45));
  NOR3_X1   g476(.A1(new_n600), .A2(new_n608), .A3(new_n636), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n448), .A2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n634), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  OAI21_X1  g481(.A(new_n188), .B1(new_n494), .B2(new_n492), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G469), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n669), .A2(new_n577), .A3(new_n495), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n613), .A2(new_n365), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(KEYINPUT41), .B(G113), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G15));
  NOR3_X1   g488(.A1(new_n670), .A2(new_n645), .A3(new_n367), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n365), .A2(new_n622), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(G116), .ZN(G18));
  NAND4_X1  g491(.A1(new_n675), .A2(new_n572), .A3(new_n312), .A4(new_n630), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G119), .ZN(G21));
  NOR4_X1   g493(.A1(new_n645), .A2(new_n600), .A3(new_n571), .A4(new_n367), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n308), .A2(new_n270), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n295), .A2(new_n296), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n187), .A3(new_n188), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n615), .A2(new_n364), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n680), .A2(new_n508), .A3(new_n671), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G122), .ZN(G24));
  NAND3_X1  g500(.A1(new_n615), .A2(new_n630), .A3(new_n683), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT106), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n615), .A2(KEYINPUT106), .A3(new_n683), .A4(new_n630), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n663), .A3(new_n675), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G125), .ZN(G27));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT107), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n695), .B1(new_n587), .B2(new_n592), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n489), .A2(KEYINPUT107), .A3(new_n495), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n696), .A2(new_n577), .A3(new_n697), .ZN(new_n698));
  NOR3_X1   g512(.A1(new_n574), .A2(new_n575), .A3(new_n367), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n698), .A2(new_n312), .A3(new_n364), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n663), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n694), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n312), .A2(new_n364), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n699), .A2(new_n696), .A3(new_n577), .A4(new_n697), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n705), .A2(KEYINPUT42), .A3(new_n663), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n702), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G131), .ZN(G33));
  INV_X1    g522(.A(new_n704), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n365), .A2(new_n709), .A3(new_n637), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G134), .ZN(G36));
  OR2_X1    g525(.A1(new_n488), .A2(KEYINPUT45), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n488), .A2(KEYINPUT45), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n712), .A2(G469), .A3(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(KEYINPUT46), .A3(new_n586), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n495), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n586), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n716), .B1(KEYINPUT46), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n577), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n630), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n616), .A2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n599), .A2(new_n608), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT43), .B1(new_n599), .B2(new_n608), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT44), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n699), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n722), .A2(KEYINPUT44), .A3(new_n727), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n720), .A2(new_n649), .A3(new_n730), .A4(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G137), .ZN(G39));
  INV_X1    g547(.A(KEYINPUT47), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n719), .B(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n312), .A2(new_n364), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n735), .A2(new_n663), .A3(new_n699), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G140), .ZN(G42));
  NAND3_X1  g552(.A1(new_n725), .A2(new_n501), .A3(new_n726), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n729), .A2(new_n670), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT115), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT115), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n741), .A2(new_n742), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n691), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n742), .A2(new_n501), .A3(new_n364), .A4(new_n657), .ZN(new_n749));
  INV_X1    g563(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n600), .A3(new_n608), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n741), .A2(new_n684), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n646), .A2(new_n366), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n671), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT50), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n755), .A2(KEYINPUT114), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n755), .B2(KEYINPUT114), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n748), .B(new_n751), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n669), .A2(new_n495), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n577), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n699), .B(new_n753), .C1(new_n735), .C2(new_n762), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(KEYINPUT51), .B1(new_n760), .B2(new_n763), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n767), .B1(new_n747), .B2(new_n365), .ZN(new_n768));
  INV_X1    g582(.A(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n747), .A2(new_n767), .A3(new_n365), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(KEYINPUT48), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT48), .ZN(new_n772));
  AOI211_X1 g586(.A(KEYINPUT117), .B(new_n703), .C1(new_n744), .C2(new_n746), .ZN(new_n773));
  OAI21_X1  g587(.A(new_n772), .B1(new_n768), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n498), .B1(new_n749), .B2(new_n610), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n753), .B2(new_n675), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(KEYINPUT116), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n771), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT118), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n598), .A2(new_n610), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n616), .A3(new_n617), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n594), .A2(new_n573), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n781), .B1(new_n782), .B2(new_n703), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT108), .ZN(new_n784));
  AND2_X1   g598(.A1(new_n631), .A2(new_n623), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n595), .A2(new_n786), .A3(new_n781), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n691), .A2(new_n663), .A3(new_n709), .ZN(new_n789));
  INV_X1    g603(.A(new_n636), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n600), .A2(new_n699), .A3(new_n571), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n634), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n789), .A2(new_n710), .A3(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n788), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT42), .B1(new_n705), .B2(new_n663), .ZN(new_n795));
  NOR4_X1   g609(.A1(new_n703), .A2(new_n704), .A3(new_n694), .A4(new_n701), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n672), .A2(new_n676), .A3(new_n678), .A4(new_n685), .ZN(new_n798));
  NOR2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n634), .B1(new_n642), .B2(new_n665), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n577), .A2(new_n696), .A3(new_n790), .A4(new_n697), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n721), .A3(new_n680), .A4(new_n656), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n800), .A2(new_n692), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n800), .A2(new_n692), .A3(KEYINPUT52), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n794), .A2(KEYINPUT53), .A3(new_n799), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT111), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n789), .A2(new_n710), .A3(new_n792), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(new_n785), .A3(new_n787), .A4(new_n784), .ZN(new_n812));
  AND4_X1   g626(.A1(new_n672), .A2(new_n676), .A3(new_n678), .A4(new_n685), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n707), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n815), .A2(KEYINPUT111), .A3(KEYINPUT53), .A4(new_n807), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n810), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT110), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n805), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n803), .A2(KEYINPUT110), .A3(new_n804), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT109), .ZN(new_n821));
  AND2_X1   g635(.A1(new_n806), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n806), .A2(new_n821), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n819), .B(new_n820), .C1(new_n822), .C2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n824), .B2(new_n815), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT54), .B1(new_n817), .B2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT53), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT112), .B1(new_n797), .B2(new_n798), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT112), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n813), .A2(new_n829), .A3(new_n707), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n827), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n831), .A3(new_n794), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n794), .A2(new_n799), .ZN(new_n833));
  INV_X1    g647(.A(new_n807), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n827), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT54), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n832), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n766), .A2(new_n779), .A3(new_n826), .A4(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(G952), .B2(G953), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n723), .B1(new_n761), .B2(KEYINPUT49), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n761), .A2(KEYINPUT49), .ZN(new_n841));
  NOR4_X1   g655(.A1(new_n646), .A2(new_n656), .A3(new_n840), .A4(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n842), .A2(new_n577), .A3(new_n366), .A4(new_n364), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(G75));
  AOI21_X1  g658(.A(new_n188), .B1(new_n832), .B2(new_n835), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT56), .B1(new_n845), .B2(G210), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n421), .A2(new_n430), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n847), .B(new_n426), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n848), .B(KEYINPUT55), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n846), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n846), .A2(new_n849), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n264), .A2(G952), .ZN(new_n852));
  NOR3_X1   g666(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(G51));
  NAND2_X1  g667(.A1(new_n832), .A2(new_n835), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(KEYINPUT54), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n837), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n586), .A2(KEYINPUT57), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n586), .A2(KEYINPUT57), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n859), .B1(new_n494), .B2(new_n492), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n845), .A2(G469), .A3(new_n712), .A4(new_n713), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n852), .B1(new_n860), .B2(new_n861), .ZN(G54));
  NAND2_X1  g676(.A1(KEYINPUT58), .A2(G475), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n863), .B(KEYINPUT119), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n845), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n531), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(new_n852), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n845), .A2(new_n531), .A3(new_n864), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT120), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n867), .A2(KEYINPUT120), .A3(new_n868), .A4(new_n869), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(G60));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n826), .A2(new_n837), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n602), .B(KEYINPUT59), .Z(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n607), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n877), .B1(new_n605), .B2(new_n606), .ZN(new_n880));
  INV_X1    g694(.A(new_n837), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n836), .B1(new_n832), .B2(new_n835), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n880), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(new_n868), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n875), .B1(new_n879), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n852), .B1(new_n856), .B2(new_n880), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n877), .B1(new_n826), .B2(new_n837), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n886), .B(KEYINPUT121), .C1(new_n607), .C2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n885), .A2(new_n888), .ZN(G63));
  NAND2_X1  g703(.A1(G217), .A2(G902), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n890), .B(KEYINPUT122), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT60), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n854), .A2(new_n628), .A3(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n854), .A2(new_n892), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n360), .B(KEYINPUT123), .Z(new_n895));
  OAI211_X1 g709(.A(new_n868), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT61), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n896), .B(new_n897), .ZN(G66));
  INV_X1    g712(.A(G224), .ZN(new_n899));
  OAI21_X1  g713(.A(G953), .B1(new_n506), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n788), .A2(new_n798), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(G953), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n847), .B1(G898), .B2(new_n264), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(G69));
  XNOR2_X1  g718(.A(new_n286), .B(new_n523), .ZN(new_n905));
  NAND2_X1  g719(.A1(G900), .A2(G953), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n800), .A2(new_n692), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n732), .A2(new_n907), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(KEYINPUT125), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n720), .A2(new_n734), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n719), .A2(KEYINPUT47), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n910), .A2(new_n663), .A3(new_n699), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n736), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n707), .B(new_n710), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NAND4_X1  g729(.A1(new_n720), .A2(new_n365), .A3(new_n649), .A4(new_n680), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n909), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n905), .B(new_n906), .C1(new_n917), .C2(G953), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n905), .B(KEYINPUT124), .ZN(new_n919));
  AND2_X1   g733(.A1(new_n737), .A2(new_n732), .ZN(new_n920));
  AND2_X1   g734(.A1(new_n610), .A2(new_n621), .ZN(new_n921));
  NOR4_X1   g735(.A1(new_n703), .A2(new_n650), .A3(new_n729), .A4(new_n921), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n660), .A2(new_n907), .ZN(new_n923));
  OR2_X1    g737(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(KEYINPUT62), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n919), .B1(new_n927), .B2(G953), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n264), .B1(G227), .B2(G900), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(G72));
  NAND3_X1  g745(.A1(new_n920), .A2(new_n926), .A3(new_n901), .ZN(new_n932));
  NAND2_X1  g746(.A1(G472), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT63), .Z(new_n934));
  NAND2_X1  g748(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n852), .B1(new_n935), .B2(new_n654), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n909), .A2(new_n915), .A3(new_n901), .A4(new_n916), .ZN(new_n937));
  AND2_X1   g751(.A1(new_n937), .A2(new_n934), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n299), .B(KEYINPUT126), .Z(new_n939));
  OAI21_X1  g753(.A(new_n936), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n299), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n941), .A2(new_n654), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n934), .B(new_n942), .C1(new_n817), .C2(new_n825), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n944));
  OR2_X1    g758(.A1(new_n943), .A2(KEYINPUT127), .ZN(new_n945));
  AOI21_X1  g759(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G57));
endmodule


