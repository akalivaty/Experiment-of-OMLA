//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 0 0 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1354, new_n1355, new_n1356, new_n1357, new_n1358, new_n1359,
    new_n1360, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  OAI21_X1  g0004(.A(G50), .B1(G58), .B2(G68), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NAND2_X1  g0006(.A1(G1), .A2(G13), .ZN(new_n207));
  NOR3_X1   g0007(.A1(new_n205), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(new_n206), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT0), .ZN(new_n214));
  AOI21_X1  g0014(.A(new_n208), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n202), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n211), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n215), .B1(new_n214), .B2(new_n213), .C1(new_n224), .C2(KEYINPUT1), .ZN(new_n225));
  AOI21_X1  g0025(.A(new_n225), .B1(KEYINPUT1), .B2(new_n224), .ZN(G361));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n227), .B(KEYINPUT2), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G226), .ZN(new_n229));
  XOR2_X1   g0029(.A(KEYINPUT64), .B(G232), .Z(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT65), .Z(new_n232));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XNOR2_X1  g0037(.A(G50), .B(G58), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G33), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n206), .A2(new_n244), .A3(KEYINPUT67), .ZN(new_n245));
  INV_X1    g0045(.A(KEYINPUT67), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G20), .B2(G33), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G150), .ZN(new_n249));
  XNOR2_X1  g0049(.A(KEYINPUT8), .B(G58), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT66), .ZN(new_n251));
  OAI21_X1  g0051(.A(new_n251), .B1(new_n244), .B2(G20), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n206), .A2(KEYINPUT66), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI221_X1 g0054(.A(new_n249), .B1(new_n206), .B2(new_n201), .C1(new_n250), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n207), .ZN(new_n257));
  AND2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(new_n217), .ZN(new_n261));
  INV_X1    g0061(.A(new_n257), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(new_n259), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n209), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(G50), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n261), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n258), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G41), .ZN(new_n268));
  INV_X1    g0068(.A(G45), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(G274), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n207), .B1(G33), .B2(G41), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n270), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n271), .B1(new_n274), .B2(new_n218), .ZN(new_n275));
  AND2_X1   g0075(.A1(KEYINPUT3), .A2(G33), .ZN(new_n276));
  NOR2_X1   g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n278), .A2(G1698), .ZN(new_n279));
  AOI22_X1  g0079(.A1(new_n279), .A2(G222), .B1(G77), .B2(new_n278), .ZN(new_n280));
  INV_X1    g0080(.A(G223), .ZN(new_n281));
  OR2_X1    g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND2_X1  g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G1698), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n280), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n275), .B1(new_n286), .B2(new_n272), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G169), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n287), .A2(G179), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n267), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(new_n258), .A2(new_n266), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT9), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(new_n293), .B1(new_n287), .B2(G190), .ZN(new_n294));
  AOI22_X1  g0094(.A1(new_n288), .A2(G200), .B1(new_n267), .B2(KEYINPUT9), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n288), .A2(G200), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT70), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n297), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OR2_X1    g0100(.A1(new_n296), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n296), .A2(new_n300), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n291), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G238), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n271), .B1(new_n274), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n279), .A2(G226), .ZN(new_n306));
  NAND2_X1  g0106(.A1(G33), .A2(G97), .ZN(new_n307));
  INV_X1    g0107(.A(G232), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n306), .B(new_n307), .C1(new_n308), .C2(new_n285), .ZN(new_n309));
  AOI211_X1 g0109(.A(KEYINPUT13), .B(new_n305), .C1(new_n309), .C2(new_n272), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n309), .A2(new_n272), .ZN(new_n312));
  INV_X1    g0112(.A(new_n305), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n311), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(G169), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT14), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(new_n310), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT71), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n305), .B1(new_n309), .B2(new_n272), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n319), .B1(new_n320), .B2(new_n311), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n317), .A2(new_n318), .A3(G179), .A4(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT14), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n323), .B(G169), .C1(new_n310), .C2(new_n314), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n245), .A2(new_n247), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(new_n217), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n254), .A2(new_n202), .B1(new_n206), .B2(G68), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n257), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g0129(.A(KEYINPUT73), .B(KEYINPUT11), .Z(new_n330));
  XNOR2_X1  g0130(.A(new_n329), .B(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n263), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(G68), .A3(new_n264), .ZN(new_n333));
  INV_X1    g0133(.A(G13), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n334), .A2(G1), .ZN(new_n335));
  INV_X1    g0135(.A(G68), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(G20), .A3(new_n336), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n337), .A2(KEYINPUT74), .A3(KEYINPUT12), .ZN(new_n338));
  OAI21_X1  g0138(.A(KEYINPUT74), .B1(new_n337), .B2(KEYINPUT12), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n337), .A2(KEYINPUT12), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(new_n331), .B(new_n333), .C1(new_n338), .C2(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n325), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G190), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n344), .B1(new_n320), .B2(new_n311), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n317), .A2(new_n321), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(KEYINPUT72), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT72), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n317), .A2(new_n348), .A3(new_n321), .A4(new_n345), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  OR2_X1    g0150(.A1(new_n310), .A2(new_n314), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n342), .B1(new_n351), .B2(G200), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n326), .A2(new_n250), .B1(new_n206), .B2(new_n202), .ZN(new_n354));
  XNOR2_X1  g0154(.A(KEYINPUT15), .B(G87), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n254), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n257), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT68), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n264), .A2(G77), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT69), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n260), .B2(new_n202), .ZN(new_n361));
  NOR3_X1   g0161(.A1(new_n259), .A2(KEYINPUT69), .A3(G77), .ZN(new_n362));
  OAI221_X1 g0162(.A(new_n358), .B1(new_n263), .B2(new_n359), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  AOI22_X1  g0163(.A1(new_n279), .A2(G232), .B1(G107), .B2(new_n278), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n304), .B2(new_n285), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n272), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n273), .A2(G244), .B1(G274), .B2(new_n270), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G169), .ZN(new_n369));
  INV_X1    g0169(.A(G179), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n369), .B1(new_n370), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n363), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n368), .A2(G190), .ZN(new_n374));
  INV_X1    g0174(.A(G200), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n374), .B1(new_n375), .B2(new_n368), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(new_n363), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n303), .A2(new_n343), .A3(new_n353), .A4(new_n378), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n250), .B1(new_n209), .B2(G20), .ZN(new_n380));
  AOI22_X1  g0180(.A1(new_n332), .A2(new_n380), .B1(new_n260), .B2(new_n250), .ZN(new_n381));
  NOR3_X1   g0181(.A1(new_n276), .A2(new_n277), .A3(G20), .ZN(new_n382));
  OAI21_X1  g0182(.A(KEYINPUT75), .B1(new_n382), .B2(KEYINPUT7), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n282), .A2(new_n206), .A3(new_n283), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT75), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT7), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n278), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n248), .A2(G159), .ZN(new_n391));
  INV_X1    g0191(.A(G58), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n336), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  OAI21_X1  g0194(.A(G20), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n391), .A2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(KEYINPUT16), .B1(new_n390), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n384), .A2(new_n386), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n388), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(G68), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(KEYINPUT16), .A3(new_n397), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(new_n257), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n381), .B1(new_n398), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G41), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(G1), .A3(G13), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(G232), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n271), .ZN(new_n409));
  INV_X1    g0209(.A(G1698), .ZN(new_n410));
  OAI211_X1 g0210(.A(G223), .B(new_n410), .C1(new_n276), .C2(new_n277), .ZN(new_n411));
  OAI211_X1 g0211(.A(G226), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n412));
  NAND2_X1  g0212(.A1(G33), .A2(G87), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  AOI211_X1 g0214(.A(G179), .B(new_n409), .C1(new_n272), .C2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n272), .ZN(new_n416));
  INV_X1    g0216(.A(new_n409), .ZN(new_n417));
  AOI21_X1  g0217(.A(G169), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(KEYINPUT76), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g0219(.A1(new_n416), .A2(new_n370), .A3(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT76), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n409), .B1(new_n414), .B2(new_n272), .ZN(new_n422));
  OAI211_X1 g0222(.A(new_n420), .B(new_n421), .C1(G169), .C2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n404), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT18), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n425), .A2(KEYINPUT77), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT77), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n396), .B1(new_n389), .B2(G68), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n257), .B(new_n402), .C1(new_n429), .C2(KEYINPUT16), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n381), .B1(new_n419), .B2(new_n423), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n431), .B2(KEYINPUT18), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT17), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT78), .ZN(new_n436));
  AND3_X1   g0236(.A1(new_n422), .A2(new_n436), .A3(new_n344), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n422), .A2(new_n344), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n436), .B1(new_n422), .B2(G200), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n435), .B1(new_n404), .B2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n381), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT16), .ZN(new_n443));
  NOR4_X1   g0243(.A1(new_n276), .A2(new_n277), .A3(new_n386), .A4(G20), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n444), .B1(KEYINPUT75), .B2(new_n399), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n336), .B1(new_n445), .B2(new_n387), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n443), .B1(new_n446), .B2(new_n396), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n396), .B1(G68), .B2(new_n400), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n262), .B1(new_n448), .B2(KEYINPUT16), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n442), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n437), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n439), .A2(new_n438), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n450), .A2(KEYINPUT17), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(KEYINPUT79), .B1(new_n441), .B2(new_n454), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n441), .A2(new_n454), .A3(KEYINPUT79), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n434), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(new_n269), .A2(G1), .ZN(new_n458));
  AND2_X1   g0258(.A1(KEYINPUT5), .A2(G41), .ZN(new_n459));
  NOR2_X1   g0259(.A1(KEYINPUT5), .A2(G41), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n461), .A2(G270), .A3(new_n406), .ZN(new_n462));
  OR2_X1    g0262(.A1(KEYINPUT5), .A2(G41), .ZN(new_n463));
  NAND2_X1  g0263(.A1(KEYINPUT5), .A2(G41), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n465), .A2(G274), .A3(new_n458), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  OAI211_X1 g0267(.A(G264), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n468));
  OAI211_X1 g0268(.A(G257), .B(new_n410), .C1(new_n276), .C2(new_n277), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n282), .A2(G303), .A3(new_n283), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n272), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n467), .A2(new_n344), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n462), .A2(new_n466), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(new_n272), .B2(new_n471), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n475), .B2(G200), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT20), .ZN(new_n477));
  INV_X1    g0277(.A(G116), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n206), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  INV_X1    g0280(.A(G97), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(G33), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n479), .B1(new_n482), .B2(new_n206), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n477), .B1(new_n483), .B2(new_n262), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n244), .A2(G97), .ZN(new_n485));
  AOI21_X1  g0285(.A(G20), .B1(new_n485), .B2(new_n480), .ZN(new_n486));
  OAI211_X1 g0286(.A(KEYINPUT20), .B(new_n257), .C1(new_n486), .C2(new_n479), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT84), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n259), .A2(new_n478), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n209), .A2(G33), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n259), .A2(new_n491), .A3(new_n207), .A4(new_n256), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n490), .B1(new_n493), .B2(new_n478), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n488), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n488), .A2(new_n494), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT84), .ZN(new_n497));
  AND3_X1   g0297(.A1(new_n476), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n475), .A2(G179), .ZN(new_n499));
  INV_X1    g0299(.A(G169), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n500), .B1(new_n467), .B2(new_n472), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT21), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n499), .A2(new_n502), .B1(new_n497), .B2(new_n495), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n467), .A2(new_n472), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G169), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(new_n497), .B2(new_n495), .ZN(new_n506));
  OAI21_X1  g0306(.A(KEYINPUT85), .B1(new_n506), .B2(KEYINPUT21), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n488), .A2(new_n489), .A3(new_n494), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n489), .B1(new_n488), .B2(new_n494), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n501), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT85), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT21), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n510), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n498), .B(new_n503), .C1(new_n507), .C2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n272), .B1(new_n458), .B2(new_n465), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(G264), .ZN(new_n516));
  INV_X1    g0316(.A(G294), .ZN(new_n517));
  NOR2_X1   g0317(.A1(new_n244), .A2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G257), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n282), .B2(new_n283), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n518), .B1(new_n520), .B2(G1698), .ZN(new_n521));
  OAI211_X1 g0321(.A(G250), .B(new_n410), .C1(new_n276), .C2(new_n277), .ZN(new_n522));
  AOI21_X1  g0322(.A(KEYINPUT86), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g0323(.A(G257), .B(G1698), .C1(new_n276), .C2(new_n277), .ZN(new_n524));
  INV_X1    g0324(.A(new_n518), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n522), .A2(new_n524), .A3(KEYINPUT86), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n272), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n516), .B(new_n466), .C1(new_n523), .C2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n375), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT86), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n532), .A2(new_n272), .A3(new_n526), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n533), .A2(new_n344), .A3(new_n516), .A4(new_n466), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n529), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(G107), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n335), .A2(G20), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n537), .B(KEYINPUT25), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n538), .B1(G107), .B2(new_n493), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT23), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n540), .B1(new_n206), .B2(G107), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n536), .A2(KEYINPUT23), .A3(G20), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n244), .A2(new_n478), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n544), .A2(new_n206), .ZN(new_n545));
  AND2_X1   g0345(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n206), .B(G87), .C1(new_n276), .C2(new_n277), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n549));
  OAI211_X1 g0349(.A(KEYINPUT24), .B(new_n546), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n257), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n543), .A2(new_n545), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(KEYINPUT22), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT22), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n284), .A2(new_n554), .A3(new_n206), .A4(G87), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n552), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(KEYINPUT24), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n539), .B1(new_n551), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n535), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n528), .A2(G169), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n533), .A2(G179), .A3(new_n516), .A4(new_n466), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n558), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n560), .A2(new_n564), .A3(KEYINPUT87), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT87), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n558), .B1(new_n529), .B2(new_n534), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n262), .B1(new_n556), .B2(KEYINPUT24), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT24), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n561), .A2(new_n562), .B1(new_n572), .B2(new_n539), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n566), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n565), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT82), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT81), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT6), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n577), .A2(new_n578), .B1(new_n481), .B2(G107), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n536), .A2(G97), .ZN(new_n580));
  NAND2_X1  g0380(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n579), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(new_n581), .ZN(new_n583));
  NOR2_X1   g0383(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n584));
  OAI211_X1 g0384(.A(G97), .B(new_n536), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n206), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(KEYINPUT80), .B1(new_n248), .B2(G77), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT80), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n588), .B(new_n202), .C1(new_n245), .C2(new_n247), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n389), .A2(G107), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n262), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n259), .A2(G97), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n593), .B1(new_n493), .B2(G97), .ZN(new_n594));
  INV_X1    g0394(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n576), .B1(new_n592), .B2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT4), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(G1698), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n284), .A2(G244), .A3(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n219), .B1(new_n282), .B2(new_n283), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n599), .B(new_n480), .C1(KEYINPUT4), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n284), .A2(G250), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n410), .B1(new_n602), .B2(KEYINPUT4), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n272), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n515), .A2(G257), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n605), .A2(new_n466), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n604), .A2(new_n606), .A3(new_n344), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n605), .A2(new_n466), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n602), .A2(KEYINPUT4), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(G1698), .ZN(new_n610));
  INV_X1    g0410(.A(new_n600), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n611), .A2(new_n597), .B1(G33), .B2(G283), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n612), .A3(new_n599), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n608), .B1(new_n613), .B2(new_n272), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n607), .B1(new_n614), .B2(G200), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n536), .B1(new_n445), .B2(new_n387), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n587), .A2(new_n589), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n582), .A2(new_n585), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(G20), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n257), .B1(new_n616), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n621), .A2(KEYINPUT82), .A3(new_n594), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n596), .A2(new_n615), .A3(new_n622), .ZN(new_n623));
  AOI21_X1  g0423(.A(G169), .B1(new_n604), .B2(new_n606), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n624), .B1(new_n370), .B2(new_n614), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n621), .A2(new_n594), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n355), .A2(new_n260), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT19), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n254), .B2(new_n481), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n284), .A2(new_n206), .A3(G68), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n206), .B1(new_n307), .B2(new_n629), .ZN(new_n632));
  OR2_X1    g0432(.A1(G87), .A2(G97), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n632), .B1(G107), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n630), .A2(new_n631), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n628), .B1(new_n635), .B2(new_n257), .ZN(new_n636));
  XNOR2_X1  g0436(.A(new_n355), .B(KEYINPUT83), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n493), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(G250), .B1(new_n269), .B2(G1), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n458), .A2(G274), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n272), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n284), .A2(G238), .A3(new_n410), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n284), .A2(G244), .A3(G1698), .ZN(new_n645));
  INV_X1    g0445(.A(new_n544), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  AOI211_X1 g0447(.A(G179), .B(new_n643), .C1(new_n647), .C2(new_n272), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n643), .B1(new_n647), .B2(new_n272), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n648), .B1(new_n500), .B2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n649), .A2(new_n375), .ZN(new_n652));
  AOI211_X1 g0452(.A(new_n344), .B(new_n643), .C1(new_n647), .C2(new_n272), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n493), .A2(G87), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n636), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n640), .A2(new_n651), .B1(new_n654), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n623), .A2(new_n627), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n514), .A2(new_n575), .A3(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n379), .A2(new_n457), .A3(new_n660), .ZN(G372));
  NAND2_X1  g0461(.A1(new_n353), .A2(new_n373), .ZN(new_n662));
  INV_X1    g0462(.A(KEYINPUT79), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n404), .A2(new_n440), .A3(new_n435), .ZN(new_n664));
  AOI21_X1  g0464(.A(KEYINPUT17), .B1(new_n450), .B2(new_n453), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n441), .A2(new_n454), .A3(KEYINPUT79), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n662), .A2(new_n343), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n415), .A2(new_n418), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  XOR2_X1   g0471(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n672));
  NOR3_X1   g0472(.A1(new_n450), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n672), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n404), .B2(new_n670), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  OR3_X1    g0476(.A1(new_n668), .A2(new_n669), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n301), .A2(new_n302), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n669), .B1(new_n668), .B2(new_n676), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n291), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n379), .A2(new_n457), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n651), .A2(new_n640), .ZN(new_n683));
  INV_X1    g0483(.A(new_n652), .ZN(new_n684));
  INV_X1    g0484(.A(new_n653), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n657), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n683), .A2(new_n625), .A3(new_n686), .A4(new_n626), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n649), .A2(new_n370), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n688), .B(KEYINPUT88), .C1(G169), .C2(new_n649), .ZN(new_n689));
  AND2_X1   g0489(.A1(new_n636), .A2(new_n639), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n688), .B1(G169), .B2(new_n649), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT88), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n690), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AOI22_X1  g0493(.A1(new_n687), .A2(KEYINPUT26), .B1(new_n689), .B2(new_n693), .ZN(new_n694));
  NOR3_X1   g0494(.A1(new_n656), .A2(new_n652), .A3(new_n653), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n695), .B1(new_n693), .B2(new_n689), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT26), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n596), .A2(new_n622), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n625), .A4(new_n698), .ZN(new_n699));
  AND2_X1   g0499(.A1(new_n694), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n503), .B1(new_n507), .B2(new_n513), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n564), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n691), .A2(new_n692), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n703), .A2(new_n640), .A3(new_n689), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n686), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n567), .ZN(new_n706));
  AND2_X1   g0506(.A1(new_n623), .A2(new_n627), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n682), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n680), .A2(new_n681), .A3(new_n710), .ZN(G369));
  NAND2_X1  g0511(.A1(new_n335), .A2(new_n206), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(KEYINPUT27), .ZN(new_n713));
  XNOR2_X1  g0513(.A(new_n713), .B(KEYINPUT91), .ZN(new_n714));
  INV_X1    g0514(.A(G213), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n715), .B1(new_n712), .B2(KEYINPUT27), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(G343), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n720), .B1(new_n495), .B2(new_n497), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n514), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n722), .B1(new_n701), .B2(new_n721), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  AOI22_X1  g0524(.A1(new_n565), .A2(new_n574), .B1(new_n558), .B2(new_n719), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n573), .B2(new_n719), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n701), .A2(new_n719), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n725), .A2(new_n729), .B1(new_n573), .B2(new_n720), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n728), .A2(new_n730), .ZN(G399));
  INV_X1    g0531(.A(new_n212), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(G41), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n633), .A2(G107), .A3(G116), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n734), .A2(G1), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(new_n205), .B2(new_n734), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT28), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n698), .A2(new_n625), .ZN(new_n739));
  OAI21_X1  g0539(.A(KEYINPUT26), .B1(new_n705), .B2(new_n739), .ZN(new_n740));
  OR2_X1    g0540(.A1(new_n687), .A2(KEYINPUT26), .ZN(new_n741));
  AND3_X1   g0541(.A1(new_n740), .A2(new_n741), .A3(new_n704), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n719), .B1(new_n742), .B2(new_n708), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n719), .B1(new_n700), .B2(new_n708), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(KEYINPUT29), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n660), .A2(KEYINPUT31), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n604), .A2(new_n606), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n533), .A2(new_n516), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n748), .A2(new_n749), .A3(new_n650), .ZN(new_n750));
  INV_X1    g0550(.A(KEYINPUT92), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(new_n504), .B2(new_n370), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n475), .A2(KEYINPUT92), .A3(G179), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n750), .A2(new_n754), .A3(KEYINPUT30), .ZN(new_n755));
  NOR3_X1   g0555(.A1(new_n475), .A2(new_n649), .A3(G179), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n756), .A2(new_n528), .A3(new_n748), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(KEYINPUT30), .B1(new_n750), .B2(new_n754), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT31), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n720), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n747), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT93), .ZN(new_n765));
  INV_X1    g0565(.A(new_n760), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n720), .A2(new_n761), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n766), .A2(new_n765), .A3(new_n767), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n764), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G330), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n746), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n738), .B1(new_n773), .B2(G1), .ZN(G364));
  NOR2_X1   g0574(.A1(new_n206), .A2(new_n344), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n370), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n206), .A2(G190), .ZN(new_n779));
  NOR2_X1   g0579(.A1(G179), .A2(G200), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G322), .A2(new_n778), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G283), .ZN(new_n784));
  INV_X1    g0584(.A(new_n779), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(G179), .A3(new_n375), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n783), .B1(new_n784), .B2(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n370), .A2(new_n375), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n775), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n776), .A2(new_n779), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n791), .A2(G326), .B1(new_n793), .B2(G311), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n789), .A2(new_n779), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g0596(.A(KEYINPUT33), .B(G317), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n284), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n206), .B1(new_n780), .B2(G190), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n794), .B(new_n798), .C1(new_n517), .C2(new_n799), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n775), .A2(new_n370), .A3(G200), .ZN(new_n801));
  OR2_X1    g0601(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(KEYINPUT96), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n788), .B(new_n800), .C1(G303), .C2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT98), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n787), .A2(new_n536), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n284), .B1(new_n777), .B2(new_n392), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n795), .A2(new_n336), .B1(new_n792), .B2(new_n202), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n790), .A2(new_n217), .ZN(new_n811));
  NOR4_X1   g0611(.A1(new_n808), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n805), .A2(G87), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n799), .B(KEYINPUT97), .Z(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(G97), .ZN(new_n815));
  XNOR2_X1  g0615(.A(KEYINPUT95), .B(G159), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n781), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT32), .ZN(new_n818));
  NAND4_X1  g0618(.A1(new_n812), .A2(new_n813), .A3(new_n815), .A4(new_n818), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n807), .A2(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n207), .B1(G20), .B2(new_n500), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n334), .A2(G20), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G45), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n734), .A2(G1), .A3(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n732), .A2(new_n278), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n828), .A2(G355), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n829), .B1(G116), .B2(new_n212), .ZN(new_n830));
  MUX2_X1   g0630(.A(new_n205), .B(new_n239), .S(G45), .Z(new_n831));
  NOR2_X1   g0631(.A1(new_n732), .A2(new_n284), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(G13), .A2(G33), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n835), .A2(G20), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n836), .A2(new_n821), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n827), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n823), .B1(KEYINPUT94), .B2(new_n839), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n840), .B1(KEYINPUT94), .B2(new_n839), .ZN(new_n841));
  INV_X1    g0641(.A(new_n836), .ZN(new_n842));
  NOR2_X1   g0642(.A1(new_n723), .A2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n724), .A2(new_n826), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n723), .A2(G330), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n841), .A2(new_n843), .B1(new_n844), .B2(new_n845), .ZN(G396));
  NOR2_X1   g0646(.A1(new_n821), .A2(new_n834), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n826), .B1(new_n202), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n805), .A2(G107), .ZN(new_n849));
  INV_X1    g0649(.A(G303), .ZN(new_n850));
  INV_X1    g0650(.A(G311), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n790), .A2(new_n850), .B1(new_n781), .B2(new_n851), .ZN(new_n852));
  AOI211_X1 g0652(.A(new_n284), .B(new_n852), .C1(G87), .C2(new_n786), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n784), .A2(new_n795), .B1(new_n777), .B2(new_n517), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n854), .B1(G116), .B2(new_n793), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n849), .A2(new_n853), .A3(new_n815), .A4(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(new_n816), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n791), .A2(G137), .B1(new_n793), .B2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(G143), .ZN(new_n859));
  INV_X1    g0659(.A(G150), .ZN(new_n860));
  OAI221_X1 g0660(.A(new_n858), .B1(new_n859), .B2(new_n777), .C1(new_n860), .C2(new_n795), .ZN(new_n861));
  XOR2_X1   g0661(.A(new_n861), .B(KEYINPUT34), .Z(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n284), .B1(new_n781), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(new_n864), .B1(G68), .B2(new_n786), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n865), .B1(new_n392), .B2(new_n799), .C1(new_n804), .C2(new_n217), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n856), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT99), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n821), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n867), .A2(new_n868), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n372), .A2(new_n719), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n363), .A2(new_n719), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n872), .B1(new_n376), .B2(new_n363), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n871), .B1(new_n873), .B2(new_n372), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n848), .B1(new_n869), .B2(new_n870), .C1(new_n874), .C2(new_n835), .ZN(new_n875));
  INV_X1    g0675(.A(new_n772), .ZN(new_n876));
  INV_X1    g0676(.A(new_n874), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n745), .B(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n827), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n876), .A2(new_n878), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n875), .B1(new_n880), .B2(new_n881), .ZN(G384));
  NOR3_X1   g0682(.A1(new_n207), .A2(new_n206), .A3(new_n478), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n883), .B1(new_n618), .B2(KEYINPUT35), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(KEYINPUT35), .B2(new_n618), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n885), .B(KEYINPUT36), .ZN(new_n886));
  NOR3_X1   g0686(.A1(new_n393), .A2(new_n205), .A3(new_n202), .ZN(new_n887));
  OR2_X1    g0687(.A1(new_n887), .A2(KEYINPUT100), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(KEYINPUT100), .B1(new_n217), .B2(G68), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n209), .B(G13), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n886), .A2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n449), .B1(KEYINPUT16), .B2(new_n448), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n381), .ZN(new_n895));
  INV_X1    g0695(.A(new_n717), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n666), .A2(new_n667), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n898), .B2(new_n434), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n431), .A2(KEYINPUT37), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n404), .A2(new_n440), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n404), .A2(new_n896), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  AOI22_X1  g0704(.A1(new_n894), .A2(new_n381), .B1(new_n671), .B2(new_n717), .ZN(new_n905));
  OAI21_X1  g0705(.A(KEYINPUT37), .B1(new_n905), .B2(new_n901), .ZN(new_n906));
  AND2_X1   g0706(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n893), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n906), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n404), .A2(new_n424), .A3(KEYINPUT18), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT77), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n425), .A2(new_n426), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n666), .A2(new_n667), .B1(new_n913), .B2(new_n427), .ZN(new_n914));
  OAI211_X1 g0714(.A(KEYINPUT38), .B(new_n909), .C1(new_n914), .C2(new_n897), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n908), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n342), .A2(new_n719), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n353), .A2(new_n343), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n325), .A2(new_n342), .A3(new_n719), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n762), .B1(new_n660), .B2(KEYINPUT31), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n766), .A2(new_n767), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n920), .B(new_n874), .C1(new_n921), .C2(new_n923), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n892), .B1(new_n916), .B2(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n924), .ZN(new_n926));
  AOI22_X1  g0726(.A1(new_n671), .A2(new_n717), .B1(new_n430), .B2(new_n381), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT102), .B1(new_n404), .B2(new_n440), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT102), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n450), .A2(new_n929), .A3(new_n453), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n927), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT37), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n904), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n441), .A2(new_n454), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n404), .B(new_n896), .C1(new_n676), .C2(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n893), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n892), .B1(new_n915), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n926), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n925), .A2(G330), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n764), .A2(new_n922), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n682), .A2(G330), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n943), .A2(KEYINPUT103), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(KEYINPUT103), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n908), .A2(new_n915), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n877), .B1(new_n764), .B2(new_n922), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n946), .A2(new_n947), .A3(new_n920), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n948), .A2(new_n892), .B1(new_n926), .B2(new_n938), .ZN(new_n949));
  NAND3_X1  g0749(.A1(new_n949), .A2(new_n682), .A3(new_n941), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n918), .A2(new_n919), .ZN(new_n952));
  AND3_X1   g0752(.A1(new_n702), .A2(new_n706), .A3(new_n707), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n694), .A2(new_n699), .ZN(new_n954));
  OAI211_X1 g0754(.A(new_n720), .B(new_n874), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  INV_X1    g0755(.A(new_n871), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n952), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n957), .A2(new_n946), .ZN(new_n958));
  INV_X1    g0758(.A(new_n676), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n958), .B1(new_n959), .B2(new_n896), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n343), .A2(new_n719), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n946), .A2(KEYINPUT101), .A3(KEYINPUT39), .ZN(new_n962));
  INV_X1    g0762(.A(KEYINPUT101), .ZN(new_n963));
  AOI21_X1  g0763(.A(KEYINPUT38), .B1(new_n933), .B2(new_n935), .ZN(new_n964));
  INV_X1    g0764(.A(new_n897), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n907), .B1(new_n457), .B2(new_n965), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n966), .B2(KEYINPUT38), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT39), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n968), .B1(new_n908), .B2(new_n915), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n962), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n960), .B1(new_n961), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n680), .A2(new_n681), .ZN(new_n973));
  OAI211_X1 g0773(.A(new_n744), .B(new_n682), .C1(KEYINPUT29), .C2(new_n745), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n972), .B(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n951), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n978), .B1(new_n209), .B2(new_n824), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n951), .A2(new_n977), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n891), .B1(new_n979), .B2(new_n980), .ZN(G367));
  NAND2_X1  g0781(.A1(new_n698), .A2(new_n719), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n707), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n698), .A2(new_n625), .A3(new_n719), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n985), .A2(new_n573), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n719), .B1(new_n986), .B2(new_n627), .ZN(new_n987));
  INV_X1    g0787(.A(new_n985), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n725), .A2(new_n729), .ZN(new_n989));
  NOR3_X1   g0789(.A1(new_n988), .A2(KEYINPUT42), .A3(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n987), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(KEYINPUT42), .B1(new_n988), .B2(new_n989), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n720), .A2(new_n657), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n696), .A2(new_n993), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n704), .A2(new_n993), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n991), .A2(new_n992), .B1(KEYINPUT43), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n996), .A2(KEYINPUT43), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n728), .A2(new_n988), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n733), .B(KEYINPUT41), .Z(new_n1002));
  NAND2_X1  g0802(.A1(new_n730), .A2(new_n985), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n1003), .A2(KEYINPUT104), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(KEYINPUT104), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT45), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1004), .A2(KEYINPUT45), .A3(new_n1005), .ZN(new_n1008));
  NOR2_X1   g0808(.A1(new_n730), .A2(new_n985), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT44), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1011), .A2(new_n727), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n726), .B1(new_n701), .B2(new_n719), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n989), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n724), .ZN(new_n1015));
  XOR2_X1   g0815(.A(new_n1015), .B(KEYINPUT105), .Z(new_n1016));
  NAND2_X1  g0816(.A1(new_n1014), .A2(new_n724), .ZN(new_n1017));
  AND3_X1   g0817(.A1(new_n1016), .A2(new_n773), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1011), .A2(new_n727), .ZN(new_n1019));
  NAND3_X1  g0819(.A1(new_n1012), .A2(new_n1018), .A3(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1002), .B1(new_n1020), .B2(new_n773), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n825), .A2(G1), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1001), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n832), .A2(new_n235), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n837), .B1(new_n212), .B2(new_n355), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n278), .B1(new_n795), .B2(new_n517), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n787), .A2(new_n481), .B1(new_n851), .B2(new_n790), .ZN(new_n1027));
  INV_X1    g0827(.A(new_n799), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1026), .B(new_n1027), .C1(G107), .C2(new_n1028), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n777), .A2(new_n850), .B1(new_n792), .B2(new_n784), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(G317), .B2(new_n782), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT46), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n804), .B2(new_n478), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n805), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1029), .A2(new_n1031), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  XOR2_X1   g0835(.A(KEYINPUT107), .B(G137), .Z(new_n1036));
  OAI22_X1  g0836(.A1(new_n1036), .A2(new_n781), .B1(new_n777), .B2(new_n860), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n786), .A2(G77), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n284), .ZN(new_n1039));
  AOI211_X1 g0839(.A(new_n1037), .B(new_n1039), .C1(G143), .C2(new_n791), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n796), .A2(new_n857), .B1(new_n793), .B2(G50), .ZN(new_n1041));
  OR2_X1    g0841(.A1(new_n1041), .A2(KEYINPUT106), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n805), .A2(G58), .B1(new_n1041), .B2(KEYINPUT106), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n814), .A2(G68), .ZN(new_n1044));
  NAND4_X1  g0844(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1035), .A2(KEYINPUT47), .A3(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1046), .A2(new_n821), .ZN(new_n1047));
  AOI21_X1  g0847(.A(KEYINPUT47), .B1(new_n1035), .B2(new_n1045), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n827), .B1(new_n1024), .B2(new_n1025), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT108), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1050), .B1(new_n842), .B2(new_n996), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1023), .A2(new_n1051), .ZN(G387));
  OAI21_X1  g0852(.A(new_n278), .B1(new_n787), .B2(new_n478), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n805), .A2(G294), .B1(G283), .B2(new_n1028), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT48), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n791), .A2(G322), .B1(new_n793), .B2(G303), .ZN(new_n1056));
  INV_X1    g0856(.A(G317), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1056), .B1(new_n851), .B2(new_n795), .C1(new_n1057), .C2(new_n777), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1054), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT49), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n1053), .B(new_n1061), .C1(G326), .C2(new_n782), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n638), .A2(new_n814), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n217), .A2(new_n777), .B1(new_n795), .B2(new_n250), .ZN(new_n1064));
  AOI211_X1 g0864(.A(new_n278), .B(new_n1064), .C1(G97), .C2(new_n786), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n805), .A2(G77), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n792), .A2(new_n336), .B1(new_n781), .B2(new_n860), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G159), .B2(new_n791), .ZN(new_n1068));
  AND4_X1   g0868(.A1(new_n1063), .A2(new_n1065), .A3(new_n1066), .A4(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n821), .B1(new_n1062), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n735), .ZN(new_n1071));
  AOI22_X1  g0871(.A1(new_n828), .A2(new_n1071), .B1(new_n536), .B2(new_n732), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n231), .A2(new_n269), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n250), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n217), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n1075), .B(KEYINPUT50), .ZN(new_n1076));
  OR2_X1    g0876(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n735), .A2(KEYINPUT109), .ZN(new_n1078));
  AOI21_X1  g0878(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n832), .B1(new_n1076), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1072), .B1(new_n1073), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n826), .B1(new_n1082), .B2(new_n837), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1070), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n726), .B2(new_n836), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1085), .B1(new_n1086), .B2(new_n1022), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1018), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n733), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n1086), .A2(new_n773), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(G393));
  INV_X1    g0891(.A(KEYINPUT113), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n988), .A2(new_n836), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT111), .ZN(new_n1094));
  AOI211_X1 g0894(.A(new_n284), .B(new_n808), .C1(G116), .C2(new_n1028), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n790), .A2(new_n1057), .B1(new_n777), .B2(new_n851), .ZN(new_n1096));
  XNOR2_X1  g0896(.A(new_n1096), .B(KEYINPUT52), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n805), .A2(G283), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n795), .A2(new_n850), .B1(new_n792), .B2(new_n517), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G322), .B2(new_n782), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1095), .A2(new_n1097), .A3(new_n1098), .A4(new_n1100), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n804), .A2(new_n336), .B1(new_n859), .B2(new_n781), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT112), .Z(new_n1103));
  INV_X1    g0903(.A(G159), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n790), .A2(new_n860), .B1(new_n777), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(new_n1105), .B(KEYINPUT51), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n814), .A2(G77), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n278), .B1(new_n786), .B2(G87), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G50), .A2(new_n796), .B1(new_n793), .B2(new_n1074), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1101), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n821), .ZN(new_n1112));
  INV_X1    g0912(.A(new_n832), .ZN(new_n1113));
  OAI221_X1 g0913(.A(new_n837), .B1(new_n481), .B2(new_n212), .C1(new_n1113), .C2(new_n242), .ZN(new_n1114));
  NAND4_X1  g0914(.A1(new_n1094), .A2(new_n827), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1020), .A2(new_n733), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1018), .B1(new_n1012), .B2(new_n1019), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1115), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1022), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT110), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1019), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1011), .A2(new_n727), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1120), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1012), .A2(KEYINPUT110), .A3(new_n1019), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1119), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1092), .B1(new_n1118), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n1022), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1088), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1129), .A2(new_n733), .A3(new_n1020), .ZN(new_n1130));
  NAND4_X1  g0930(.A1(new_n1128), .A2(new_n1130), .A3(KEYINPUT113), .A4(new_n1115), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1126), .A2(new_n1131), .ZN(G390));
  OR2_X1    g0932(.A1(new_n971), .A2(new_n835), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n847), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n827), .B1(new_n1074), .B2(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n777), .A2(new_n478), .B1(new_n792), .B2(new_n481), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n284), .B(new_n1136), .C1(G68), .C2(new_n786), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n795), .A2(new_n536), .B1(new_n781), .B2(new_n517), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G283), .B2(new_n791), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1137), .A2(new_n813), .A3(new_n1107), .A4(new_n1139), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n787), .A2(new_n217), .B1(new_n863), .B2(new_n777), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n284), .B1(new_n1036), .B2(new_n795), .ZN(new_n1142));
  INV_X1    g0942(.A(G128), .ZN(new_n1143));
  INV_X1    g0943(.A(G125), .ZN(new_n1144));
  OAI22_X1  g0944(.A1(new_n790), .A2(new_n1143), .B1(new_n781), .B2(new_n1144), .ZN(new_n1145));
  NOR3_X1   g0945(.A1(new_n1141), .A2(new_n1142), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n814), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(KEYINPUT54), .B(G143), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(new_n1148), .B(KEYINPUT116), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1146), .B1(new_n1104), .B2(new_n1147), .C1(new_n792), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n805), .A2(G150), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT53), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1140), .B1(new_n1151), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1135), .B1(new_n1154), .B2(new_n821), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1133), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n961), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n871), .B1(new_n745), .B2(new_n874), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1157), .B1(new_n1158), .B2(new_n952), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1159), .B(new_n962), .C1(new_n969), .C2(new_n970), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n967), .A2(new_n961), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n873), .A2(new_n372), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n871), .B1(new_n743), .B2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1161), .B1(new_n952), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n771), .A2(G330), .A3(new_n874), .A4(new_n920), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1160), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT114), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1160), .A2(new_n1167), .A3(new_n1164), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n947), .A2(G330), .A3(new_n920), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1167), .B1(new_n1160), .B2(new_n1164), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1166), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1156), .B1(new_n1173), .B2(new_n1119), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n680), .A2(new_n974), .A3(new_n681), .A4(new_n942), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1158), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n770), .A2(new_n768), .ZN(new_n1178));
  OAI211_X1 g0978(.A(G330), .B(new_n874), .C1(new_n1178), .C2(new_n921), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1179), .A2(new_n952), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1177), .B1(new_n1180), .B2(new_n1170), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n947), .A2(G330), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n952), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n1163), .A3(new_n1165), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1176), .B1(new_n1181), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1186), .A2(KEYINPUT114), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1187), .A2(new_n1168), .A3(new_n1170), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1185), .B1(new_n1188), .B2(new_n1166), .ZN(new_n1189));
  OAI211_X1 g0989(.A(new_n1166), .B(new_n1185), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(KEYINPUT115), .B2(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1181), .A2(new_n1184), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1176), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1173), .A2(KEYINPUT115), .A3(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(new_n733), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1175), .B1(new_n1191), .B2(new_n1196), .ZN(G378));
  NOR2_X1   g0997(.A1(new_n267), .A2(new_n717), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT55), .ZN(new_n1199));
  INV_X1    g0999(.A(new_n1199), .ZN(new_n1200));
  XOR2_X1   g1000(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1201));
  NAND2_X1  g1001(.A1(new_n303), .A2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n303), .A2(new_n1201), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1200), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  OR2_X1    g1005(.A1(new_n303), .A2(new_n1201), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1206), .A2(new_n1199), .A3(new_n1202), .ZN(new_n1207));
  AND2_X1   g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n949), .B2(G330), .ZN(new_n1209));
  AND4_X1   g1009(.A1(G330), .A2(new_n925), .A3(new_n939), .A4(new_n1208), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n972), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n915), .A2(new_n937), .A3(new_n968), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(KEYINPUT101), .A2(new_n1212), .B1(new_n946), .B2(KEYINPUT39), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n963), .B(new_n968), .C1(new_n908), .C2(new_n915), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n961), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n957), .A2(new_n946), .B1(new_n676), .B2(new_n717), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(new_n1208), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n940), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n949), .A2(G330), .A3(new_n1208), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1219), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1211), .A2(new_n1022), .A3(new_n1221), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n827), .B1(G50), .B2(new_n1134), .ZN(new_n1223));
  OAI211_X1 g1023(.A(new_n244), .B(new_n268), .C1(new_n787), .C2(new_n816), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n795), .A2(new_n863), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n790), .A2(new_n1144), .B1(new_n777), .B2(new_n1143), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(G137), .C2(new_n793), .ZN(new_n1227));
  OAI221_X1 g1027(.A(new_n1227), .B1(new_n860), .B2(new_n1147), .C1(new_n804), .C2(new_n1150), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1228), .A2(KEYINPUT59), .ZN(new_n1229));
  AOI211_X1 g1029(.A(new_n1224), .B(new_n1229), .C1(G124), .C2(new_n782), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(KEYINPUT59), .B2(new_n1228), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n284), .A2(G41), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G50), .B(new_n1232), .C1(new_n244), .C2(new_n268), .ZN(new_n1233));
  OAI22_X1  g1033(.A1(new_n787), .A2(new_n392), .B1(new_n478), .B2(new_n790), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n536), .B2(new_n777), .ZN(new_n1235));
  OAI22_X1  g1035(.A1(new_n795), .A2(new_n481), .B1(new_n781), .B2(new_n784), .ZN(new_n1236));
  NOR3_X1   g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n638), .A2(new_n793), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1237), .A2(new_n1044), .A3(new_n1066), .A4(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT58), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1233), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1231), .B(new_n1241), .C1(new_n1240), .C2(new_n1239), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1223), .B1(new_n1242), .B2(new_n821), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n1208), .B2(new_n835), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1222), .A2(KEYINPUT118), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT118), .B1(new_n1222), .B2(new_n1244), .ZN(new_n1246));
  NOR2_X1   g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1190), .A2(new_n1193), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1211), .A2(KEYINPUT57), .A3(new_n1221), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1250), .A2(new_n733), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1211), .A2(new_n1221), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1247), .B1(new_n1251), .B2(new_n1254), .ZN(G375));
  NAND3_X1  g1055(.A1(new_n1181), .A2(new_n1176), .A3(new_n1184), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1257), .A2(new_n1002), .A3(new_n1185), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1192), .A2(new_n1022), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n826), .B1(new_n336), .B2(new_n847), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n804), .A2(new_n481), .B1(new_n850), .B2(new_n781), .ZN(new_n1261));
  XOR2_X1   g1061(.A(new_n1261), .B(KEYINPUT120), .Z(new_n1262));
  OAI22_X1  g1062(.A1(new_n478), .A2(new_n795), .B1(new_n777), .B2(new_n784), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n790), .A2(new_n517), .B1(new_n792), .B2(new_n536), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1038), .A2(KEYINPUT119), .A3(new_n278), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT119), .B1(new_n1038), .B2(new_n278), .ZN(new_n1267));
  OAI211_X1 g1067(.A(new_n1063), .B(new_n1265), .C1(new_n1266), .C2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n814), .A2(G50), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1104), .A2(new_n804), .B1(new_n1150), .B2(new_n795), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n284), .B1(new_n787), .B2(new_n392), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n790), .A2(new_n863), .B1(new_n792), .B2(new_n860), .ZN(new_n1273));
  OAI22_X1  g1073(.A1(new_n1036), .A2(new_n777), .B1(new_n781), .B2(new_n1143), .ZN(new_n1274));
  NOR4_X1   g1074(.A1(new_n1271), .A2(new_n1272), .A3(new_n1273), .A4(new_n1274), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1262), .A2(new_n1269), .B1(new_n1270), .B2(new_n1275), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1260), .B1(new_n822), .B2(new_n1276), .C1(new_n920), .C2(new_n835), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1259), .A2(new_n1277), .ZN(new_n1278));
  OR2_X1    g1078(.A1(new_n1258), .A2(new_n1278), .ZN(G381));
  NAND4_X1  g1079(.A1(new_n1126), .A2(new_n1131), .A3(new_n1023), .A4(new_n1051), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1280), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(G375), .A2(G378), .ZN(new_n1282));
  INV_X1    g1082(.A(G396), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1283), .B(new_n1087), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1284), .A2(G381), .A3(G384), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1281), .A2(new_n1282), .A3(new_n1285), .ZN(G407));
  OR3_X1    g1086(.A1(new_n715), .A2(KEYINPUT121), .A3(G343), .ZN(new_n1287));
  OAI21_X1  g1087(.A(KEYINPUT121), .B1(new_n715), .B2(G343), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  XOR2_X1   g1089(.A(new_n1289), .B(KEYINPUT122), .Z(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1282), .A2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  AOI21_X1  g1093(.A(new_n1252), .B1(new_n1190), .B2(new_n1193), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1250), .B(new_n733), .C1(KEYINPUT57), .C2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(G378), .A2(new_n1295), .A3(new_n1247), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1190), .A2(KEYINPUT115), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1173), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1297), .B1(new_n1298), .B2(new_n1185), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n734), .B1(new_n1189), .B2(KEYINPUT115), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1174), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1301));
  AND2_X1   g1101(.A1(new_n1222), .A2(new_n1244), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1294), .ZN(new_n1303));
  OAI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1002), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1301), .A2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1296), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1290), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1194), .A2(new_n733), .ZN(new_n1308));
  OR2_X1    g1108(.A1(new_n1256), .A2(KEYINPUT60), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1256), .A2(KEYINPUT60), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1309), .B2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(G384), .ZN(new_n1312));
  OR3_X1    g1112(.A1(new_n1311), .A2(new_n1312), .A3(new_n1278), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1312), .B1(new_n1311), .B2(new_n1278), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1313), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT63), .ZN(new_n1317));
  OAI21_X1  g1117(.A(KEYINPUT124), .B1(new_n1307), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1291), .B1(new_n1296), .B2(new_n1305), .ZN(new_n1319));
  INV_X1    g1119(.A(KEYINPUT124), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1319), .A2(new_n1320), .A3(KEYINPUT63), .A4(new_n1316), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1318), .A2(new_n1321), .ZN(new_n1322));
  NAND2_X1  g1122(.A1(G390), .A2(G387), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(G393), .A2(G396), .ZN(new_n1324));
  INV_X1    g1124(.A(KEYINPUT123), .ZN(new_n1325));
  AND3_X1   g1125(.A1(new_n1324), .A2(new_n1325), .A3(new_n1284), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1325), .B1(new_n1324), .B2(new_n1284), .ZN(new_n1327));
  NOR2_X1   g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  AND3_X1   g1128(.A1(new_n1323), .A2(new_n1328), .A3(new_n1280), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1323), .B2(new_n1280), .ZN(new_n1330));
  NOR2_X1   g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1289), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1296), .B2(new_n1305), .ZN(new_n1333));
  AND2_X1   g1133(.A1(new_n1332), .A2(G2897), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1313), .A2(new_n1314), .A3(new_n1334), .ZN(new_n1335));
  AOI22_X1  g1135(.A1(new_n1313), .A2(new_n1314), .B1(G2897), .B2(new_n1291), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(KEYINPUT63), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1306), .A2(new_n1289), .A3(new_n1316), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1338), .A2(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT61), .ZN(new_n1341));
  NAND4_X1  g1141(.A1(new_n1322), .A2(new_n1331), .A3(new_n1340), .A4(new_n1341), .ZN(new_n1342));
  OAI21_X1  g1142(.A(new_n1341), .B1(new_n1319), .B2(new_n1337), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1313), .A2(KEYINPUT62), .A3(new_n1314), .ZN(new_n1344));
  AOI211_X1 g1144(.A(new_n1291), .B(new_n1344), .C1(new_n1296), .C2(new_n1305), .ZN(new_n1345));
  AOI21_X1  g1145(.A(KEYINPUT62), .B1(new_n1333), .B2(new_n1316), .ZN(new_n1346));
  AOI21_X1  g1146(.A(new_n1345), .B1(new_n1346), .B2(KEYINPUT125), .ZN(new_n1347));
  INV_X1    g1147(.A(KEYINPUT62), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1339), .A2(new_n1348), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT125), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1349), .A2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1343), .B1(new_n1347), .B2(new_n1351), .ZN(new_n1352));
  OAI21_X1  g1152(.A(new_n1342), .B1(new_n1352), .B2(new_n1331), .ZN(G405));
  NAND2_X1  g1153(.A1(G375), .A2(new_n1301), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT126), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1354), .A2(new_n1355), .A3(new_n1296), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(G375), .A2(KEYINPUT126), .A3(new_n1301), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1356), .A2(new_n1316), .A3(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT127), .ZN(new_n1359));
  AOI211_X1 g1159(.A(new_n1359), .B(new_n1316), .C1(new_n1356), .C2(new_n1357), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1355), .B1(G375), .B2(new_n1301), .ZN(new_n1361));
  AOI21_X1  g1161(.A(G378), .B1(new_n1295), .B2(new_n1247), .ZN(new_n1362));
  OAI21_X1  g1162(.A(new_n1357), .B1(new_n1361), .B2(new_n1362), .ZN(new_n1363));
  AOI21_X1  g1163(.A(KEYINPUT127), .B1(new_n1363), .B2(new_n1315), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1358), .B1(new_n1360), .B2(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(new_n1331), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  OAI211_X1 g1167(.A(new_n1331), .B(new_n1358), .C1(new_n1360), .C2(new_n1364), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1367), .A2(new_n1368), .ZN(G402));
endmodule


