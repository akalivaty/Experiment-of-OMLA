

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n674, n675, n676, n677, n678, n679, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797;

  NOR2_X1 U375 ( .A1(n658), .A2(n706), .ZN(n685) );
  NAND2_X1 U376 ( .A1(n384), .A2(n381), .ZN(n658) );
  NOR2_X1 U377 ( .A1(n644), .A2(n655), .ZN(n383) );
  XNOR2_X1 U378 ( .A(n353), .B(n674), .ZN(G51) );
  NAND2_X1 U379 ( .A1(n672), .A2(n678), .ZN(n353) );
  XNOR2_X1 U380 ( .A(n354), .B(n681), .ZN(G60) );
  NAND2_X1 U381 ( .A1(n679), .A2(n678), .ZN(n354) );
  XNOR2_X2 U382 ( .A(n362), .B(n482), .ZN(n777) );
  XOR2_X1 U383 ( .A(G104), .B(KEYINPUT12), .Z(n455) );
  NOR2_X1 U384 ( .A1(n682), .A2(n795), .ZN(n609) );
  INV_X2 U385 ( .A(G953), .ZN(n787) );
  AND2_X2 U386 ( .A1(n580), .A2(n579), .ZN(n586) );
  NAND2_X2 U387 ( .A1(n683), .A2(n535), .ZN(n536) );
  OR2_X2 U388 ( .A1(n693), .A2(G902), .ZN(n444) );
  XNOR2_X2 U389 ( .A(n538), .B(n537), .ZN(n742) );
  OR2_X2 U390 ( .A1(n554), .A2(n625), .ZN(n538) );
  NOR2_X1 U391 ( .A1(n742), .A2(n539), .ZN(n540) );
  NOR2_X1 U392 ( .A1(G953), .A2(G237), .ZN(n461) );
  NOR2_X1 U393 ( .A1(n726), .A2(n728), .ZN(n595) );
  NAND2_X1 U394 ( .A1(n528), .A2(n560), .ZN(n726) );
  XNOR2_X1 U395 ( .A(n483), .B(n481), .ZN(n362) );
  INV_X1 U396 ( .A(KEYINPUT92), .ZN(n364) );
  NOR2_X1 U397 ( .A1(n634), .A2(n633), .ZN(n635) );
  AND2_X1 U398 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U399 ( .A(KEYINPUT41), .B(n595), .Z(n741) );
  OR2_X1 U400 ( .A1(n599), .A2(n373), .ZN(n370) );
  NOR2_X1 U401 ( .A1(n503), .A2(n594), .ZN(n505) );
  BUF_X1 U402 ( .A(n503), .Z(n501) );
  XNOR2_X1 U403 ( .A(n500), .B(n499), .ZN(n503) );
  AND2_X1 U404 ( .A1(n410), .A2(n373), .ZN(n372) );
  NOR2_X2 U405 ( .A1(n658), .A2(n706), .ZN(n355) );
  BUF_X1 U406 ( .A(n784), .Z(n356) );
  XNOR2_X1 U407 ( .A(n471), .B(n395), .ZN(n784) );
  XNOR2_X1 U408 ( .A(n490), .B(n394), .ZN(n471) );
  BUF_X1 U409 ( .A(n513), .Z(n357) );
  AND2_X4 U410 ( .A1(n652), .A2(n643), .ZN(n646) );
  NOR2_X2 U411 ( .A1(n644), .A2(n379), .ZN(n378) );
  XNOR2_X2 U412 ( .A(n646), .B(KEYINPUT75), .ZN(n644) );
  XNOR2_X2 U413 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n783) );
  XNOR2_X1 U414 ( .A(n587), .B(KEYINPUT64), .ZN(n588) );
  INV_X1 U415 ( .A(G134), .ZN(n394) );
  INV_X1 U416 ( .A(KEYINPUT91), .ZN(n363) );
  XOR2_X1 U417 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n411) );
  XNOR2_X1 U418 ( .A(G131), .B(G140), .ZN(n459) );
  XOR2_X1 U419 ( .A(n498), .B(KEYINPUT96), .Z(n499) );
  XNOR2_X1 U420 ( .A(n466), .B(n465), .ZN(n528) );
  XNOR2_X1 U421 ( .A(n464), .B(KEYINPUT13), .ZN(n465) );
  INV_X1 U422 ( .A(G475), .ZN(n464) );
  XNOR2_X1 U423 ( .A(n375), .B(n374), .ZN(n482) );
  XNOR2_X1 U424 ( .A(G119), .B(G116), .ZN(n374) );
  XNOR2_X1 U425 ( .A(n397), .B(G113), .ZN(n375) );
  INV_X1 U426 ( .A(KEYINPUT3), .ZN(n397) );
  NOR2_X1 U427 ( .A1(n645), .A2(KEYINPUT66), .ZN(n382) );
  XNOR2_X1 U428 ( .A(G116), .B(G122), .ZN(n470) );
  INV_X1 U429 ( .A(G107), .ZN(n472) );
  XNOR2_X1 U430 ( .A(n784), .B(n396), .ZN(n442) );
  NOR2_X1 U431 ( .A1(n453), .A2(n368), .ZN(n367) );
  NOR2_X1 U432 ( .A1(n410), .A2(n373), .ZN(n368) );
  INV_X1 U433 ( .A(G237), .ZN(n409) );
  NAND2_X1 U434 ( .A1(n496), .A2(n387), .ZN(n386) );
  NAND2_X1 U435 ( .A1(KEYINPUT2), .A2(n388), .ZN(n387) );
  XNOR2_X1 U436 ( .A(KEYINPUT70), .B(G137), .ZN(n395) );
  XNOR2_X1 U437 ( .A(n783), .B(G101), .ZN(n487) );
  XNOR2_X1 U438 ( .A(KEYINPUT17), .B(KEYINPUT93), .ZN(n484) );
  XNOR2_X1 U439 ( .A(KEYINPUT18), .B(KEYINPUT95), .ZN(n489) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n445) );
  INV_X1 U441 ( .A(KEYINPUT0), .ZN(n376) );
  OR2_X1 U442 ( .A1(n662), .A2(G902), .ZN(n407) );
  XNOR2_X1 U443 ( .A(KEYINPUT5), .B(G131), .ZN(n399) );
  XNOR2_X1 U444 ( .A(KEYINPUT101), .B(KEYINPUT102), .ZN(n398) );
  XNOR2_X1 U445 ( .A(G137), .B(G119), .ZN(n418) );
  XNOR2_X1 U446 ( .A(n423), .B(n422), .ZN(n424) );
  INV_X1 U447 ( .A(KEYINPUT97), .ZN(n422) );
  XNOR2_X1 U448 ( .A(G128), .B(G140), .ZN(n423) );
  XNOR2_X1 U449 ( .A(n463), .B(n462), .ZN(n675) );
  XNOR2_X1 U450 ( .A(n785), .B(n392), .ZN(n462) );
  XNOR2_X1 U451 ( .A(G143), .B(G113), .ZN(n457) );
  NOR2_X1 U452 ( .A1(n369), .A2(n366), .ZN(n527) );
  XOR2_X1 U453 ( .A(KEYINPUT16), .B(G122), .Z(n481) );
  NAND2_X1 U454 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U455 ( .A(n475), .B(n474), .ZN(n686) );
  XNOR2_X1 U456 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U457 ( .A(n675), .B(KEYINPUT59), .ZN(n676) );
  INV_X1 U458 ( .A(n369), .ZN(n365) );
  XNOR2_X1 U459 ( .A(n501), .B(n525), .ZN(n593) );
  INV_X1 U460 ( .A(n593), .ZN(n724) );
  AND2_X1 U461 ( .A1(n365), .A2(n367), .ZN(n358) );
  OR2_X1 U462 ( .A1(n496), .A2(KEYINPUT66), .ZN(n359) );
  NAND2_X1 U463 ( .A1(n390), .A2(KEYINPUT66), .ZN(n360) );
  NAND2_X1 U464 ( .A1(n361), .A2(n380), .ZN(n384) );
  NAND2_X1 U465 ( .A1(n389), .A2(n378), .ZN(n361) );
  XNOR2_X1 U466 ( .A(n505), .B(n504), .ZN(n616) );
  XNOR2_X1 U467 ( .A(n566), .B(n363), .ZN(n582) );
  XNOR2_X2 U468 ( .A(n536), .B(n364), .ZN(n566) );
  NOR2_X2 U469 ( .A1(n656), .A2(n657), .ZN(n706) );
  XNOR2_X2 U470 ( .A(n619), .B(KEYINPUT79), .ZN(n760) );
  XNOR2_X1 U471 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U472 ( .A(n427), .B(n426), .ZN(n530) );
  XNOR2_X2 U473 ( .A(n432), .B(n431), .ZN(n553) );
  INV_X2 U474 ( .A(n553), .ZN(n712) );
  BUF_X2 U475 ( .A(n655), .Z(n656) );
  XNOR2_X2 U476 ( .A(n437), .B(n436), .ZN(n483) );
  NAND2_X1 U477 ( .A1(n724), .A2(n367), .ZN(n366) );
  NAND2_X1 U478 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U479 ( .A1(n599), .A2(n372), .ZN(n371) );
  INV_X1 U480 ( .A(KEYINPUT30), .ZN(n373) );
  INV_X1 U481 ( .A(n357), .ZN(n539) );
  XNOR2_X2 U482 ( .A(n377), .B(n376), .ZN(n513) );
  NAND2_X1 U483 ( .A1(n616), .A2(n509), .ZN(n377) );
  INV_X1 U484 ( .A(n655), .ZN(n389) );
  INV_X1 U485 ( .A(n385), .ZN(n379) );
  NAND2_X1 U486 ( .A1(n385), .A2(n360), .ZN(n380) );
  NAND2_X1 U487 ( .A1(n359), .A2(n386), .ZN(n385) );
  INV_X1 U488 ( .A(KEYINPUT66), .ZN(n388) );
  INV_X1 U489 ( .A(KEYINPUT2), .ZN(n390) );
  XOR2_X1 U490 ( .A(KEYINPUT109), .B(n447), .Z(n391) );
  AND2_X1 U491 ( .A1(G214), .A2(n461), .ZN(n392) );
  XOR2_X1 U492 ( .A(n639), .B(KEYINPUT110), .Z(n393) );
  AND2_X1 U493 ( .A1(n566), .A2(n573), .ZN(n572) );
  NAND2_X1 U494 ( .A1(n572), .A2(n571), .ZN(n578) );
  INV_X1 U495 ( .A(n713), .ZN(n510) );
  INV_X1 U496 ( .A(KEYINPUT19), .ZN(n504) );
  BUF_X1 U497 ( .A(n355), .Z(n690) );
  XNOR2_X1 U498 ( .A(n478), .B(n477), .ZN(n560) );
  XNOR2_X1 U499 ( .A(n592), .B(n591), .ZN(n682) );
  XNOR2_X2 U500 ( .A(G143), .B(G128), .ZN(n490) );
  XNOR2_X1 U501 ( .A(n487), .B(G146), .ZN(n396) );
  XNOR2_X1 U502 ( .A(n399), .B(n398), .ZN(n402) );
  NAND2_X1 U503 ( .A1(G210), .A2(n461), .ZN(n400) );
  XNOR2_X1 U504 ( .A(n400), .B(KEYINPUT100), .ZN(n401) );
  XNOR2_X1 U505 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U506 ( .A(n482), .B(n403), .ZN(n404) );
  XNOR2_X1 U507 ( .A(n442), .B(n404), .ZN(n662) );
  INV_X1 U508 ( .A(KEYINPUT103), .ZN(n405) );
  XNOR2_X1 U509 ( .A(n405), .B(G472), .ZN(n406) );
  XNOR2_X2 U510 ( .A(n407), .B(n406), .ZN(n518) );
  INV_X1 U511 ( .A(KEYINPUT107), .ZN(n408) );
  XNOR2_X1 U512 ( .A(n518), .B(n408), .ZN(n599) );
  INV_X1 U513 ( .A(G902), .ZN(n476) );
  NAND2_X1 U514 ( .A1(n476), .A2(n409), .ZN(n497) );
  AND2_X1 U515 ( .A1(n497), .A2(G214), .ZN(n594) );
  INV_X1 U516 ( .A(n594), .ZN(n410) );
  XNOR2_X2 U517 ( .A(G146), .B(G125), .ZN(n485) );
  XNOR2_X1 U518 ( .A(n411), .B(n485), .ZN(n460) );
  XNOR2_X1 U519 ( .A(n460), .B(KEYINPUT23), .ZN(n412) );
  NAND2_X1 U520 ( .A1(n412), .A2(KEYINPUT72), .ZN(n416) );
  INV_X1 U521 ( .A(n412), .ZN(n414) );
  INV_X1 U522 ( .A(KEYINPUT72), .ZN(n413) );
  NAND2_X1 U523 ( .A1(n414), .A2(n413), .ZN(n415) );
  NAND2_X1 U524 ( .A1(n416), .A2(n415), .ZN(n427) );
  NAND2_X1 U525 ( .A1(G234), .A2(n787), .ZN(n417) );
  XOR2_X1 U526 ( .A(KEYINPUT8), .B(n417), .Z(n467) );
  NAND2_X1 U527 ( .A1(n467), .A2(G221), .ZN(n421) );
  XOR2_X1 U528 ( .A(KEYINPUT24), .B(G110), .Z(n419) );
  XNOR2_X1 U529 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U530 ( .A(n421), .B(n420), .ZN(n425) );
  NAND2_X1 U531 ( .A1(n530), .A2(n476), .ZN(n432) );
  XOR2_X1 U532 ( .A(KEYINPUT98), .B(KEYINPUT25), .Z(n430) );
  XNOR2_X1 U533 ( .A(G902), .B(KEYINPUT15), .ZN(n645) );
  NAND2_X1 U534 ( .A1(G234), .A2(n645), .ZN(n428) );
  XNOR2_X1 U535 ( .A(KEYINPUT20), .B(n428), .ZN(n433) );
  NAND2_X1 U536 ( .A1(n433), .A2(G217), .ZN(n429) );
  XNOR2_X1 U537 ( .A(n430), .B(n429), .ZN(n431) );
  AND2_X1 U538 ( .A1(n433), .A2(G221), .ZN(n435) );
  XNOR2_X1 U539 ( .A(KEYINPUT99), .B(KEYINPUT21), .ZN(n434) );
  XNOR2_X1 U540 ( .A(n435), .B(n434), .ZN(n713) );
  AND2_X2 U541 ( .A1(n553), .A2(n510), .ZN(n709) );
  XNOR2_X2 U542 ( .A(G107), .B(G104), .ZN(n437) );
  XNOR2_X2 U543 ( .A(G110), .B(KEYINPUT74), .ZN(n436) );
  INV_X1 U544 ( .A(n459), .ZN(n439) );
  NAND2_X1 U545 ( .A1(G227), .A2(n787), .ZN(n438) );
  XNOR2_X1 U546 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U547 ( .A(n483), .B(n440), .ZN(n441) );
  XNOR2_X1 U548 ( .A(n442), .B(n441), .ZN(n693) );
  INV_X1 U549 ( .A(G469), .ZN(n443) );
  XNOR2_X2 U550 ( .A(n444), .B(n443), .ZN(n602) );
  XNOR2_X1 U551 ( .A(n445), .B(KEYINPUT14), .ZN(n448) );
  NAND2_X1 U552 ( .A1(G902), .A2(n448), .ZN(n506) );
  NOR2_X1 U553 ( .A1(G900), .A2(n506), .ZN(n446) );
  NAND2_X1 U554 ( .A1(G953), .A2(n446), .ZN(n447) );
  NAND2_X1 U555 ( .A1(G952), .A2(n448), .ZN(n738) );
  INV_X1 U556 ( .A(n738), .ZN(n449) );
  NAND2_X1 U557 ( .A1(n449), .A2(n787), .ZN(n508) );
  NAND2_X1 U558 ( .A1(n391), .A2(n508), .ZN(n450) );
  XNOR2_X1 U559 ( .A(n450), .B(KEYINPUT80), .ZN(n596) );
  INV_X1 U560 ( .A(n596), .ZN(n451) );
  NOR2_X1 U561 ( .A1(n602), .A2(n451), .ZN(n452) );
  NAND2_X1 U562 ( .A1(n709), .A2(n452), .ZN(n453) );
  XNOR2_X1 U563 ( .A(KEYINPUT11), .B(KEYINPUT104), .ZN(n454) );
  XNOR2_X1 U564 ( .A(n455), .B(n454), .ZN(n456) );
  XOR2_X1 U565 ( .A(n456), .B(G122), .Z(n458) );
  XNOR2_X1 U566 ( .A(n458), .B(n457), .ZN(n463) );
  XNOR2_X1 U567 ( .A(n460), .B(n459), .ZN(n785) );
  NOR2_X1 U568 ( .A1(G902), .A2(n675), .ZN(n466) );
  INV_X1 U569 ( .A(n528), .ZN(n480) );
  XOR2_X1 U570 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n469) );
  NAND2_X1 U571 ( .A1(G217), .A2(n467), .ZN(n468) );
  XNOR2_X1 U572 ( .A(n469), .B(n468), .ZN(n475) );
  XNOR2_X1 U573 ( .A(n471), .B(n470), .ZN(n473) );
  NAND2_X1 U574 ( .A1(n686), .A2(n476), .ZN(n478) );
  INV_X1 U575 ( .A(G478), .ZN(n477) );
  INV_X1 U576 ( .A(n560), .ZN(n479) );
  NAND2_X1 U577 ( .A1(n480), .A2(n479), .ZN(n541) );
  XNOR2_X1 U578 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U579 ( .A(n487), .B(n486), .ZN(n494) );
  NAND2_X1 U580 ( .A1(n787), .A2(G224), .ZN(n488) );
  XNOR2_X1 U581 ( .A(n489), .B(n488), .ZN(n492) );
  INV_X1 U582 ( .A(n490), .ZN(n491) );
  XNOR2_X1 U583 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U584 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U585 ( .A(n495), .B(n777), .ZN(n667) );
  INV_X1 U586 ( .A(n645), .ZN(n496) );
  NOR2_X1 U587 ( .A1(n667), .A2(n496), .ZN(n500) );
  NAND2_X1 U588 ( .A1(n497), .A2(G210), .ZN(n498) );
  NOR2_X1 U589 ( .A1(n541), .A2(n501), .ZN(n502) );
  NAND2_X1 U590 ( .A1(n358), .A2(n502), .ZN(n613) );
  XNOR2_X1 U591 ( .A(n613), .B(G143), .ZN(G45) );
  OR2_X1 U592 ( .A1(n787), .A2(G898), .ZN(n779) );
  OR2_X1 U593 ( .A1(n506), .A2(n779), .ZN(n507) );
  NAND2_X1 U594 ( .A1(n508), .A2(n507), .ZN(n509) );
  INV_X1 U595 ( .A(n726), .ZN(n511) );
  AND2_X1 U596 ( .A1(n511), .A2(n510), .ZN(n512) );
  NAND2_X1 U597 ( .A1(n513), .A2(n512), .ZN(n516) );
  INV_X1 U598 ( .A(KEYINPUT68), .ZN(n514) );
  XNOR2_X1 U599 ( .A(n514), .B(KEYINPUT22), .ZN(n515) );
  XNOR2_X1 U600 ( .A(n516), .B(n515), .ZN(n531) );
  BUF_X1 U601 ( .A(n531), .Z(n522) );
  INV_X1 U602 ( .A(KEYINPUT1), .ZN(n517) );
  XNOR2_X2 U603 ( .A(n602), .B(n517), .ZN(n708) );
  XNOR2_X1 U604 ( .A(n708), .B(KEYINPUT94), .ZN(n630) );
  XNOR2_X1 U605 ( .A(n518), .B(KEYINPUT6), .ZN(n625) );
  XNOR2_X1 U606 ( .A(n625), .B(KEYINPUT78), .ZN(n519) );
  AND2_X1 U607 ( .A1(n519), .A2(n712), .ZN(n520) );
  AND2_X1 U608 ( .A1(n630), .A2(n520), .ZN(n521) );
  NAND2_X1 U609 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U610 ( .A(n523), .B(KEYINPUT32), .ZN(n535) );
  XOR2_X1 U611 ( .A(G119), .B(KEYINPUT127), .Z(n524) );
  XNOR2_X1 U612 ( .A(n535), .B(n524), .ZN(G21) );
  INV_X1 U613 ( .A(KEYINPUT38), .ZN(n525) );
  INV_X1 U614 ( .A(KEYINPUT39), .ZN(n526) );
  XNOR2_X1 U615 ( .A(n527), .B(n526), .ZN(n590) );
  INV_X1 U616 ( .A(n590), .ZN(n529) );
  XNOR2_X1 U617 ( .A(n528), .B(KEYINPUT105), .ZN(n561) );
  NOR2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n764) );
  INV_X1 U619 ( .A(n764), .ZN(n610) );
  OR2_X1 U620 ( .A1(n529), .A2(n610), .ZN(n648) );
  XNOR2_X1 U621 ( .A(n648), .B(G134), .ZN(G36) );
  INV_X1 U622 ( .A(n708), .ZN(n640) );
  AND2_X2 U623 ( .A1(n531), .A2(n640), .ZN(n549) );
  INV_X1 U624 ( .A(n599), .ZN(n532) );
  NAND2_X1 U625 ( .A1(n549), .A2(n532), .ZN(n533) );
  XNOR2_X1 U626 ( .A(n533), .B(KEYINPUT67), .ZN(n534) );
  NAND2_X1 U627 ( .A1(n534), .A2(n712), .ZN(n683) );
  NAND2_X1 U628 ( .A1(n709), .A2(n708), .ZN(n554) );
  XOR2_X1 U629 ( .A(KEYINPUT108), .B(KEYINPUT33), .Z(n537) );
  XNOR2_X1 U630 ( .A(n540), .B(KEYINPUT34), .ZN(n543) );
  XNOR2_X1 U631 ( .A(n541), .B(KEYINPUT77), .ZN(n542) );
  NAND2_X1 U632 ( .A1(n543), .A2(n542), .ZN(n547) );
  XNOR2_X1 U633 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n545) );
  INV_X1 U634 ( .A(KEYINPUT76), .ZN(n544) );
  XNOR2_X1 U635 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X2 U636 ( .A(n547), .B(n546), .ZN(n796) );
  NAND2_X1 U637 ( .A1(n582), .A2(n796), .ZN(n548) );
  NAND2_X1 U638 ( .A1(n548), .A2(KEYINPUT73), .ZN(n580) );
  BUF_X1 U639 ( .A(n549), .Z(n550) );
  NAND2_X1 U640 ( .A1(n550), .A2(n625), .ZN(n551) );
  XNOR2_X1 U641 ( .A(n551), .B(KEYINPUT89), .ZN(n552) );
  AND2_X1 U642 ( .A1(n553), .A2(n552), .ZN(n751) );
  INV_X1 U643 ( .A(n518), .ZN(n557) );
  OR2_X1 U644 ( .A1(n554), .A2(n557), .ZN(n719) );
  NOR2_X1 U645 ( .A1(n719), .A2(n539), .ZN(n556) );
  INV_X1 U646 ( .A(KEYINPUT31), .ZN(n555) );
  XNOR2_X1 U647 ( .A(n556), .B(n555), .ZN(n765) );
  NAND2_X1 U648 ( .A1(n709), .A2(n557), .ZN(n558) );
  OR2_X1 U649 ( .A1(n539), .A2(n558), .ZN(n559) );
  NOR2_X1 U650 ( .A1(n602), .A2(n559), .ZN(n754) );
  OR2_X1 U651 ( .A1(n765), .A2(n754), .ZN(n564) );
  NAND2_X1 U652 ( .A1(n561), .A2(n560), .ZN(n563) );
  INV_X1 U653 ( .A(KEYINPUT106), .ZN(n562) );
  XNOR2_X1 U654 ( .A(n563), .B(n562), .ZN(n627) );
  BUF_X1 U655 ( .A(n627), .Z(n762) );
  OR2_X1 U656 ( .A1(n762), .A2(n764), .ZN(n727) );
  AND2_X1 U657 ( .A1(n564), .A2(n727), .ZN(n565) );
  NOR2_X2 U658 ( .A1(n751), .A2(n565), .ZN(n573) );
  INV_X1 U659 ( .A(n796), .ZN(n567) );
  NAND2_X1 U660 ( .A1(n567), .A2(KEYINPUT90), .ZN(n570) );
  INV_X1 U661 ( .A(KEYINPUT73), .ZN(n568) );
  AND2_X1 U662 ( .A1(n568), .A2(KEYINPUT44), .ZN(n569) );
  INV_X1 U663 ( .A(n573), .ZN(n576) );
  INV_X1 U664 ( .A(KEYINPUT44), .ZN(n574) );
  NAND2_X1 U665 ( .A1(n574), .A2(KEYINPUT90), .ZN(n575) );
  OR2_X1 U666 ( .A1(n576), .A2(n575), .ZN(n577) );
  NAND2_X1 U667 ( .A1(n578), .A2(n577), .ZN(n579) );
  NOR2_X1 U668 ( .A1(KEYINPUT44), .A2(KEYINPUT73), .ZN(n581) );
  NAND2_X1 U669 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U670 ( .A1(n583), .A2(KEYINPUT90), .ZN(n584) );
  NAND2_X1 U671 ( .A1(n584), .A2(n796), .ZN(n585) );
  NAND2_X1 U672 ( .A1(n586), .A2(n585), .ZN(n589) );
  XNOR2_X1 U673 ( .A(KEYINPUT85), .B(KEYINPUT45), .ZN(n587) );
  XNOR2_X2 U674 ( .A(n589), .B(n588), .ZN(n655) );
  NAND2_X1 U675 ( .A1(n590), .A2(n627), .ZN(n592) );
  XNOR2_X1 U676 ( .A(KEYINPUT111), .B(KEYINPUT40), .ZN(n591) );
  NAND2_X1 U677 ( .A1(n724), .A2(n410), .ZN(n728) );
  AND2_X1 U678 ( .A1(n510), .A2(n596), .ZN(n597) );
  NAND2_X1 U679 ( .A1(n597), .A2(n712), .ZN(n598) );
  XNOR2_X1 U680 ( .A(n598), .B(KEYINPUT71), .ZN(n624) );
  NAND2_X1 U681 ( .A1(n624), .A2(n599), .ZN(n601) );
  INV_X1 U682 ( .A(KEYINPUT28), .ZN(n600) );
  XNOR2_X1 U683 ( .A(n601), .B(n600), .ZN(n604) );
  INV_X1 U684 ( .A(n602), .ZN(n603) );
  AND2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n618) );
  NAND2_X1 U686 ( .A1(n741), .A2(n618), .ZN(n607) );
  INV_X1 U687 ( .A(KEYINPUT112), .ZN(n605) );
  XNOR2_X1 U688 ( .A(n605), .B(KEYINPUT42), .ZN(n606) );
  XNOR2_X1 U689 ( .A(n607), .B(n606), .ZN(n795) );
  XNOR2_X1 U690 ( .A(KEYINPUT88), .B(KEYINPUT46), .ZN(n608) );
  XNOR2_X1 U691 ( .A(n609), .B(n608), .ZN(n636) );
  NAND2_X1 U692 ( .A1(KEYINPUT47), .A2(n610), .ZN(n611) );
  OR2_X1 U693 ( .A1(n627), .A2(n611), .ZN(n612) );
  XOR2_X1 U694 ( .A(KEYINPUT83), .B(n612), .Z(n614) );
  NAND2_X1 U695 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U696 ( .A(n615), .B(KEYINPUT82), .ZN(n634) );
  BUF_X1 U697 ( .A(n616), .Z(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n619) );
  INV_X1 U699 ( .A(KEYINPUT47), .ZN(n620) );
  NAND2_X1 U700 ( .A1(n727), .A2(n620), .ZN(n621) );
  NAND2_X1 U701 ( .A1(n760), .A2(n621), .ZN(n623) );
  OR2_X2 U702 ( .A1(n760), .A2(KEYINPUT47), .ZN(n622) );
  NAND2_X1 U703 ( .A1(n623), .A2(n622), .ZN(n632) );
  NAND2_X1 U704 ( .A1(n624), .A2(n410), .ZN(n626) );
  NOR2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n628), .A2(n627), .ZN(n639) );
  NOR2_X1 U707 ( .A1(n639), .A2(n501), .ZN(n629) );
  XNOR2_X1 U708 ( .A(n629), .B(KEYINPUT36), .ZN(n631) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n767) );
  NAND2_X1 U710 ( .A1(n632), .A2(n767), .ZN(n633) );
  NAND2_X1 U711 ( .A1(n635), .A2(n636), .ZN(n638) );
  XNOR2_X1 U712 ( .A(KEYINPUT87), .B(KEYINPUT48), .ZN(n637) );
  XNOR2_X2 U713 ( .A(n638), .B(n637), .ZN(n652) );
  NAND2_X1 U714 ( .A1(n393), .A2(n640), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n641), .B(KEYINPUT43), .ZN(n642) );
  NAND2_X1 U716 ( .A1(n642), .A2(n501), .ZN(n770) );
  AND2_X1 U717 ( .A1(n770), .A2(n648), .ZN(n643) );
  NOR2_X1 U718 ( .A1(n390), .A2(KEYINPUT81), .ZN(n647) );
  NAND2_X1 U719 ( .A1(n646), .A2(n647), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n770), .A2(KEYINPUT81), .ZN(n650) );
  AND2_X1 U721 ( .A1(n648), .A2(KEYINPUT2), .ZN(n649) );
  NOR2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U723 ( .A1(n652), .A2(n651), .ZN(n653) );
  AND2_X1 U724 ( .A1(n654), .A2(n653), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n355), .A2(G217), .ZN(n659) );
  XOR2_X1 U726 ( .A(n530), .B(n659), .Z(n661) );
  INV_X1 U727 ( .A(G952), .ZN(n660) );
  NAND2_X1 U728 ( .A1(n660), .A2(G953), .ZN(n678) );
  INV_X1 U729 ( .A(n678), .ZN(n696) );
  NOR2_X1 U730 ( .A1(n661), .A2(n696), .ZN(G66) );
  NAND2_X1 U731 ( .A1(n355), .A2(G472), .ZN(n664) );
  XOR2_X1 U732 ( .A(KEYINPUT62), .B(n662), .Z(n663) );
  XNOR2_X1 U733 ( .A(n664), .B(n663), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n665), .A2(n678), .ZN(n666) );
  XNOR2_X1 U735 ( .A(n666), .B(KEYINPUT63), .ZN(G57) );
  INV_X1 U736 ( .A(KEYINPUT56), .ZN(n674) );
  NAND2_X1 U737 ( .A1(n685), .A2(G210), .ZN(n671) );
  BUF_X1 U738 ( .A(n667), .Z(n669) );
  XNOR2_X1 U739 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n669), .B(n668), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(n672) );
  INV_X1 U742 ( .A(KEYINPUT60), .ZN(n681) );
  NAND2_X1 U743 ( .A1(n685), .A2(G475), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n677), .B(n676), .ZN(n679) );
  XOR2_X1 U745 ( .A(n682), .B(G131), .Z(G33) );
  BUF_X1 U746 ( .A(n683), .Z(n684) );
  XNOR2_X1 U747 ( .A(n684), .B(G110), .ZN(G12) );
  NAND2_X1 U748 ( .A1(n690), .A2(G478), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n686), .B(KEYINPUT123), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n688), .B(n687), .ZN(n689) );
  NOR2_X1 U751 ( .A1(n689), .A2(n696), .ZN(G63) );
  NAND2_X1 U752 ( .A1(n690), .A2(G469), .ZN(n695) );
  XOR2_X1 U753 ( .A(KEYINPUT122), .B(KEYINPUT57), .Z(n691) );
  XNOR2_X1 U754 ( .A(n691), .B(KEYINPUT58), .ZN(n692) );
  XNOR2_X1 U755 ( .A(n693), .B(n692), .ZN(n694) );
  XNOR2_X1 U756 ( .A(n695), .B(n694), .ZN(n697) );
  NOR2_X1 U757 ( .A1(n697), .A2(n696), .ZN(G54) );
  INV_X1 U758 ( .A(n646), .ZN(n698) );
  NOR2_X1 U759 ( .A1(n698), .A2(n656), .ZN(n699) );
  NOR2_X1 U760 ( .A1(n699), .A2(KEYINPUT2), .ZN(n701) );
  INV_X1 U761 ( .A(KEYINPUT84), .ZN(n700) );
  NOR2_X1 U762 ( .A1(n701), .A2(n700), .ZN(n705) );
  NOR2_X1 U763 ( .A1(KEYINPUT2), .A2(KEYINPUT84), .ZN(n702) );
  NAND2_X1 U764 ( .A1(n646), .A2(n702), .ZN(n703) );
  INV_X1 U765 ( .A(n656), .ZN(n772) );
  NOR2_X1 U766 ( .A1(n703), .A2(n772), .ZN(n704) );
  NOR2_X1 U767 ( .A1(n705), .A2(n704), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n748) );
  NOR2_X1 U769 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U770 ( .A(KEYINPUT50), .B(KEYINPUT115), .ZN(n710) );
  XNOR2_X1 U771 ( .A(n711), .B(n710), .ZN(n716) );
  NAND2_X1 U772 ( .A1(n713), .A2(n712), .ZN(n714) );
  XOR2_X1 U773 ( .A(KEYINPUT49), .B(n714), .Z(n715) );
  NAND2_X1 U774 ( .A1(n716), .A2(n715), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n717), .A2(n518), .ZN(n718) );
  XOR2_X1 U776 ( .A(KEYINPUT116), .B(n718), .Z(n720) );
  AND2_X1 U777 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U778 ( .A(n721), .B(KEYINPUT117), .Z(n722) );
  XNOR2_X1 U779 ( .A(KEYINPUT51), .B(n722), .ZN(n723) );
  NAND2_X1 U780 ( .A1(n723), .A2(n741), .ZN(n735) );
  NOR2_X1 U781 ( .A1(n724), .A2(n410), .ZN(n725) );
  NOR2_X1 U782 ( .A1(n726), .A2(n725), .ZN(n731) );
  INV_X1 U783 ( .A(n727), .ZN(n729) );
  NOR2_X1 U784 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U785 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U786 ( .A1(n742), .A2(n732), .ZN(n733) );
  XOR2_X1 U787 ( .A(KEYINPUT118), .B(n733), .Z(n734) );
  NAND2_X1 U788 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U789 ( .A(n736), .B(KEYINPUT119), .ZN(n737) );
  XNOR2_X1 U790 ( .A(n737), .B(KEYINPUT52), .ZN(n739) );
  NOR2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XOR2_X1 U792 ( .A(KEYINPUT120), .B(n740), .Z(n746) );
  INV_X1 U793 ( .A(n741), .ZN(n743) );
  NOR2_X1 U794 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U795 ( .A1(n744), .A2(G953), .ZN(n745) );
  NAND2_X1 U796 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U797 ( .A1(n748), .A2(n747), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n749) );
  XNOR2_X1 U799 ( .A(n750), .B(n749), .ZN(G75) );
  XOR2_X1 U800 ( .A(G101), .B(n751), .Z(G3) );
  XOR2_X1 U801 ( .A(G104), .B(KEYINPUT113), .Z(n753) );
  NAND2_X1 U802 ( .A1(n754), .A2(n762), .ZN(n752) );
  XNOR2_X1 U803 ( .A(n753), .B(n752), .ZN(G6) );
  XOR2_X1 U804 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n756) );
  NAND2_X1 U805 ( .A1(n754), .A2(n764), .ZN(n755) );
  XNOR2_X1 U806 ( .A(n756), .B(n755), .ZN(n757) );
  XNOR2_X1 U807 ( .A(G107), .B(n757), .ZN(G9) );
  XOR2_X1 U808 ( .A(G128), .B(KEYINPUT29), .Z(n759) );
  NAND2_X1 U809 ( .A1(n764), .A2(n760), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n759), .B(n758), .ZN(G30) );
  NAND2_X1 U811 ( .A1(n762), .A2(n760), .ZN(n761) );
  XNOR2_X1 U812 ( .A(n761), .B(G146), .ZN(G48) );
  NAND2_X1 U813 ( .A1(n762), .A2(n765), .ZN(n763) );
  XNOR2_X1 U814 ( .A(n763), .B(G113), .ZN(G15) );
  NAND2_X1 U815 ( .A1(n765), .A2(n764), .ZN(n766) );
  XNOR2_X1 U816 ( .A(n766), .B(G116), .ZN(G18) );
  INV_X1 U817 ( .A(n767), .ZN(n768) );
  XNOR2_X1 U818 ( .A(G125), .B(n768), .ZN(n769) );
  XNOR2_X1 U819 ( .A(n769), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U820 ( .A(n770), .B(G140), .ZN(n771) );
  XNOR2_X1 U821 ( .A(KEYINPUT114), .B(n771), .ZN(G42) );
  NAND2_X1 U822 ( .A1(n772), .A2(n787), .ZN(n776) );
  NAND2_X1 U823 ( .A1(G953), .A2(G224), .ZN(n773) );
  XNOR2_X1 U824 ( .A(KEYINPUT61), .B(n773), .ZN(n774) );
  NAND2_X1 U825 ( .A1(n774), .A2(G898), .ZN(n775) );
  NAND2_X1 U826 ( .A1(n776), .A2(n775), .ZN(n782) );
  XOR2_X1 U827 ( .A(G101), .B(KEYINPUT124), .Z(n778) );
  XNOR2_X1 U828 ( .A(n777), .B(n778), .ZN(n780) );
  NAND2_X1 U829 ( .A1(n780), .A2(n779), .ZN(n781) );
  XOR2_X1 U830 ( .A(n782), .B(n781), .Z(G69) );
  XNOR2_X1 U831 ( .A(n783), .B(n356), .ZN(n786) );
  XNOR2_X1 U832 ( .A(n786), .B(n785), .ZN(n789) );
  XNOR2_X1 U833 ( .A(n646), .B(n789), .ZN(n788) );
  NAND2_X1 U834 ( .A1(n788), .A2(n787), .ZN(n794) );
  XOR2_X1 U835 ( .A(G227), .B(n789), .Z(n790) );
  NAND2_X1 U836 ( .A1(n790), .A2(G900), .ZN(n791) );
  XOR2_X1 U837 ( .A(KEYINPUT125), .B(n791), .Z(n792) );
  NAND2_X1 U838 ( .A1(G953), .A2(n792), .ZN(n793) );
  NAND2_X1 U839 ( .A1(n794), .A2(n793), .ZN(G72) );
  XOR2_X1 U840 ( .A(G137), .B(n795), .Z(G39) );
  XNOR2_X1 U841 ( .A(G122), .B(KEYINPUT126), .ZN(n797) );
  XNOR2_X1 U842 ( .A(n797), .B(n796), .ZN(G24) );
endmodule

