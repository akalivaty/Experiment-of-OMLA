//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 1 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:55 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1218, new_n1219,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G68), .A3(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT64), .Z(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XOR2_X1   g0014(.A(new_n214), .B(KEYINPUT0), .Z(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(new_n210), .ZN(new_n217));
  INV_X1    g0017(.A(G68), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n202), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n219), .A2(G50), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n215), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  INV_X1    g0025(.A(G257), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n223), .B1(new_n224), .B2(new_n225), .C1(new_n205), .C2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n230));
  NAND3_X1  g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n227), .A2(KEYINPUT65), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n212), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n234));
  OR2_X1    g0034(.A1(new_n233), .A2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g0035(.A1(new_n222), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n236), .B(KEYINPUT66), .Z(G361));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(KEYINPUT2), .B(G226), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(G264), .B(G270), .Z(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n242), .B(new_n245), .ZN(G358));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XNOR2_X1  g0050(.A(G107), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n249), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n210), .A3(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n216), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n209), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G50), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n255), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(G50), .B2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n257), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT8), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n268), .A2(G20), .ZN(new_n269));
  NOR2_X1   g0069(.A1(G20), .A2(G33), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n267), .A2(new_n269), .B1(G150), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g0071(.A(G20), .B1(new_n203), .B2(G68), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n263), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n262), .B1(KEYINPUT69), .B2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(KEYINPUT69), .B2(new_n273), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT9), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT72), .ZN(new_n278));
  XNOR2_X1  g0078(.A(new_n277), .B(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT68), .ZN(new_n280));
  AND2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n280), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT3), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(new_n268), .ZN(new_n285));
  NAND2_X1  g0085(.A1(KEYINPUT3), .A2(G33), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n285), .A2(KEYINPUT68), .A3(new_n286), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n288), .A2(G222), .A3(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G77), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n288), .A2(G1698), .ZN(new_n292));
  INV_X1    g0092(.A(G223), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n290), .B1(new_n291), .B2(new_n288), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(G33), .A2(G41), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G1), .A3(G13), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n300), .A2(new_n296), .A3(G274), .ZN(new_n301));
  XNOR2_X1  g0101(.A(KEYINPUT67), .B(G226), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n296), .A3(new_n299), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n298), .A2(new_n301), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(G200), .ZN(new_n305));
  OR2_X1    g0105(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n306));
  INV_X1    g0106(.A(new_n304), .ZN(new_n307));
  AOI22_X1  g0107(.A1(new_n307), .A2(G190), .B1(new_n276), .B2(new_n275), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(KEYINPUT73), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n279), .A2(new_n306), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT10), .ZN(new_n311));
  OAI21_X1  g0111(.A(new_n275), .B1(new_n307), .B2(G169), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n304), .A2(G179), .ZN(new_n313));
  NOR2_X1   g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n311), .A2(new_n315), .ZN(new_n316));
  NAND4_X1  g0116(.A1(new_n283), .A2(new_n287), .A3(G232), .A4(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n283), .A2(new_n287), .A3(G226), .A4(new_n289), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n317), .B(new_n318), .C1(new_n268), .C2(new_n205), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n297), .ZN(new_n320));
  INV_X1    g0120(.A(G238), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n296), .A2(new_n299), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n301), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n320), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n323), .B1(new_n319), .B2(new_n297), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT13), .ZN(new_n328));
  AOI21_X1  g0128(.A(KEYINPUT74), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(KEYINPUT74), .A3(KEYINPUT13), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(G169), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT14), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT14), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n330), .A2(new_n334), .A3(G169), .A4(new_n331), .ZN(new_n335));
  INV_X1    g0135(.A(G179), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n336), .B1(new_n327), .B2(new_n328), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n326), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n255), .A2(new_n218), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT12), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n341), .A2(KEYINPUT76), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT76), .B1(new_n341), .B2(new_n342), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n201), .A2(G20), .A3(G33), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT75), .ZN(new_n346));
  INV_X1    g0146(.A(new_n269), .ZN(new_n347));
  OAI22_X1  g0147(.A1(new_n347), .A2(new_n291), .B1(new_n210), .B2(G68), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n257), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  AND2_X1   g0149(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n349), .A2(KEYINPUT11), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n343), .A2(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n330), .A2(G200), .A3(new_n331), .ZN(new_n354));
  INV_X1    g0154(.A(G190), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n327), .B2(new_n328), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n352), .B1(new_n326), .B2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n258), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n267), .A2(new_n259), .ZN(new_n362));
  OAI22_X1  g0162(.A1(new_n361), .A2(new_n362), .B1(new_n261), .B2(new_n267), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n270), .A2(G159), .ZN(new_n364));
  NAND2_X1  g0164(.A1(G58), .A2(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n210), .B1(new_n219), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n364), .B1(new_n366), .B2(KEYINPUT77), .ZN(new_n367));
  AND2_X1   g0167(.A1(G58), .A2(G68), .ZN(new_n368));
  NOR2_X1   g0168(.A1(G58), .A2(G68), .ZN(new_n369));
  OAI211_X1 g0169(.A(KEYINPUT77), .B(G20), .C1(new_n368), .C2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  OAI21_X1  g0171(.A(KEYINPUT78), .B1(new_n367), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n368), .B2(new_n369), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT77), .ZN(new_n374));
  AOI22_X1  g0174(.A1(new_n373), .A2(new_n374), .B1(G159), .B2(new_n270), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT78), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n376), .A3(new_n370), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n281), .A2(new_n282), .ZN(new_n378));
  AOI21_X1  g0178(.A(KEYINPUT7), .B1(new_n378), .B2(new_n210), .ZN(new_n379));
  AND4_X1   g0179(.A1(KEYINPUT7), .A2(new_n285), .A3(new_n210), .A4(new_n286), .ZN(new_n380));
  OAI21_X1  g0180(.A(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n372), .A2(KEYINPUT16), .A3(new_n377), .A4(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n257), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT16), .ZN(new_n384));
  INV_X1    g0184(.A(new_n380), .ZN(new_n385));
  AOI21_X1  g0185(.A(G20), .B1(new_n283), .B2(new_n287), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n385), .B1(new_n386), .B2(KEYINPUT7), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n387), .A2(G68), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n372), .A2(new_n377), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n383), .B1(new_n390), .B2(KEYINPUT79), .ZN(new_n391));
  AND2_X1   g0191(.A1(new_n372), .A2(new_n377), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n387), .A2(G68), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT16), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT79), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n363), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g0197(.A(KEYINPUT3), .B(G33), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n293), .A2(new_n289), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(G226), .C2(new_n289), .ZN(new_n400));
  NAND2_X1  g0200(.A1(G33), .A2(G87), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n296), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n301), .B1(new_n239), .B2(new_n322), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n402), .B1(KEYINPUT80), .B2(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(G169), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(G179), .B2(new_n406), .ZN(new_n409));
  OAI21_X1  g0209(.A(KEYINPUT18), .B1(new_n397), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n363), .ZN(new_n411));
  INV_X1    g0211(.A(new_n383), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n394), .B2(new_n395), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n390), .A2(KEYINPUT79), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT18), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n406), .A2(G179), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(new_n407), .B2(new_n406), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n415), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n410), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n404), .A2(new_n355), .A3(new_n405), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n422), .B1(new_n406), .B2(G200), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n411), .B(new_n423), .C1(new_n413), .C2(new_n414), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT17), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n397), .A2(KEYINPUT17), .A3(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n421), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n267), .B1(KEYINPUT70), .B2(new_n270), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(KEYINPUT70), .B2(new_n270), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT15), .B(G87), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n433), .A2(new_n347), .B1(new_n210), .B2(new_n291), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n257), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n435), .B(KEYINPUT71), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(G77), .B2(new_n261), .ZN(new_n438));
  INV_X1    g0238(.A(G244), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n301), .B1(new_n439), .B2(new_n322), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n288), .A2(G232), .A3(new_n289), .ZN(new_n441));
  OAI221_X1 g0241(.A(new_n441), .B1(new_n206), .B2(new_n288), .C1(new_n292), .C2(new_n321), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n440), .B1(new_n442), .B2(new_n297), .ZN(new_n443));
  OAI22_X1  g0243(.A1(new_n436), .A2(new_n438), .B1(new_n443), .B2(G169), .ZN(new_n444));
  AND2_X1   g0244(.A1(new_n443), .A2(new_n336), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n436), .A2(new_n438), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n443), .A2(G190), .ZN(new_n449));
  INV_X1    g0249(.A(G200), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n448), .B(new_n449), .C1(new_n450), .C2(new_n443), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  NOR4_X1   g0252(.A1(new_n316), .A2(new_n360), .A3(new_n430), .A4(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT82), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n261), .B2(G97), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n255), .A2(KEYINPUT82), .A3(new_n205), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n209), .A2(G33), .ZN(new_n458));
  XNOR2_X1  g0258(.A(new_n458), .B(KEYINPUT83), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n258), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n457), .B1(new_n205), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n387), .A2(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n270), .A2(G77), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G97), .A2(G107), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n207), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(KEYINPUT81), .B2(KEYINPUT6), .ZN(new_n466));
  NOR2_X1   g0266(.A1(KEYINPUT81), .A2(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n207), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n205), .A2(KEYINPUT6), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n466), .A2(G20), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n462), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n461), .B1(new_n471), .B2(new_n257), .ZN(new_n472));
  NAND2_X1  g0272(.A1(G33), .A2(G283), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G244), .B(new_n289), .C1(new_n281), .C2(new_n282), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT4), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n283), .A2(new_n287), .A3(G250), .A4(G1698), .ZN(new_n478));
  NOR3_X1   g0278(.A1(new_n476), .A2(new_n439), .A3(G1698), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n283), .A2(new_n287), .A3(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n297), .ZN(new_n482));
  XNOR2_X1  g0282(.A(KEYINPUT5), .B(G41), .ZN(new_n483));
  INV_X1    g0283(.A(G45), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G1), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n483), .A2(G274), .A3(new_n296), .A4(new_n485), .ZN(new_n486));
  AND2_X1   g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  NOR2_X1   g0287(.A1(KEYINPUT5), .A2(G41), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(new_n296), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n486), .B1(new_n490), .B2(new_n226), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n482), .A2(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n493), .A2(G190), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(new_n481), .B2(new_n297), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(G200), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n472), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(G274), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n485), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n225), .B1(new_n484), .B2(G1), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n499), .A2(new_n296), .A3(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n321), .A2(new_n289), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n439), .A2(G1698), .ZN(new_n504));
  OAI211_X1 g0304(.A(new_n503), .B(new_n504), .C1(new_n281), .C2(new_n282), .ZN(new_n505));
  AND2_X1   g0305(.A1(KEYINPUT84), .A2(G116), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT84), .A2(G116), .ZN(new_n507));
  OAI21_X1  g0307(.A(G33), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT85), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n296), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n505), .A2(KEYINPUT85), .A3(new_n508), .ZN(new_n512));
  AOI211_X1 g0312(.A(KEYINPUT86), .B(new_n502), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n509), .A2(new_n510), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n515), .A2(new_n297), .A3(new_n512), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n514), .B1(new_n516), .B2(new_n501), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n407), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n505), .A2(KEYINPUT85), .A3(new_n508), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT85), .B1(new_n505), .B2(new_n508), .ZN(new_n520));
  NOR3_X1   g0320(.A1(new_n519), .A2(new_n520), .A3(new_n296), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT86), .B1(new_n521), .B2(new_n502), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(new_n514), .A3(new_n501), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n522), .A2(new_n336), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n398), .A2(new_n210), .A3(G68), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n347), .A2(new_n205), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n525), .B1(new_n526), .B2(KEYINPUT19), .ZN(new_n527));
  INV_X1    g0327(.A(new_n207), .ZN(new_n528));
  NAND3_X1  g0328(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n528), .A2(new_n224), .B1(new_n210), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n257), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n433), .A2(new_n255), .ZN(new_n532));
  OAI211_X1 g0332(.A(new_n531), .B(new_n532), .C1(new_n460), .C2(new_n433), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n518), .A2(new_n524), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(G200), .B1(new_n513), .B2(new_n517), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n522), .A2(G190), .A3(new_n523), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(new_n532), .ZN(new_n537));
  INV_X1    g0337(.A(new_n460), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n537), .B1(G87), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n536), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n461), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n470), .A2(new_n463), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n542), .B1(G107), .B2(new_n387), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n543), .B2(new_n263), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n495), .A2(new_n336), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n493), .A2(new_n407), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n497), .A2(new_n534), .A3(new_n540), .A4(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n289), .A2(G250), .ZN(new_n549));
  OAI21_X1  g0349(.A(KEYINPUT89), .B1(new_n378), .B2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G294), .ZN(new_n551));
  NOR2_X1   g0351(.A1(new_n268), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n226), .A2(new_n289), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n398), .B2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT89), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n398), .A2(new_n555), .A3(G250), .A4(new_n289), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n550), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n297), .ZN(new_n558));
  INV_X1    g0358(.A(G264), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n490), .A2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n558), .A2(new_n355), .A3(new_n486), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT90), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n558), .A2(new_n486), .A3(new_n561), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n450), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n560), .B1(new_n557), .B2(new_n297), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT90), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n566), .A2(new_n567), .A3(new_n355), .A4(new_n486), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n210), .B(G87), .C1(new_n281), .C2(new_n282), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT22), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n283), .A2(new_n287), .ZN(new_n572));
  OR3_X1    g0372(.A1(new_n224), .A2(KEYINPUT22), .A3(G20), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n571), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n508), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT23), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(new_n210), .B2(G107), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n578));
  AOI22_X1  g0378(.A1(new_n575), .A2(new_n210), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT24), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n574), .A2(new_n579), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n263), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n255), .A2(new_n206), .ZN(new_n585));
  XOR2_X1   g0385(.A(new_n585), .B(KEYINPUT25), .Z(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n206), .B2(new_n460), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n569), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n564), .A2(new_n407), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n566), .A2(new_n336), .A3(new_n486), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n590), .B(new_n591), .C1(new_n584), .C2(new_n587), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT88), .ZN(new_n594));
  INV_X1    g0394(.A(G116), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n594), .B1(new_n460), .B2(new_n595), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n506), .A2(new_n507), .A3(new_n210), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI211_X1 g0398(.A(new_n473), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(KEYINPUT20), .A3(new_n257), .A4(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT20), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n257), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n601), .B1(new_n602), .B2(new_n597), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n254), .A2(G1), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n597), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n459), .A2(KEYINPUT88), .A3(new_n258), .A4(G116), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n596), .A2(new_n604), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G303), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n609), .B1(new_n283), .B2(new_n287), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n559), .A2(G1698), .ZN(new_n611));
  OAI221_X1 g0411(.A(new_n611), .B1(G257), .B2(G1698), .C1(new_n281), .C2(new_n282), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n297), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n489), .A2(G270), .A3(new_n296), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n615), .A2(KEYINPUT87), .A3(new_n486), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT87), .B1(new_n615), .B2(new_n486), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n614), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n608), .B1(G200), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n615), .A2(new_n486), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT87), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n615), .A2(KEYINPUT87), .A3(new_n486), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(G190), .A3(new_n614), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n608), .A2(G169), .A3(new_n618), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT21), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n608), .A2(KEYINPUT21), .A3(G169), .A4(new_n618), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n608), .A2(G179), .A3(new_n614), .A4(new_n624), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n626), .A2(new_n629), .A3(new_n630), .A4(new_n631), .ZN(new_n632));
  NOR3_X1   g0432(.A1(new_n548), .A2(new_n593), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n453), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g0434(.A(new_n634), .B(KEYINPUT91), .Z(G372));
  NAND2_X1  g0435(.A1(new_n516), .A2(new_n501), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n407), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n524), .A2(new_n533), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(G200), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n536), .A2(new_n539), .A3(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n589), .A2(new_n497), .A3(new_n547), .A4(new_n641), .ZN(new_n642));
  AND3_X1   g0442(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n592), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n639), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n646), .A2(new_n638), .A3(new_n641), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT26), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n646), .A2(new_n534), .A3(new_n540), .A4(KEYINPUT26), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n453), .A2(new_n652), .ZN(new_n653));
  AOI22_X1  g0453(.A1(new_n359), .A2(new_n446), .B1(new_n339), .B2(new_n352), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n421), .B1(new_n654), .B2(new_n428), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n314), .B1(new_n655), .B2(new_n311), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n653), .A2(new_n656), .ZN(G369));
  NAND2_X1  g0457(.A1(new_n605), .A2(new_n210), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n608), .A2(new_n663), .ZN(new_n664));
  OR2_X1    g0464(.A1(new_n632), .A2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n643), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(new_n664), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n668), .B(KEYINPUT92), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(G330), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n589), .A2(new_n592), .ZN(new_n672));
  INV_X1    g0472(.A(new_n663), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n588), .B2(new_n673), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n674), .B1(new_n592), .B2(new_n673), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n671), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g0476(.A1(new_n592), .A2(new_n663), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n643), .A2(new_n663), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n672), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n676), .A2(new_n677), .A3(new_n679), .ZN(G399));
  INV_X1    g0480(.A(new_n213), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n681), .A2(G41), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n528), .A2(new_n224), .A3(new_n595), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n682), .A2(new_n209), .A3(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n684), .B1(new_n221), .B2(new_n682), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT28), .Z(new_n686));
  OR3_X1    g0486(.A1(new_n647), .A2(KEYINPUT95), .A3(new_n648), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT95), .B1(new_n647), .B2(new_n648), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n646), .A2(new_n534), .A3(new_n540), .ZN(new_n689));
  OAI211_X1 g0489(.A(new_n687), .B(new_n688), .C1(KEYINPUT26), .C2(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n663), .B1(new_n690), .B2(new_n645), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT29), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT96), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n691), .A2(KEYINPUT96), .A3(KEYINPUT29), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n663), .B1(new_n645), .B2(new_n651), .ZN(new_n696));
  OR2_X1    g0496(.A1(new_n696), .A2(KEYINPUT29), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n694), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n614), .B(G179), .C1(new_n616), .C2(new_n617), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n624), .A2(KEYINPUT93), .A3(G179), .A4(new_n614), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n513), .A2(new_n517), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n495), .A2(new_n566), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n564), .A2(new_n336), .A3(new_n636), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n495), .B1(new_n614), .B2(new_n624), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  AOI21_X1  g0512(.A(G179), .B1(new_n516), .B2(new_n501), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n713), .A2(new_n493), .A3(new_n618), .A4(new_n564), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(KEYINPUT30), .ZN(new_n715));
  NOR3_X1   g0515(.A1(new_n705), .A2(new_n513), .A3(new_n517), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n715), .A2(new_n703), .A3(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n712), .A2(new_n663), .A3(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT31), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT94), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n717), .A4(new_n663), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  AND4_X1   g0523(.A1(new_n497), .A2(new_n534), .A3(new_n540), .A4(new_n547), .ZN(new_n724));
  INV_X1    g0524(.A(new_n632), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n724), .A2(new_n725), .A3(new_n672), .A4(new_n673), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n721), .B1(new_n720), .B2(new_n722), .ZN(new_n728));
  OAI21_X1  g0528(.A(G330), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n698), .A2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n686), .B1(new_n730), .B2(G1), .ZN(G364));
  NOR2_X1   g0531(.A1(new_n254), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n209), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n682), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n671), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G330), .B2(new_n669), .ZN(new_n737));
  NOR2_X1   g0537(.A1(G13), .A2(G33), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(G20), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n216), .B1(G20), .B2(new_n407), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n681), .A2(new_n398), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(G45), .B2(new_n220), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n744), .B1(G45), .B2(new_n249), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n681), .A2(new_n572), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n746), .A2(G355), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(G116), .B2(new_n213), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n742), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n749), .A2(new_n735), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n210), .A2(G179), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G190), .A2(G200), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(G159), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n355), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n336), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G20), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n756), .A2(KEYINPUT32), .B1(new_n760), .B2(new_n205), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n751), .A2(new_n355), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n761), .B1(G107), .B2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n210), .A2(new_n336), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G200), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT98), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n768), .A2(new_n355), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(G190), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n764), .B1(new_n770), .B2(new_n201), .C1(new_n218), .C2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n751), .A2(G190), .A3(G200), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  AOI22_X1  g0575(.A1(new_n756), .A2(KEYINPUT32), .B1(G87), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n765), .A2(new_n752), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n572), .B1(G77), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT97), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n765), .A2(new_n780), .A3(new_n757), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n765), .B2(new_n757), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n776), .B(new_n779), .C1(new_n783), .C2(new_n202), .ZN(new_n784));
  XNOR2_X1  g0584(.A(KEYINPUT33), .B(G317), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G326), .A2(new_n769), .B1(new_n771), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n774), .B(KEYINPUT99), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n609), .B2(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(new_n783), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G322), .ZN(new_n791));
  INV_X1    g0591(.A(new_n753), .ZN(new_n792));
  AOI22_X1  g0592(.A1(G311), .A2(new_n778), .B1(new_n792), .B2(G329), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n763), .A2(G283), .B1(new_n759), .B2(G294), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n791), .A2(new_n572), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  OAI22_X1  g0595(.A1(new_n773), .A2(new_n784), .B1(new_n789), .B2(new_n795), .ZN(new_n796));
  OR2_X1    g0596(.A1(new_n796), .A2(KEYINPUT100), .ZN(new_n797));
  INV_X1    g0597(.A(new_n741), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n798), .B1(new_n796), .B2(KEYINPUT100), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n750), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n740), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n800), .B1(new_n668), .B2(new_n801), .ZN(new_n802));
  AND2_X1   g0602(.A1(new_n737), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(G396));
  NOR3_X1   g0604(.A1(new_n444), .A2(new_n445), .A3(new_n663), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n451), .B1(new_n448), .B2(new_n673), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n805), .B1(new_n806), .B2(new_n447), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n696), .B(new_n807), .ZN(new_n808));
  AOI21_X1  g0608(.A(new_n735), .B1(new_n808), .B2(new_n729), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n729), .B2(new_n808), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n798), .A2(new_n739), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n735), .B1(G77), .B2(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n790), .A2(G143), .B1(G159), .B2(new_n778), .ZN(new_n813));
  INV_X1    g0613(.A(G137), .ZN(new_n814));
  INV_X1    g0614(.A(G150), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n813), .B1(new_n770), .B2(new_n814), .C1(new_n815), .C2(new_n772), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT34), .Z(new_n817));
  INV_X1    g0617(.A(G132), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n398), .B1(new_n753), .B2(new_n818), .C1(new_n760), .C2(new_n202), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(G68), .B2(new_n763), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n201), .B2(new_n788), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n762), .A2(new_n224), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n506), .A2(new_n507), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n572), .B1(new_n823), .B2(new_n753), .C1(new_n824), .C2(new_n777), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n822), .B(new_n825), .C1(G97), .C2(new_n759), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n551), .B2(new_n783), .ZN(new_n827));
  AOI22_X1  g0627(.A1(new_n769), .A2(G303), .B1(G107), .B2(new_n787), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI21_X1  g0629(.A(new_n828), .B1(new_n829), .B2(new_n772), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n817), .A2(new_n821), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n812), .B1(new_n831), .B2(new_n741), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n739), .B2(new_n807), .ZN(new_n833));
  AND2_X1   g0633(.A1(new_n810), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(G384));
  NAND3_X1  g0635(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT35), .ZN(new_n837));
  OAI211_X1 g0637(.A(G116), .B(new_n217), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  XNOR2_X1  g0639(.A(new_n839), .B(KEYINPUT36), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n221), .A2(G77), .A3(new_n365), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n201), .A2(G68), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n209), .B(G13), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n840), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n732), .A2(new_n209), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT38), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n415), .A2(new_n418), .ZN(new_n847));
  INV_X1    g0647(.A(new_n661), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n415), .A2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(KEYINPUT37), .ZN(new_n850));
  NAND4_X1  g0650(.A1(new_n847), .A2(new_n849), .A3(new_n850), .A4(new_n424), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n372), .A2(new_n377), .A3(new_n381), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n853), .A2(KEYINPUT101), .ZN(new_n854));
  AOI21_X1  g0654(.A(KEYINPUT16), .B1(new_n853), .B2(KEYINPUT101), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n383), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n418), .B1(new_n363), .B2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(new_n424), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT102), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n857), .A2(KEYINPUT102), .A3(new_n424), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n848), .B1(new_n856), .B2(new_n363), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n852), .B1(new_n863), .B2(KEYINPUT37), .ZN(new_n864));
  INV_X1    g0664(.A(new_n862), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n865), .B1(new_n420), .B2(new_n428), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n846), .B1(new_n864), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n865), .B1(new_n858), .B2(new_n859), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n850), .B1(new_n869), .B2(new_n861), .ZN(new_n870));
  OAI211_X1 g0670(.A(KEYINPUT38), .B(new_n866), .C1(new_n870), .C2(new_n852), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n652), .A2(new_n673), .A3(new_n807), .ZN(new_n873));
  INV_X1    g0673(.A(new_n805), .ZN(new_n874));
  AND2_X1   g0674(.A1(new_n352), .A2(new_n663), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n353), .A2(new_n359), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n352), .B(new_n663), .C1(new_n339), .C2(new_n358), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n873), .A2(new_n874), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n872), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n421), .B2(new_n848), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n424), .B1(new_n397), .B2(new_n409), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n397), .A2(new_n661), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n884), .A2(KEYINPUT103), .A3(new_n851), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n883), .B1(new_n420), .B2(new_n428), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT103), .B1(new_n884), .B2(new_n851), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n846), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n871), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n893));
  AND2_X1   g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n339), .A2(new_n352), .A3(new_n673), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n881), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n453), .A2(new_n695), .A3(new_n694), .A4(new_n697), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n656), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n453), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT104), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n722), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n673), .B1(new_n707), .B2(new_n711), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n904), .A2(KEYINPUT104), .A3(KEYINPUT31), .A4(new_n717), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n726), .A2(new_n903), .A3(new_n720), .A4(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT105), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AND2_X1   g0708(.A1(new_n903), .A2(new_n905), .ZN(new_n909));
  AOI22_X1  g0709(.A1(new_n633), .A2(new_n673), .B1(new_n719), .B2(new_n718), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n909), .A2(KEYINPUT105), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n901), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  INV_X1    g0712(.A(KEYINPUT40), .ZN(new_n913));
  INV_X1    g0713(.A(new_n878), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n875), .B(new_n358), .C1(new_n339), .C2(new_n352), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n807), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n911), .B2(new_n908), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n872), .A2(new_n913), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n806), .A2(new_n447), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(new_n874), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n920), .B1(new_n877), .B2(new_n878), .ZN(new_n921));
  AOI21_X1  g0721(.A(KEYINPUT105), .B1(new_n909), .B2(new_n910), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n906), .A2(new_n907), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(new_n871), .B2(new_n889), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n918), .B1(new_n925), .B2(new_n913), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n912), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n912), .A2(new_n926), .ZN(new_n928));
  INV_X1    g0728(.A(G330), .ZN(new_n929));
  NOR3_X1   g0729(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n845), .B1(new_n900), .B2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT106), .ZN(new_n932));
  OAI22_X1  g0732(.A1(new_n931), .A2(new_n932), .B1(new_n900), .B2(new_n930), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n931), .A2(new_n932), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n844), .B1(new_n933), .B2(new_n934), .ZN(G367));
  INV_X1    g0735(.A(new_n743), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n742), .B1(new_n213), .B2(new_n433), .C1(new_n936), .C2(new_n245), .ZN(new_n937));
  AND2_X1   g0737(.A1(new_n937), .A2(new_n735), .ZN(new_n938));
  INV_X1    g0738(.A(G317), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n378), .B1(new_n753), .B2(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n760), .A2(new_n206), .B1(new_n762), .B2(new_n205), .ZN(new_n941));
  AOI211_X1 g0741(.A(new_n940), .B(new_n941), .C1(G283), .C2(new_n778), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n774), .A2(new_n824), .ZN(new_n943));
  OAI221_X1 g0743(.A(new_n942), .B1(KEYINPUT46), .B2(new_n943), .C1(new_n609), .C2(new_n783), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n770), .B2(new_n823), .C1(new_n551), .C2(new_n772), .ZN(new_n946));
  OAI22_X1  g0746(.A1(new_n777), .A2(new_n201), .B1(new_n753), .B2(new_n814), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n947), .B1(G58), .B2(new_n775), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n948), .B1(new_n218), .B2(new_n760), .C1(new_n815), .C2(new_n783), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n572), .B1(G77), .B2(new_n763), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT110), .ZN(new_n951));
  INV_X1    g0751(.A(G143), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n951), .B1(new_n770), .B2(new_n952), .C1(new_n754), .C2(new_n772), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n944), .A2(new_n946), .B1(new_n949), .B2(new_n953), .ZN(new_n954));
  XNOR2_X1  g0754(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n954), .B(new_n955), .ZN(new_n956));
  OR2_X1    g0756(.A1(new_n539), .A2(new_n673), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n957), .A2(new_n638), .A3(new_n641), .ZN(new_n958));
  INV_X1    g0758(.A(new_n957), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n958), .A2(KEYINPUT107), .B1(new_n639), .B2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(KEYINPUT107), .B2(new_n958), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT108), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n938), .B1(new_n798), .B2(new_n956), .C1(new_n963), .C2(new_n801), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n679), .A2(new_n677), .ZN(new_n965));
  OAI211_X1 g0765(.A(new_n497), .B(new_n547), .C1(new_n472), .C2(new_n673), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n646), .A2(new_n663), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT44), .Z(new_n970));
  NOR2_X1   g0770(.A1(new_n965), .A2(new_n968), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n973), .B(new_n676), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n679), .B1(new_n675), .B2(new_n678), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT109), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n977), .B1(new_n671), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n670), .B(new_n978), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n979), .B1(new_n980), .B2(new_n977), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n730), .B1(new_n975), .B2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n682), .B(KEYINPUT41), .Z(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n734), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n679), .A2(new_n968), .ZN(new_n986));
  OR2_X1    g0786(.A1(new_n986), .A2(KEYINPUT42), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n547), .B1(new_n966), .B2(new_n592), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n986), .A2(KEYINPUT42), .B1(new_n673), .B2(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(new_n963), .A2(KEYINPUT43), .B1(new_n987), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n963), .A2(KEYINPUT43), .ZN(new_n991));
  XOR2_X1   g0791(.A(new_n990), .B(new_n991), .Z(new_n992));
  OR2_X1    g0792(.A1(new_n676), .A2(new_n968), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n964), .B1(new_n985), .B2(new_n994), .ZN(G387));
  INV_X1    g0795(.A(new_n981), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n734), .ZN(new_n997));
  OR2_X1    g0797(.A1(new_n242), .A2(new_n484), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n998), .A2(new_n743), .B1(new_n683), .B2(new_n746), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n267), .A2(new_n201), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT50), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n484), .B1(new_n218), .B2(new_n291), .ZN(new_n1002));
  NOR3_X1   g0802(.A1(new_n1001), .A2(new_n683), .A3(new_n1002), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n999), .A2(new_n1003), .B1(G107), .B2(new_n213), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n682), .B(new_n734), .C1(new_n1004), .C2(new_n742), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n267), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n754), .A2(new_n770), .B1(new_n772), .B2(new_n1006), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n433), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G97), .A2(new_n763), .B1(new_n759), .B2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n291), .B2(new_n774), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n783), .A2(new_n201), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n398), .B1(new_n753), .B2(new_n815), .C1(new_n218), .C2(new_n777), .ZN(new_n1012));
  NOR4_X1   g0812(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n790), .A2(G317), .B1(G303), .B2(new_n778), .ZN(new_n1014));
  INV_X1    g0814(.A(G322), .ZN(new_n1015));
  OAI221_X1 g0815(.A(new_n1014), .B1(new_n770), .B2(new_n1015), .C1(new_n823), .C2(new_n772), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT48), .ZN(new_n1017));
  OR2_X1    g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n775), .A2(G294), .B1(new_n759), .B2(G283), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT49), .Z(new_n1022));
  OR2_X1    g0822(.A1(new_n1022), .A2(KEYINPUT112), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n398), .B1(new_n792), .B2(G326), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1024), .B1(new_n824), .B2(new_n762), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n1022), .B2(KEYINPUT112), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1013), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1005), .B1(new_n675), .B2(new_n801), .C1(new_n1027), .C2(new_n798), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n997), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n996), .A2(new_n730), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n682), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n996), .A2(new_n730), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G393));
  NAND2_X1  g0833(.A1(new_n974), .A2(new_n734), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n936), .A2(new_n252), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n742), .B1(new_n213), .B2(new_n205), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n735), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n769), .A2(G150), .B1(G159), .B2(new_n790), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT51), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n398), .B1(new_n753), .B2(new_n952), .C1(new_n1006), .C2(new_n777), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n760), .A2(new_n291), .B1(new_n762), .B2(new_n224), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n1040), .B(new_n1041), .C1(G68), .C2(new_n775), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n201), .B2(new_n772), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n769), .A2(G317), .B1(G311), .B2(new_n790), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT52), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n763), .A2(G107), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n829), .B2(new_n774), .C1(new_n760), .C2(new_n824), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n777), .A2(new_n551), .B1(new_n753), .B2(new_n1015), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n288), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n609), .B2(new_n772), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1039), .A2(new_n1043), .B1(new_n1045), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1037), .B1(new_n1051), .B2(new_n741), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n968), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1052), .B1(new_n1053), .B2(new_n801), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1034), .A2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n996), .A2(new_n730), .A3(new_n974), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1056), .A2(new_n682), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1030), .A2(new_n975), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1055), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G390));
  OAI211_X1 g0860(.A(G330), .B(new_n921), .C1(new_n922), .C2(new_n923), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT113), .ZN(new_n1063));
  OAI21_X1  g0863(.A(new_n1063), .B1(new_n879), .B2(new_n896), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n805), .B1(new_n696), .B2(new_n807), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n914), .A2(new_n915), .ZN(new_n1066));
  OAI211_X1 g0866(.A(KEYINPUT113), .B(new_n895), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1068), .B1(new_n892), .B2(new_n893), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n805), .B1(new_n691), .B2(new_n919), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n890), .B(new_n895), .C1(new_n1070), .C2(new_n1066), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1062), .B1(new_n1069), .B2(new_n1072), .ZN(new_n1073));
  OR3_X1    g0873(.A1(new_n729), .A2(new_n920), .A3(new_n1066), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1074), .B(new_n1071), .C1(new_n894), .C2(new_n1068), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n929), .B1(new_n911), .B2(new_n908), .ZN(new_n1078));
  AND2_X1   g0878(.A1(new_n1078), .A2(new_n807), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1066), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n1070), .B(new_n1074), .C1(new_n1079), .C2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1066), .B1(new_n729), .B2(new_n920), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1061), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1065), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1083), .A2(KEYINPUT114), .A3(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(KEYINPUT114), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1081), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n453), .A2(new_n1078), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n898), .A2(new_n656), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1087), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT115), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1077), .A2(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1076), .A2(KEYINPUT115), .A3(new_n1091), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n682), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n892), .A2(new_n893), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1096), .A2(new_n738), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n735), .B1(new_n267), .B2(new_n811), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT116), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n760), .A2(new_n754), .B1(new_n762), .B2(new_n201), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT54), .B(G143), .ZN(new_n1101));
  INV_X1    g0901(.A(G125), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n777), .A2(new_n1101), .B1(new_n753), .B2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g0903(.A1(new_n1100), .A2(new_n1103), .A3(new_n572), .ZN(new_n1104));
  INV_X1    g0904(.A(G128), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1104), .B1(new_n770), .B2(new_n1105), .C1(new_n814), .C2(new_n772), .ZN(new_n1106));
  OR3_X1    g0906(.A1(new_n774), .A2(KEYINPUT53), .A3(new_n815), .ZN(new_n1107));
  OAI21_X1  g0907(.A(KEYINPUT53), .B1(new_n774), .B2(new_n815), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1107), .B(new_n1108), .C1(new_n783), .C2(new_n818), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n790), .A2(G116), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(G97), .A2(new_n778), .B1(new_n792), .B2(G294), .ZN(new_n1111));
  AOI22_X1  g0911(.A1(new_n763), .A2(G68), .B1(new_n759), .B2(G77), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1110), .A2(new_n572), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n769), .A2(G283), .B1(G87), .B2(new_n787), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1114), .B1(new_n206), .B2(new_n772), .ZN(new_n1115));
  OAI22_X1  g0915(.A1(new_n1106), .A2(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1099), .B1(new_n741), .B2(new_n1116), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1097), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1118), .B1(new_n1076), .B2(new_n733), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(KEYINPUT117), .ZN(new_n1120));
  INV_X1    g0920(.A(KEYINPUT117), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1121), .B(new_n1118), .C1(new_n1076), .C2(new_n733), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1095), .A2(new_n1120), .A3(new_n1122), .ZN(G378));
  OAI221_X1 g0923(.A(new_n880), .B1(new_n421), .B2(new_n848), .C1(new_n1096), .C2(new_n895), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n275), .A2(new_n848), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n311), .A2(new_n315), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1127), .B1(new_n311), .B2(new_n315), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1126), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1127), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n316), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(new_n1128), .A3(new_n1125), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n872), .A2(new_n913), .A3(new_n917), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n913), .B1(new_n890), .B2(new_n917), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(G330), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1135), .B1(new_n926), .B2(G330), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1124), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1135), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n890), .A2(new_n917), .ZN(new_n1143));
  AOI21_X1  g0943(.A(KEYINPUT40), .B1(new_n868), .B2(new_n871), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n1143), .A2(KEYINPUT40), .B1(new_n1144), .B2(new_n917), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1142), .B1(new_n1145), .B2(new_n929), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1146), .A2(new_n897), .A3(new_n1138), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1141), .A2(KEYINPUT121), .A3(new_n1147), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT121), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(new_n897), .A3(new_n1149), .A4(new_n1138), .ZN(new_n1150));
  NAND3_X1  g0950(.A1(new_n1148), .A2(new_n734), .A3(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n735), .B1(G50), .B2(new_n811), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n759), .A2(G150), .B1(new_n778), .B2(G137), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n774), .B2(new_n1101), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n1102), .A2(new_n770), .B1(new_n772), .B2(new_n818), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(G128), .C2(new_n790), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1157), .A2(KEYINPUT59), .ZN(new_n1159));
  AOI211_X1 g0959(.A(G33), .B(G41), .C1(new_n792), .C2(G124), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n754), .B2(new_n762), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT119), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1158), .A2(new_n1159), .A3(new_n1162), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n760), .A2(new_n218), .B1(new_n777), .B2(new_n433), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G107), .B2(new_n790), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n770), .B2(new_n595), .ZN(new_n1166));
  OR2_X1    g0966(.A1(new_n398), .A2(G41), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G283), .B2(new_n792), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n202), .B2(new_n762), .C1(new_n291), .C2(new_n774), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT118), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1166), .B(new_n1170), .C1(G97), .C2(new_n771), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1172));
  OAI211_X1 g0972(.A(new_n1167), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n1171), .A2(KEYINPUT58), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n1163), .A2(new_n1172), .A3(new_n1173), .A4(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1152), .B1(new_n1175), .B2(new_n741), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n1135), .B2(new_n739), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT120), .Z(new_n1178));
  AND2_X1   g0978(.A1(new_n1151), .A2(new_n1178), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1073), .A2(new_n1075), .A3(new_n1087), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n1090), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1148), .A2(new_n1181), .A3(new_n1150), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1141), .A2(KEYINPUT122), .A3(new_n1147), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1146), .A2(new_n897), .A3(new_n1186), .A4(new_n1138), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n1181), .A3(KEYINPUT57), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n682), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1179), .B1(new_n1184), .B2(new_n1189), .ZN(G375));
  OAI211_X1 g0990(.A(new_n1089), .B(new_n1081), .C1(new_n1086), .C2(new_n1085), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1091), .A2(new_n1191), .A3(new_n984), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1066), .A2(new_n738), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n735), .B1(G68), .B2(new_n811), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n769), .A2(G132), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n754), .B2(new_n788), .C1(new_n772), .C2(new_n1101), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n398), .B1(new_n777), .B2(new_n815), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1197), .B1(G128), .B2(new_n792), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n763), .A2(G58), .B1(new_n759), .B2(G50), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n814), .C2(new_n783), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n769), .A2(G294), .B1(G97), .B2(new_n787), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1201), .B1(new_n824), .B2(new_n772), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n790), .A2(G283), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G107), .A2(new_n778), .B1(new_n792), .B2(G303), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(G77), .A2(new_n763), .B1(new_n759), .B2(new_n1008), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1203), .A2(new_n572), .A3(new_n1204), .A4(new_n1205), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n1196), .A2(new_n1200), .B1(new_n1202), .B2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1194), .B1(new_n1207), .B2(new_n741), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n1087), .A2(new_n734), .B1(new_n1193), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1192), .A2(new_n1209), .ZN(G381));
  OR2_X1    g1010(.A1(G393), .A2(G396), .ZN(new_n1211));
  OR3_X1    g1011(.A1(new_n1211), .A2(G381), .A3(G384), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1119), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1095), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1059), .B(new_n964), .C1(new_n985), .C2(new_n994), .ZN(new_n1216));
  OR4_X1    g1016(.A1(G375), .A2(new_n1212), .A3(new_n1215), .A4(new_n1216), .ZN(G407));
  NAND2_X1  g1017(.A1(new_n662), .A2(G213), .ZN(new_n1218));
  OR3_X1    g1018(.A1(G375), .A2(new_n1215), .A3(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(G407), .A2(G213), .A3(new_n1219), .ZN(G409));
  INV_X1    g1020(.A(new_n1087), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT60), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1221), .A2(new_n1222), .A3(new_n1089), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1191), .A2(KEYINPUT60), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(new_n1224), .ZN(new_n1225));
  AND2_X1   g1025(.A1(new_n1091), .A2(new_n682), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1225), .A2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1227), .A2(new_n1209), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n834), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1227), .A2(G384), .A3(new_n1209), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n662), .A2(G213), .A3(G2897), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1229), .A2(new_n1230), .A3(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1231), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1227), .B2(new_n1209), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1209), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n834), .B(new_n1235), .C1(new_n1225), .C2(new_n1226), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1232), .A2(new_n1237), .ZN(new_n1238));
  OAI211_X1 g1038(.A(G378), .B(new_n1179), .C1(new_n1184), .C2(new_n1189), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1185), .A2(new_n734), .A3(new_n1187), .ZN(new_n1240));
  OAI211_X1 g1040(.A(new_n1178), .B(new_n1240), .C1(new_n1182), .C2(new_n983), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1214), .A2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1239), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1238), .B1(new_n1243), .B2(new_n1218), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT124), .B1(new_n1244), .B2(KEYINPUT61), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT124), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  AOI22_X1  g1047(.A1(new_n1239), .A2(new_n1242), .B1(G213), .B2(new_n662), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1246), .B(new_n1247), .C1(new_n1248), .C2(new_n1238), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1248), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(KEYINPUT62), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT62), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1248), .A2(new_n1253), .A3(new_n1250), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1245), .A2(new_n1249), .A3(new_n1252), .A4(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(G390), .A2(G387), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1216), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(G393), .A2(G396), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n1211), .A3(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1211), .A2(new_n1258), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1216), .A3(new_n1256), .ZN(new_n1261));
  AND3_X1   g1061(.A1(new_n1259), .A2(KEYINPUT125), .A3(new_n1261), .ZN(new_n1262));
  AOI21_X1  g1062(.A(KEYINPUT125), .B1(new_n1259), .B2(new_n1261), .ZN(new_n1263));
  NOR2_X1   g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1255), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1251), .A2(KEYINPUT63), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT63), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1248), .A2(new_n1267), .A3(new_n1250), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  AND3_X1   g1069(.A1(new_n1259), .A2(new_n1247), .A3(new_n1261), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1244), .A2(KEYINPUT123), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1244), .A2(KEYINPUT123), .ZN(new_n1272));
  OAI211_X1 g1072(.A(new_n1269), .B(new_n1270), .C1(new_n1271), .C2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1265), .A2(new_n1273), .ZN(G405));
  NAND2_X1  g1074(.A1(G375), .A2(new_n1214), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1275), .A2(new_n1239), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1276), .A2(new_n1277), .A3(new_n1250), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1250), .A2(new_n1277), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1275), .A2(new_n1239), .A3(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1264), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(KEYINPUT127), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1278), .A2(new_n1280), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1283), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1284));
  INV_X1    g1084(.A(KEYINPUT127), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1264), .A2(new_n1278), .A3(new_n1285), .A4(new_n1280), .ZN(new_n1286));
  AND3_X1   g1086(.A1(new_n1282), .A2(new_n1284), .A3(new_n1286), .ZN(G402));
endmodule


