

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731;

  XNOR2_X1 U366 ( .A(n408), .B(n441), .ZN(n445) );
  XNOR2_X1 U367 ( .A(n406), .B(G146), .ZN(n469) );
  NAND2_X1 U368 ( .A1(n437), .A2(n436), .ZN(n441) );
  OR2_X1 U369 ( .A1(n463), .A2(n697), .ZN(n364) );
  XOR2_X1 U370 ( .A(G475), .B(n498), .Z(n535) );
  INV_X2 U371 ( .A(G953), .ZN(n718) );
  XNOR2_X2 U372 ( .A(n514), .B(n404), .ZN(n355) );
  NOR2_X1 U373 ( .A1(n685), .A2(n696), .ZN(n376) );
  NOR2_X1 U374 ( .A1(n616), .A2(n696), .ZN(n375) );
  NOR2_X1 U375 ( .A1(n607), .A2(n606), .ZN(n352) );
  NAND2_X2 U376 ( .A1(n358), .A2(n359), .ZN(n525) );
  BUF_X4 U377 ( .A(n646), .Z(n343) );
  NOR2_X2 U378 ( .A1(n401), .A2(n597), .ZN(n579) );
  XNOR2_X2 U379 ( .A(n386), .B(n700), .ZN(n463) );
  INV_X1 U380 ( .A(G125), .ZN(n406) );
  NAND2_X1 U381 ( .A1(n577), .A2(n360), .ZN(n601) );
  AND2_X1 U382 ( .A1(n516), .A2(n426), .ZN(n532) );
  NOR2_X1 U383 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U384 ( .A(n531), .B(KEYINPUT38), .ZN(n657) );
  NAND2_X1 U385 ( .A1(n371), .A2(n656), .ZN(n385) );
  AND2_X1 U386 ( .A1(n370), .A2(n383), .ZN(n359) );
  OR2_X1 U387 ( .A1(n613), .A2(G902), .ZN(n428) );
  XOR2_X2 U388 ( .A(G137), .B(G140), .Z(n369) );
  XNOR2_X1 U389 ( .A(n451), .B(n450), .ZN(n697) );
  XOR2_X1 U390 ( .A(G128), .B(G143), .Z(n344) );
  XNOR2_X1 U391 ( .A(n428), .B(n347), .ZN(n646) );
  NOR2_X1 U392 ( .A1(G953), .A2(G237), .ZN(n485) );
  XNOR2_X1 U393 ( .A(n391), .B(n390), .ZN(n511) );
  INV_X1 U394 ( .A(KEYINPUT105), .ZN(n390) );
  XNOR2_X1 U395 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n567) );
  OR2_X1 U396 ( .A1(G902), .A2(G237), .ZN(n459) );
  INV_X1 U397 ( .A(n518), .ZN(n427) );
  XNOR2_X1 U398 ( .A(n395), .B(n462), .ZN(n394) );
  XNOR2_X1 U399 ( .A(n461), .B(n346), .ZN(n395) );
  XNOR2_X1 U400 ( .A(KEYINPUT71), .B(G113), .ZN(n448) );
  XNOR2_X1 U401 ( .A(n425), .B(n351), .ZN(n555) );
  XNOR2_X1 U402 ( .A(n366), .B(n368), .ZN(n365) );
  NAND2_X1 U403 ( .A1(n504), .A2(G221), .ZN(n368) );
  XNOR2_X1 U404 ( .A(n367), .B(n471), .ZN(n366) );
  NAND2_X1 U405 ( .A1(n397), .A2(n396), .ZN(n420) );
  AND2_X1 U406 ( .A1(n356), .A2(n589), .ZN(n361) );
  INV_X1 U407 ( .A(KEYINPUT46), .ZN(n417) );
  INV_X1 U408 ( .A(KEYINPUT88), .ZN(n578) );
  INV_X1 U409 ( .A(KEYINPUT66), .ZN(n404) );
  XOR2_X1 U410 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n460) );
  AND2_X1 U411 ( .A1(n418), .A2(n416), .ZN(n547) );
  NOR2_X1 U412 ( .A1(n543), .A2(n419), .ZN(n418) );
  XNOR2_X1 U413 ( .A(n542), .B(n417), .ZN(n416) );
  NAND2_X1 U414 ( .A1(n420), .A2(n545), .ZN(n419) );
  INV_X1 U415 ( .A(KEYINPUT67), .ZN(n433) );
  XNOR2_X1 U416 ( .A(n411), .B(n410), .ZN(n602) );
  INV_X1 U417 ( .A(KEYINPUT87), .ZN(n410) );
  NAND2_X1 U418 ( .A1(n413), .A2(n412), .ZN(n411) );
  XNOR2_X1 U419 ( .A(n469), .B(KEYINPUT10), .ZN(n489) );
  XOR2_X1 U420 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n487) );
  XOR2_X1 U421 ( .A(G113), .B(G131), .Z(n484) );
  XNOR2_X1 U422 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U423 ( .A(n369), .B(G104), .ZN(n380) );
  XNOR2_X1 U424 ( .A(KEYINPUT64), .B(G101), .ZN(n442) );
  XNOR2_X1 U425 ( .A(KEYINPUT17), .B(KEYINPUT93), .ZN(n452) );
  XOR2_X1 U426 ( .A(KEYINPUT77), .B(KEYINPUT18), .Z(n453) );
  NAND2_X1 U427 ( .A1(G237), .A2(G234), .ZN(n465) );
  XNOR2_X1 U428 ( .A(n393), .B(KEYINPUT69), .ZN(n523) );
  INV_X1 U429 ( .A(KEYINPUT0), .ZN(n399) );
  NAND2_X1 U430 ( .A1(n407), .A2(G902), .ZN(n383) );
  NAND2_X1 U431 ( .A1(n447), .A2(n382), .ZN(n381) );
  INV_X1 U432 ( .A(G902), .ZN(n382) );
  XNOR2_X1 U433 ( .A(KEYINPUT24), .B(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U434 ( .A(G119), .B(G128), .ZN(n470) );
  XNOR2_X1 U435 ( .A(n475), .B(n405), .ZN(n504) );
  INV_X1 U436 ( .A(KEYINPUT8), .ZN(n405) );
  XOR2_X1 U437 ( .A(G122), .B(G116), .Z(n501) );
  XNOR2_X1 U438 ( .A(G134), .B(G107), .ZN(n500) );
  AND2_X1 U439 ( .A1(n517), .A2(n427), .ZN(n426) );
  INV_X1 U440 ( .A(KEYINPUT6), .ZN(n392) );
  XNOR2_X1 U441 ( .A(n613), .B(n612), .ZN(n614) );
  XNOR2_X1 U442 ( .A(KEYINPUT3), .B(G119), .ZN(n387) );
  XNOR2_X1 U443 ( .A(n448), .B(n389), .ZN(n388) );
  INV_X1 U444 ( .A(G116), .ZN(n389) );
  NOR2_X1 U445 ( .A1(n673), .A2(KEYINPUT83), .ZN(n674) );
  XNOR2_X1 U446 ( .A(n576), .B(KEYINPUT32), .ZN(n729) );
  XNOR2_X1 U447 ( .A(n424), .B(n423), .ZN(n422) );
  INV_X1 U448 ( .A(KEYINPUT60), .ZN(n373) );
  INV_X1 U449 ( .A(n420), .ZN(n637) );
  INV_X1 U450 ( .A(n360), .ZN(n625) );
  NOR2_X1 U451 ( .A1(n553), .A2(n371), .ZN(n345) );
  AND2_X1 U452 ( .A1(n485), .A2(G210), .ZN(n346) );
  XOR2_X1 U453 ( .A(n464), .B(G472), .Z(n347) );
  XNOR2_X1 U454 ( .A(n458), .B(KEYINPUT81), .ZN(n348) );
  AND2_X1 U455 ( .A1(n600), .A2(n599), .ZN(n349) );
  INV_X1 U456 ( .A(n447), .ZN(n407) );
  NOR2_X1 U457 ( .A1(n665), .A2(n401), .ZN(n350) );
  XOR2_X1 U458 ( .A(KEYINPUT86), .B(KEYINPUT39), .Z(n351) );
  NOR2_X1 U459 ( .A1(G952), .A2(n718), .ZN(n696) );
  NOR2_X1 U460 ( .A1(n607), .A2(n606), .ZN(n353) );
  XNOR2_X2 U461 ( .A(n400), .B(n399), .ZN(n354) );
  NOR2_X2 U462 ( .A1(n607), .A2(n606), .ZN(n414) );
  XNOR2_X1 U463 ( .A(n400), .B(n399), .ZN(n593) );
  XNOR2_X1 U464 ( .A(G140), .B(G143), .ZN(n483) );
  XOR2_X1 U465 ( .A(n479), .B(n478), .Z(n356) );
  NOR2_X2 U466 ( .A1(n695), .A2(G902), .ZN(n479) );
  XNOR2_X1 U467 ( .A(n477), .B(KEYINPUT25), .ZN(n478) );
  XNOR2_X1 U468 ( .A(n398), .B(KEYINPUT36), .ZN(n397) );
  NAND2_X1 U469 ( .A1(n358), .A2(n359), .ZN(n357) );
  OR2_X1 U470 ( .A1(n445), .A2(n381), .ZN(n358) );
  INV_X1 U471 ( .A(n572), .ZN(n396) );
  NAND2_X1 U472 ( .A1(n361), .A2(n343), .ZN(n360) );
  BUF_X1 U473 ( .A(n682), .Z(n362) );
  NAND2_X1 U474 ( .A1(n463), .A2(n697), .ZN(n363) );
  NAND2_X1 U475 ( .A1(n364), .A2(n363), .ZN(n377) );
  NOR2_X1 U476 ( .A1(n575), .A2(n647), .ZN(n589) );
  XNOR2_X1 U477 ( .A(n377), .B(n457), .ZN(n682) );
  NAND2_X1 U478 ( .A1(n353), .A2(G475), .ZN(n690) );
  NAND2_X1 U479 ( .A1(n727), .A2(KEYINPUT44), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n712), .B(n365), .ZN(n695) );
  XNOR2_X1 U481 ( .A(n474), .B(n473), .ZN(n367) );
  XNOR2_X1 U482 ( .A(n489), .B(n369), .ZN(n712) );
  NAND2_X1 U483 ( .A1(n445), .A2(n407), .ZN(n370) );
  INV_X1 U484 ( .A(n371), .ZN(n531) );
  XNOR2_X2 U485 ( .A(n415), .B(n348), .ZN(n371) );
  XNOR2_X1 U486 ( .A(n605), .B(KEYINPUT45), .ZN(n403) );
  NAND2_X1 U487 ( .A1(n414), .A2(G210), .ZN(n684) );
  XNOR2_X1 U488 ( .A(n372), .B(KEYINPUT72), .ZN(n604) );
  NAND2_X1 U489 ( .A1(n586), .A2(n587), .ZN(n372) );
  AND2_X2 U490 ( .A1(n403), .A2(n402), .ZN(n673) );
  XNOR2_X2 U491 ( .A(KEYINPUT15), .B(G902), .ZN(n606) );
  NAND2_X1 U492 ( .A1(n430), .A2(n610), .ZN(n611) );
  XNOR2_X1 U493 ( .A(n374), .B(n373), .ZN(G60) );
  NAND2_X1 U494 ( .A1(n691), .A2(n610), .ZN(n374) );
  XNOR2_X1 U495 ( .A(n375), .B(n617), .ZN(G57) );
  XNOR2_X1 U496 ( .A(n380), .B(n440), .ZN(n409) );
  XNOR2_X1 U497 ( .A(n376), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U498 ( .A1(n727), .A2(KEYINPUT44), .ZN(n585) );
  XNOR2_X2 U499 ( .A(n378), .B(KEYINPUT33), .ZN(n401) );
  NOR2_X2 U500 ( .A1(n592), .A2(n588), .ZN(n378) );
  XNOR2_X2 U501 ( .A(n379), .B(KEYINPUT76), .ZN(n592) );
  NAND2_X1 U502 ( .A1(n355), .A2(n647), .ZN(n379) );
  XNOR2_X2 U503 ( .A(n525), .B(KEYINPUT1), .ZN(n647) );
  OR2_X2 U504 ( .A1(n462), .A2(n384), .ZN(n437) );
  INV_X1 U505 ( .A(n449), .ZN(n384) );
  XNOR2_X2 U506 ( .A(n715), .B(G146), .ZN(n462) );
  NAND2_X1 U507 ( .A1(n435), .A2(n434), .ZN(n715) );
  XNOR2_X2 U508 ( .A(n385), .B(KEYINPUT19), .ZN(n563) );
  NOR2_X1 U509 ( .A1(n548), .A2(n385), .ZN(n398) );
  XNOR2_X1 U510 ( .A(n386), .B(n409), .ZN(n408) );
  XNOR2_X2 U511 ( .A(n711), .B(n442), .ZN(n386) );
  XNOR2_X2 U512 ( .A(n388), .B(n387), .ZN(n700) );
  XNOR2_X2 U513 ( .A(n499), .B(KEYINPUT4), .ZN(n711) );
  XNOR2_X2 U514 ( .A(G128), .B(G143), .ZN(n499) );
  NAND2_X2 U515 ( .A1(n563), .A2(n562), .ZN(n400) );
  NOR2_X1 U516 ( .A1(n523), .A2(n588), .ZN(n391) );
  XNOR2_X2 U517 ( .A(n343), .B(n392), .ZN(n588) );
  AND2_X1 U518 ( .A1(n482), .A2(n643), .ZN(n393) );
  XNOR2_X1 U519 ( .A(n463), .B(n394), .ZN(n613) );
  XNOR2_X2 U520 ( .A(n673), .B(KEYINPUT2), .ZN(n607) );
  NOR2_X1 U521 ( .A1(n670), .A2(n401), .ZN(n671) );
  INV_X1 U522 ( .A(n717), .ZN(n402) );
  AND2_X1 U523 ( .A1(n403), .A2(n718), .ZN(n707) );
  NAND2_X1 U524 ( .A1(n355), .A2(n357), .ZN(n596) );
  NOR2_X1 U525 ( .A1(n647), .A2(n355), .ZN(n648) );
  NOR2_X1 U526 ( .A1(n618), .A2(n349), .ZN(n412) );
  NAND2_X1 U527 ( .A1(n414), .A2(G472), .ZN(n615) );
  NAND2_X1 U528 ( .A1(n352), .A2(G469), .ZN(n608) );
  NAND2_X1 U529 ( .A1(n353), .A2(G217), .ZN(n424) );
  NAND2_X1 U530 ( .A1(n352), .A2(G478), .ZN(n692) );
  NAND2_X1 U531 ( .A1(n682), .A2(n606), .ZN(n415) );
  XNOR2_X1 U532 ( .A(n421), .B(KEYINPUT121), .ZN(G66) );
  NAND2_X1 U533 ( .A1(n422), .A2(n610), .ZN(n421) );
  INV_X1 U534 ( .A(n695), .ZN(n423) );
  NAND2_X1 U535 ( .A1(n532), .A2(n657), .ZN(n425) );
  XNOR2_X1 U536 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U537 ( .A(n690), .B(n689), .ZN(n691) );
  INV_X1 U538 ( .A(n729), .ZN(n577) );
  XNOR2_X1 U539 ( .A(n601), .B(n578), .ZN(n587) );
  NOR2_X2 U540 ( .A1(n575), .A2(n574), .ZN(n576) );
  INV_X1 U541 ( .A(n593), .ZN(n597) );
  AND2_X1 U542 ( .A1(n601), .A2(KEYINPUT44), .ZN(n429) );
  INV_X1 U543 ( .A(n696), .ZN(n610) );
  XNOR2_X1 U544 ( .A(n609), .B(n608), .ZN(n430) );
  INV_X1 U545 ( .A(n726), .ZN(n540) );
  NAND2_X1 U546 ( .A1(n541), .A2(n540), .ZN(n542) );
  INV_X1 U547 ( .A(KEYINPUT65), .ZN(n584) );
  XNOR2_X1 U548 ( .A(n460), .B(G137), .ZN(n461) );
  INV_X1 U549 ( .A(KEYINPUT70), .ZN(n446) );
  XNOR2_X1 U550 ( .A(n446), .B(G469), .ZN(n447) );
  XNOR2_X1 U551 ( .A(n615), .B(n614), .ZN(n616) );
  XNOR2_X1 U552 ( .A(KEYINPUT58), .B(KEYINPUT118), .ZN(n444) );
  XNOR2_X2 U553 ( .A(G131), .B(G134), .ZN(n432) );
  INV_X1 U554 ( .A(n432), .ZN(n431) );
  NAND2_X1 U555 ( .A1(n431), .A2(KEYINPUT67), .ZN(n435) );
  NAND2_X1 U556 ( .A1(n433), .A2(n432), .ZN(n434) );
  XOR2_X1 U557 ( .A(G110), .B(G107), .Z(n449) );
  NAND2_X1 U558 ( .A1(n462), .A2(n384), .ZN(n436) );
  NAND2_X1 U559 ( .A1(G227), .A2(n718), .ZN(n439) );
  INV_X1 U560 ( .A(KEYINPUT95), .ZN(n438) );
  XNOR2_X1 U561 ( .A(n445), .B(KEYINPUT57), .ZN(n443) );
  XNOR2_X1 U562 ( .A(n444), .B(n443), .ZN(n609) );
  INV_X1 U563 ( .A(n647), .ZN(n572) );
  XOR2_X1 U564 ( .A(G104), .B(G122), .Z(n490) );
  XOR2_X1 U565 ( .A(n490), .B(KEYINPUT75), .Z(n451) );
  XNOR2_X1 U566 ( .A(n449), .B(KEYINPUT16), .ZN(n450) );
  XNOR2_X1 U567 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U568 ( .A(n469), .B(n454), .Z(n456) );
  NAND2_X1 U569 ( .A1(G224), .A2(n718), .ZN(n455) );
  XNOR2_X1 U570 ( .A(n456), .B(n455), .ZN(n457) );
  NAND2_X1 U571 ( .A1(n459), .A2(G210), .ZN(n458) );
  NAND2_X1 U572 ( .A1(G214), .A2(n459), .ZN(n656) );
  XNOR2_X1 U573 ( .A(KEYINPUT73), .B(KEYINPUT99), .ZN(n464) );
  XNOR2_X1 U574 ( .A(KEYINPUT14), .B(n465), .ZN(n467) );
  NAND2_X1 U575 ( .A1(G902), .A2(n467), .ZN(n558) );
  OR2_X1 U576 ( .A1(n718), .A2(n558), .ZN(n466) );
  NOR2_X1 U577 ( .A1(G900), .A2(n466), .ZN(n468) );
  NAND2_X1 U578 ( .A1(G952), .A2(n467), .ZN(n669) );
  NOR2_X1 U579 ( .A1(G953), .A2(n669), .ZN(n560) );
  NOR2_X1 U580 ( .A1(n468), .A2(n560), .ZN(n518) );
  XNOR2_X1 U581 ( .A(n470), .B(KEYINPUT23), .ZN(n471) );
  INV_X1 U582 ( .A(n472), .ZN(n474) );
  XNOR2_X1 U583 ( .A(G110), .B(KEYINPUT85), .ZN(n473) );
  NAND2_X1 U584 ( .A1(G234), .A2(n718), .ZN(n475) );
  NAND2_X1 U585 ( .A1(G234), .A2(n606), .ZN(n476) );
  XNOR2_X1 U586 ( .A(KEYINPUT20), .B(n476), .ZN(n480) );
  NAND2_X1 U587 ( .A1(n480), .A2(G217), .ZN(n477) );
  XNOR2_X2 U588 ( .A(n479), .B(n478), .ZN(n642) );
  NOR2_X1 U589 ( .A1(n518), .A2(n642), .ZN(n482) );
  NAND2_X1 U590 ( .A1(n480), .A2(G221), .ZN(n481) );
  XOR2_X1 U591 ( .A(KEYINPUT21), .B(n481), .Z(n643) );
  XNOR2_X1 U592 ( .A(n484), .B(n483), .ZN(n495) );
  NAND2_X1 U593 ( .A1(n485), .A2(G214), .ZN(n486) );
  XNOR2_X1 U594 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U595 ( .A(n488), .B(KEYINPUT101), .Z(n493) );
  INV_X1 U596 ( .A(n489), .ZN(n491) );
  XNOR2_X1 U597 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U598 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U599 ( .A(n495), .B(n494), .ZN(n686) );
  NOR2_X1 U600 ( .A1(G902), .A2(n686), .ZN(n497) );
  XNOR2_X1 U601 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n496) );
  XNOR2_X1 U602 ( .A(n497), .B(n496), .ZN(n498) );
  INV_X1 U603 ( .A(n535), .ZN(n512) );
  XNOR2_X1 U604 ( .A(n344), .B(KEYINPUT7), .ZN(n503) );
  XNOR2_X1 U605 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U606 ( .A(n503), .B(n502), .ZN(n508) );
  XOR2_X1 U607 ( .A(KEYINPUT9), .B(KEYINPUT103), .Z(n506) );
  NAND2_X1 U608 ( .A1(G217), .A2(n504), .ZN(n505) );
  XNOR2_X1 U609 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U610 ( .A(n508), .B(n507), .ZN(n693) );
  NOR2_X1 U611 ( .A1(G902), .A2(n693), .ZN(n509) );
  XOR2_X1 U612 ( .A(n509), .B(KEYINPUT104), .Z(n510) );
  XOR2_X1 U613 ( .A(G478), .B(n510), .Z(n534) );
  NAND2_X1 U614 ( .A1(n512), .A2(n534), .ZN(n631) );
  INV_X1 U615 ( .A(n631), .ZN(n513) );
  NAND2_X1 U616 ( .A1(n511), .A2(n513), .ZN(n548) );
  NOR2_X1 U617 ( .A1(n534), .A2(n512), .ZN(n554) );
  NOR2_X1 U618 ( .A1(n513), .A2(n554), .ZN(n662) );
  NAND2_X1 U619 ( .A1(KEYINPUT47), .A2(n662), .ZN(n521) );
  XOR2_X1 U620 ( .A(n643), .B(KEYINPUT97), .Z(n565) );
  NAND2_X1 U621 ( .A1(n565), .A2(n642), .ZN(n514) );
  INV_X1 U622 ( .A(n596), .ZN(n517) );
  INV_X1 U623 ( .A(n343), .ZN(n569) );
  NAND2_X1 U624 ( .A1(n569), .A2(n656), .ZN(n515) );
  XOR2_X1 U625 ( .A(KEYINPUT30), .B(n515), .Z(n516) );
  NOR2_X1 U626 ( .A1(n535), .A2(n534), .ZN(n580) );
  NAND2_X1 U627 ( .A1(n532), .A2(n580), .ZN(n519) );
  NOR2_X1 U628 ( .A1(n519), .A2(n531), .ZN(n520) );
  XNOR2_X1 U629 ( .A(n520), .B(KEYINPUT107), .ZN(n728) );
  NAND2_X1 U630 ( .A1(n521), .A2(n728), .ZN(n522) );
  XOR2_X1 U631 ( .A(KEYINPUT82), .B(n522), .Z(n530) );
  NOR2_X1 U632 ( .A1(n523), .A2(n343), .ZN(n524) );
  XNOR2_X1 U633 ( .A(n524), .B(KEYINPUT28), .ZN(n527) );
  XNOR2_X1 U634 ( .A(n357), .B(KEYINPUT108), .ZN(n526) );
  NAND2_X1 U635 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U636 ( .A(KEYINPUT109), .B(n528), .ZN(n537) );
  NAND2_X1 U637 ( .A1(n563), .A2(n537), .ZN(n629) );
  NAND2_X1 U638 ( .A1(KEYINPUT47), .A2(n629), .ZN(n529) );
  NAND2_X1 U639 ( .A1(n530), .A2(n529), .ZN(n543) );
  NOR2_X1 U640 ( .A1(n631), .A2(n555), .ZN(n533) );
  XNOR2_X1 U641 ( .A(n533), .B(KEYINPUT40), .ZN(n730) );
  INV_X1 U642 ( .A(n730), .ZN(n541) );
  XOR2_X1 U643 ( .A(KEYINPUT110), .B(KEYINPUT42), .Z(n539) );
  NAND2_X1 U644 ( .A1(n535), .A2(n534), .ZN(n660) );
  NAND2_X1 U645 ( .A1(n657), .A2(n656), .ZN(n661) );
  NOR2_X1 U646 ( .A1(n660), .A2(n661), .ZN(n536) );
  XOR2_X1 U647 ( .A(KEYINPUT41), .B(n536), .Z(n641) );
  NAND2_X1 U648 ( .A1(n641), .A2(n537), .ZN(n538) );
  XNOR2_X1 U649 ( .A(n539), .B(n538), .ZN(n726) );
  XOR2_X1 U650 ( .A(n662), .B(KEYINPUT84), .Z(n600) );
  NOR2_X1 U651 ( .A1(n629), .A2(KEYINPUT47), .ZN(n544) );
  NAND2_X1 U652 ( .A1(n600), .A2(n544), .ZN(n545) );
  XNOR2_X1 U653 ( .A(KEYINPUT48), .B(KEYINPUT68), .ZN(n546) );
  XNOR2_X1 U654 ( .A(n547), .B(n546), .ZN(n557) );
  INV_X1 U655 ( .A(n548), .ZN(n549) );
  NAND2_X1 U656 ( .A1(n549), .A2(n656), .ZN(n550) );
  NOR2_X1 U657 ( .A1(n647), .A2(n550), .ZN(n552) );
  XNOR2_X1 U658 ( .A(KEYINPUT106), .B(KEYINPUT43), .ZN(n551) );
  XNOR2_X1 U659 ( .A(n552), .B(n551), .ZN(n553) );
  INV_X1 U660 ( .A(n554), .ZN(n634) );
  NOR2_X1 U661 ( .A1(n555), .A2(n634), .ZN(n639) );
  NOR2_X1 U662 ( .A1(n345), .A2(n639), .ZN(n556) );
  NAND2_X1 U663 ( .A1(n557), .A2(n556), .ZN(n717) );
  INV_X1 U664 ( .A(G898), .ZN(n705) );
  NAND2_X1 U665 ( .A1(G953), .A2(n705), .ZN(n701) );
  NOR2_X1 U666 ( .A1(n558), .A2(n701), .ZN(n559) );
  NOR2_X1 U667 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U668 ( .A(n561), .B(KEYINPUT94), .Z(n562) );
  INV_X1 U669 ( .A(n660), .ZN(n564) );
  AND2_X1 U670 ( .A1(n565), .A2(n564), .ZN(n566) );
  NAND2_X1 U671 ( .A1(n354), .A2(n566), .ZN(n568) );
  XNOR2_X2 U672 ( .A(n568), .B(n567), .ZN(n575) );
  XNOR2_X1 U673 ( .A(KEYINPUT80), .B(n588), .ZN(n570) );
  NAND2_X1 U674 ( .A1(n570), .A2(n356), .ZN(n571) );
  XNOR2_X1 U675 ( .A(n573), .B(KEYINPUT79), .ZN(n574) );
  XNOR2_X1 U676 ( .A(n579), .B(KEYINPUT34), .ZN(n582) );
  XNOR2_X1 U677 ( .A(n580), .B(KEYINPUT78), .ZN(n581) );
  NAND2_X1 U678 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X2 U679 ( .A(n583), .B(KEYINPUT35), .ZN(n727) );
  XNOR2_X1 U680 ( .A(n585), .B(n584), .ZN(n586) );
  INV_X1 U681 ( .A(n588), .ZN(n591) );
  NAND2_X1 U682 ( .A1(n589), .A2(n642), .ZN(n590) );
  NOR2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n618) );
  XOR2_X1 U684 ( .A(KEYINPUT100), .B(KEYINPUT31), .Z(n595) );
  NOR2_X1 U685 ( .A1(n592), .A2(n343), .ZN(n653) );
  NAND2_X1 U686 ( .A1(n653), .A2(n354), .ZN(n594) );
  XNOR2_X1 U687 ( .A(n595), .B(n594), .ZN(n635) );
  NOR2_X1 U688 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U689 ( .A1(n598), .A2(n343), .ZN(n620) );
  NAND2_X1 U690 ( .A1(n635), .A2(n620), .ZN(n599) );
  NOR2_X1 U691 ( .A1(n602), .A2(n429), .ZN(n603) );
  NAND2_X1 U692 ( .A1(n604), .A2(n603), .ZN(n605) );
  XNOR2_X1 U693 ( .A(n611), .B(KEYINPUT119), .ZN(G54) );
  XOR2_X1 U694 ( .A(KEYINPUT62), .B(KEYINPUT91), .Z(n612) );
  XNOR2_X1 U695 ( .A(KEYINPUT89), .B(KEYINPUT63), .ZN(n617) );
  XOR2_X1 U696 ( .A(G101), .B(n618), .Z(G3) );
  NOR2_X1 U697 ( .A1(n631), .A2(n620), .ZN(n619) );
  XOR2_X1 U698 ( .A(G104), .B(n619), .Z(G6) );
  NOR2_X1 U699 ( .A1(n620), .A2(n634), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n622) );
  XNOR2_X1 U701 ( .A(G107), .B(KEYINPUT111), .ZN(n621) );
  XNOR2_X1 U702 ( .A(n622), .B(n621), .ZN(n623) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(G9) );
  XOR2_X1 U704 ( .A(n625), .B(G110), .Z(G12) );
  NOR2_X1 U705 ( .A1(n629), .A2(n634), .ZN(n627) );
  XNOR2_X1 U706 ( .A(KEYINPUT29), .B(KEYINPUT112), .ZN(n626) );
  XNOR2_X1 U707 ( .A(n627), .B(n626), .ZN(n628) );
  XNOR2_X1 U708 ( .A(G128), .B(n628), .ZN(G30) );
  NOR2_X1 U709 ( .A1(n631), .A2(n629), .ZN(n630) );
  XOR2_X1 U710 ( .A(G146), .B(n630), .Z(G48) );
  NOR2_X1 U711 ( .A1(n635), .A2(n631), .ZN(n633) );
  XNOR2_X1 U712 ( .A(G113), .B(KEYINPUT113), .ZN(n632) );
  XNOR2_X1 U713 ( .A(n633), .B(n632), .ZN(G15) );
  NOR2_X1 U714 ( .A1(n635), .A2(n634), .ZN(n636) );
  XOR2_X1 U715 ( .A(G116), .B(n636), .Z(G18) );
  XNOR2_X1 U716 ( .A(G125), .B(n637), .ZN(n638) );
  XNOR2_X1 U717 ( .A(n638), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U718 ( .A(G134), .B(n639), .Z(n640) );
  XNOR2_X1 U719 ( .A(KEYINPUT114), .B(n640), .ZN(G36) );
  XOR2_X1 U720 ( .A(G140), .B(n345), .Z(G42) );
  INV_X1 U721 ( .A(n641), .ZN(n670) );
  NOR2_X1 U722 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U723 ( .A(n644), .B(KEYINPUT49), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n343), .A2(n645), .ZN(n650) );
  XNOR2_X1 U725 ( .A(n648), .B(KEYINPUT50), .ZN(n649) );
  NOR2_X1 U726 ( .A1(n650), .A2(n649), .ZN(n651) );
  XOR2_X1 U727 ( .A(KEYINPUT115), .B(n651), .Z(n652) );
  NOR2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  XOR2_X1 U729 ( .A(KEYINPUT51), .B(n654), .Z(n655) );
  NOR2_X1 U730 ( .A1(n670), .A2(n655), .ZN(n666) );
  NOR2_X1 U731 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U732 ( .A(n658), .B(KEYINPUT116), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n664) );
  NOR2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U735 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U736 ( .A1(n666), .A2(n350), .ZN(n667) );
  XNOR2_X1 U737 ( .A(n667), .B(KEYINPUT52), .ZN(n668) );
  NOR2_X1 U738 ( .A1(n669), .A2(n668), .ZN(n672) );
  NOR2_X1 U739 ( .A1(n672), .A2(n671), .ZN(n676) );
  XOR2_X1 U740 ( .A(KEYINPUT2), .B(n674), .Z(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U742 ( .A1(n677), .A2(G953), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n678), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U744 ( .A(KEYINPUT90), .B(KEYINPUT55), .Z(n680) );
  XNOR2_X1 U745 ( .A(KEYINPUT117), .B(KEYINPUT54), .ZN(n679) );
  XNOR2_X1 U746 ( .A(n680), .B(n679), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n362), .B(n681), .ZN(n683) );
  XNOR2_X1 U748 ( .A(KEYINPUT59), .B(KEYINPUT92), .ZN(n688) );
  XNOR2_X1 U749 ( .A(n686), .B(KEYINPUT120), .ZN(n687) );
  XNOR2_X1 U750 ( .A(n688), .B(n687), .ZN(n689) );
  XNOR2_X1 U751 ( .A(n693), .B(n692), .ZN(n694) );
  NOR2_X1 U752 ( .A1(n696), .A2(n694), .ZN(G63) );
  XNOR2_X1 U753 ( .A(G101), .B(n697), .ZN(n698) );
  XNOR2_X1 U754 ( .A(n698), .B(KEYINPUT123), .ZN(n699) );
  XNOR2_X1 U755 ( .A(n700), .B(n699), .ZN(n702) );
  NAND2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n710) );
  NAND2_X1 U757 ( .A1(G953), .A2(G224), .ZN(n703) );
  XOR2_X1 U758 ( .A(KEYINPUT61), .B(n703), .Z(n704) );
  NOR2_X1 U759 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(KEYINPUT122), .ZN(n708) );
  NOR2_X1 U761 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n710), .B(n709), .ZN(G69) );
  XOR2_X1 U763 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n714) );
  XNOR2_X1 U764 ( .A(n712), .B(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n714), .B(n713), .ZN(n716) );
  XOR2_X1 U766 ( .A(n716), .B(n715), .Z(n720) );
  XNOR2_X1 U767 ( .A(n720), .B(n717), .ZN(n719) );
  NAND2_X1 U768 ( .A1(n719), .A2(n718), .ZN(n725) );
  XNOR2_X1 U769 ( .A(G227), .B(n720), .ZN(n721) );
  NAND2_X1 U770 ( .A1(n721), .A2(G900), .ZN(n722) );
  XNOR2_X1 U771 ( .A(KEYINPUT126), .B(n722), .ZN(n723) );
  NAND2_X1 U772 ( .A1(n723), .A2(G953), .ZN(n724) );
  NAND2_X1 U773 ( .A1(n725), .A2(n724), .ZN(G72) );
  XOR2_X1 U774 ( .A(G137), .B(n726), .Z(G39) );
  XOR2_X1 U775 ( .A(n727), .B(G122), .Z(G24) );
  XNOR2_X1 U776 ( .A(G143), .B(n728), .ZN(G45) );
  XOR2_X1 U777 ( .A(G119), .B(n729), .Z(G21) );
  XNOR2_X1 U778 ( .A(G131), .B(KEYINPUT127), .ZN(n731) );
  XNOR2_X1 U779 ( .A(n731), .B(n730), .ZN(G33) );
endmodule

