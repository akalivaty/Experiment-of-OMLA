//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1306, new_n1307, new_n1308,
    new_n1309, new_n1310, new_n1311, new_n1313, new_n1314, new_n1315,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1412, new_n1413,
    new_n1414, new_n1415, new_n1416, new_n1417;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n218));
  INV_X1    g0018(.A(G226), .ZN(new_n219));
  INV_X1    g0019(.A(G116), .ZN(new_n220));
  INV_X1    g0020(.A(G270), .ZN(new_n221));
  OAI221_X1 g0021(.A(new_n218), .B1(new_n202), .B2(new_n219), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  INV_X1    g0043(.A(G41), .ZN(new_n244));
  INV_X1    g0044(.A(G45), .ZN(new_n245));
  AOI21_X1  g0045(.A(G1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(G33), .A2(G41), .ZN(new_n247));
  NAND3_X1  g0047(.A1(new_n247), .A2(G1), .A3(G13), .ZN(new_n248));
  AND4_X1   g0048(.A1(KEYINPUT64), .A2(new_n246), .A3(new_n248), .A4(G274), .ZN(new_n249));
  INV_X1    g0049(.A(G274), .ZN(new_n250));
  AND2_X1   g0050(.A1(G1), .A2(G13), .ZN(new_n251));
  AOI21_X1  g0051(.A(new_n250), .B1(new_n251), .B2(new_n247), .ZN(new_n252));
  AOI21_X1  g0052(.A(KEYINPUT64), .B1(new_n252), .B2(new_n246), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n249), .A2(new_n253), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n248), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n254), .B1(G226), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT3), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n264), .A2(G223), .B1(new_n267), .B2(G77), .ZN(new_n268));
  INV_X1    g0068(.A(G222), .ZN(new_n269));
  XNOR2_X1  g0069(.A(KEYINPUT3), .B(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n259), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n268), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  AND2_X1   g0072(.A1(G33), .A2(G41), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(new_n215), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n258), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT68), .B1(new_n277), .B2(G190), .ZN(new_n278));
  NAND3_X1  g0078(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n215), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n280), .B1(new_n206), .B2(G20), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n281), .A2(G50), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n282), .B1(G50), .B2(new_n283), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  AOI22_X1  g0085(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT8), .B(G58), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT65), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G58), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(KEYINPUT65), .A3(KEYINPUT8), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n207), .A2(G33), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n286), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n284), .B1(new_n280), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT9), .ZN(new_n296));
  XNOR2_X1  g0096(.A(new_n295), .B(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n276), .A2(G200), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n278), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n299), .A2(KEYINPUT10), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT10), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n278), .A2(new_n297), .A3(new_n301), .A4(new_n298), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(new_n280), .ZN(new_n304));
  INV_X1    g0104(.A(new_n287), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n285), .B1(G20), .B2(G77), .ZN(new_n306));
  XNOR2_X1  g0106(.A(KEYINPUT15), .B(G87), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n307), .A2(new_n293), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n304), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n281), .A2(G77), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(G77), .B2(new_n283), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  XNOR2_X1  g0112(.A(new_n312), .B(KEYINPUT66), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n254), .B1(G244), .B2(new_n257), .ZN(new_n314));
  AOI22_X1  g0114(.A1(new_n264), .A2(G238), .B1(new_n267), .B2(G107), .ZN(new_n315));
  INV_X1    g0115(.A(G232), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n315), .B1(new_n316), .B2(new_n271), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n317), .A2(new_n274), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G200), .ZN(new_n320));
  INV_X1    g0120(.A(G190), .ZN(new_n321));
  OAI211_X1 g0121(.A(new_n313), .B(new_n320), .C1(new_n321), .C2(new_n319), .ZN(new_n322));
  INV_X1    g0122(.A(G169), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n312), .ZN(new_n325));
  INV_X1    g0125(.A(G179), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n314), .A2(new_n326), .A3(new_n318), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT67), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g0131(.A(new_n295), .B1(new_n276), .B2(new_n323), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n332), .B1(G179), .B2(new_n276), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n322), .A2(KEYINPUT67), .A3(new_n328), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n303), .A2(new_n331), .A3(new_n333), .A4(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT73), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n292), .A2(new_n283), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n292), .B2(new_n281), .ZN(new_n338));
  INV_X1    g0138(.A(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(KEYINPUT7), .B1(new_n267), .B2(new_n207), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n262), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n263), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G68), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(G68), .ZN(new_n344));
  NOR2_X1   g0144(.A1(new_n290), .A2(new_n344), .ZN(new_n345));
  OAI21_X1  g0145(.A(G20), .B1(new_n345), .B2(new_n201), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n285), .A2(G159), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n343), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n304), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n341), .A2(KEYINPUT72), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT72), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n267), .A2(new_n354), .A3(KEYINPUT7), .A4(new_n207), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n262), .A2(new_n207), .A3(new_n263), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT7), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(G68), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n346), .A2(KEYINPUT16), .A3(new_n347), .ZN(new_n361));
  INV_X1    g0161(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n339), .B1(new_n352), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G200), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n248), .A2(G232), .A3(new_n255), .ZN(new_n366));
  NOR2_X1   g0166(.A1(G223), .A2(G1698), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n367), .B1(new_n219), .B2(G1698), .ZN(new_n368));
  AOI22_X1  g0168(.A1(new_n368), .A2(new_n270), .B1(G33), .B2(G87), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n366), .B1(new_n369), .B2(new_n248), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n365), .B1(new_n370), .B2(new_n254), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n219), .A2(G1698), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n372), .B1(G223), .B2(G1698), .ZN(new_n373));
  INV_X1    g0173(.A(G87), .ZN(new_n374));
  OAI22_X1  g0174(.A1(new_n373), .A2(new_n267), .B1(new_n261), .B2(new_n374), .ZN(new_n375));
  AOI22_X1  g0175(.A1(new_n375), .A2(new_n274), .B1(G232), .B2(new_n257), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT64), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n248), .A2(G274), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n377), .B1(new_n378), .B2(new_n255), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n252), .A2(KEYINPUT64), .A3(new_n246), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n376), .A2(new_n321), .A3(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n371), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(KEYINPUT17), .B1(new_n364), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n344), .B1(new_n358), .B2(new_n341), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n351), .B1(new_n385), .B2(new_n348), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n363), .A2(new_n280), .A3(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n387), .A2(new_n383), .A3(KEYINPUT17), .A4(new_n338), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n336), .B1(new_n384), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n386), .A2(new_n280), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n361), .B1(new_n359), .B2(G68), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n338), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT18), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n376), .A2(G179), .A3(new_n381), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n370), .A2(new_n254), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n395), .B1(new_n396), .B2(new_n323), .ZN(new_n397));
  AND3_X1   g0197(.A1(new_n393), .A2(new_n394), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n394), .B1(new_n393), .B2(new_n397), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT17), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n371), .A2(new_n382), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n393), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n403), .A2(KEYINPUT73), .A3(new_n388), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n390), .A2(new_n400), .A3(new_n404), .ZN(new_n405));
  XOR2_X1   g0205(.A(KEYINPUT70), .B(KEYINPUT13), .Z(new_n406));
  NAND2_X1  g0206(.A1(new_n219), .A2(new_n259), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n316), .A2(G1698), .ZN(new_n408));
  OAI211_X1 g0208(.A(new_n407), .B(new_n408), .C1(new_n265), .C2(new_n266), .ZN(new_n409));
  NAND2_X1  g0209(.A1(G33), .A2(G97), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n274), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT69), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n248), .B1(new_n409), .B2(new_n410), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT69), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G238), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n256), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n379), .B2(new_n380), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n406), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n414), .A2(new_n415), .ZN(new_n422));
  AOI211_X1 g0222(.A(KEYINPUT69), .B(new_n248), .C1(new_n409), .C2(new_n410), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n420), .B(new_n406), .C1(new_n422), .C2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(G169), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n426), .A2(KEYINPUT14), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n420), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n428), .A2(KEYINPUT71), .A3(KEYINPUT13), .ZN(new_n429));
  AOI21_X1  g0229(.A(KEYINPUT71), .B1(new_n428), .B2(KEYINPUT13), .ZN(new_n430));
  OAI211_X1 g0230(.A(G179), .B(new_n424), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n406), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(new_n424), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT14), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n434), .A2(new_n435), .A3(G169), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n427), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n281), .A2(G68), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT12), .ZN(new_n439));
  INV_X1    g0239(.A(new_n283), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(new_n344), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n283), .A2(KEYINPUT12), .A3(G68), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n438), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT11), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n285), .A2(G50), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n445), .B1(new_n207), .B2(G68), .ZN(new_n446));
  INV_X1    g0246(.A(G77), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n293), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n280), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n443), .B1(new_n444), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n450), .B1(new_n444), .B2(new_n449), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n437), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n451), .B1(new_n434), .B2(G200), .ZN(new_n453));
  OAI211_X1 g0253(.A(G190), .B(new_n424), .C1(new_n429), .C2(new_n430), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(G244), .B(new_n259), .C1(new_n265), .C2(new_n266), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT75), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  OR2_X1    g0261(.A1(new_n457), .A2(new_n458), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n457), .A2(KEYINPUT75), .A3(new_n458), .ZN(new_n463));
  OAI211_X1 g0263(.A(G250), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n464));
  NAND2_X1  g0264(.A1(G33), .A2(G283), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g0266(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(new_n274), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n245), .A2(G1), .ZN(new_n469));
  AND2_X1   g0269(.A1(KEYINPUT5), .A2(G41), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n472), .A2(G257), .A3(new_n248), .ZN(new_n473));
  XNOR2_X1  g0273(.A(KEYINPUT5), .B(G41), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n252), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT76), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n473), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n476), .B1(new_n473), .B2(new_n475), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n468), .A2(new_n480), .A3(new_n321), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n465), .B(new_n464), .C1(new_n457), .C2(new_n458), .ZN(new_n482));
  AOI21_X1  g0282(.A(KEYINPUT75), .B1(new_n457), .B2(new_n458), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n248), .B1(new_n484), .B2(new_n463), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n473), .A2(new_n475), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT76), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n477), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n481), .B1(new_n489), .B2(G200), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n283), .A2(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n261), .A2(G1), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n440), .A2(new_n280), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(G97), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(G107), .B1(new_n340), .B2(new_n342), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  AND2_X1   g0297(.A1(G97), .A2(G107), .ZN(new_n498));
  NOR2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n497), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G107), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT6), .A3(G97), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g0303(.A1(new_n503), .A2(G20), .B1(G77), .B2(new_n285), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n280), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT74), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n505), .A2(KEYINPUT74), .A3(new_n280), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n495), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n490), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT74), .B1(new_n505), .B2(new_n280), .ZN(new_n512));
  AOI211_X1 g0312(.A(new_n507), .B(new_n304), .C1(new_n496), .C2(new_n504), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n494), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n468), .A2(new_n480), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(new_n323), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n468), .A2(new_n480), .A3(new_n326), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT19), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n207), .B1(new_n410), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n499), .A2(new_n374), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n207), .B(G68), .C1(new_n265), .C2(new_n266), .ZN(new_n523));
  INV_X1    g0323(.A(G97), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n519), .B1(new_n293), .B2(new_n524), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n522), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  AOI22_X1  g0326(.A1(new_n526), .A2(new_n280), .B1(new_n440), .B2(new_n307), .ZN(new_n527));
  INV_X1    g0327(.A(new_n307), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n493), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  OAI211_X1 g0330(.A(G244), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n531));
  OAI211_X1 g0331(.A(G238), .B(new_n259), .C1(new_n265), .C2(new_n266), .ZN(new_n532));
  NAND2_X1  g0332(.A1(G33), .A2(G116), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n274), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n248), .A2(G274), .A3(new_n469), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n206), .A2(G45), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(G250), .C1(new_n273), .C2(new_n215), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n535), .A2(new_n326), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n539), .B1(new_n534), .B2(new_n274), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n530), .B(new_n541), .C1(G169), .C2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n542), .A2(KEYINPUT78), .A3(G190), .ZN(new_n544));
  AOI21_X1  g0344(.A(KEYINPUT78), .B1(new_n542), .B2(G190), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n526), .A2(new_n280), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n307), .A2(new_n440), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n493), .A2(G87), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n547), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT77), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n550), .B(new_n551), .C1(new_n365), .C2(new_n542), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n527), .B(new_n549), .C1(new_n542), .C2(new_n365), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT77), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n546), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n511), .A2(new_n518), .A3(new_n543), .A4(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  OAI211_X1 g0357(.A(G264), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(KEYINPUT79), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT79), .ZN(new_n560));
  NAND4_X1  g0360(.A1(new_n270), .A2(new_n560), .A3(G264), .A4(G1698), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n267), .A2(G303), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n270), .A2(G257), .A3(new_n259), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n559), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(new_n274), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n472), .A2(new_n248), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n475), .B1(new_n566), .B2(new_n221), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  AOI22_X1  g0369(.A1(new_n279), .A2(new_n215), .B1(G20), .B2(new_n220), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n465), .B(new_n207), .C1(G33), .C2(new_n524), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT20), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(KEYINPUT20), .A3(new_n571), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n283), .A2(G116), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n493), .B2(G116), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n323), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n569), .A2(new_n579), .A3(KEYINPUT21), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT80), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n569), .A2(new_n579), .A3(KEYINPUT80), .A4(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n569), .A2(new_n579), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  AND3_X1   g0386(.A1(new_n565), .A2(G179), .A3(new_n568), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n576), .A2(new_n578), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n585), .A2(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n588), .B1(new_n569), .B2(G200), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n590), .B1(new_n321), .B2(new_n569), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n584), .A2(new_n589), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  OAI211_X1 g0393(.A(G257), .B(G1698), .C1(new_n265), .C2(new_n266), .ZN(new_n594));
  OAI211_X1 g0394(.A(G250), .B(new_n259), .C1(new_n265), .C2(new_n266), .ZN(new_n595));
  NAND2_X1  g0395(.A1(G33), .A2(G294), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n274), .B1(new_n469), .B2(new_n474), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n274), .A2(new_n597), .B1(new_n598), .B2(G264), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n475), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(G169), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n597), .A2(new_n274), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n598), .A2(G264), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT82), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n599), .A2(KEYINPUT82), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n606), .A2(new_n607), .A3(G179), .A4(new_n475), .ZN(new_n608));
  NOR2_X1   g0408(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n270), .A2(new_n207), .A3(G87), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n610), .A2(KEYINPUT22), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT22), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n270), .A2(new_n612), .A3(new_n207), .A4(G87), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g0414(.A(KEYINPUT23), .B1(new_n207), .B2(G107), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT23), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n616), .A2(new_n501), .A3(G20), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n618));
  NAND2_X1  g0418(.A1(KEYINPUT81), .A2(KEYINPUT24), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n615), .A2(new_n617), .A3(new_n618), .A4(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n609), .B1(new_n614), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n609), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n623), .B(new_n620), .C1(new_n611), .C2(new_n613), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n280), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT25), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n283), .A2(new_n626), .A3(G107), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n626), .B1(new_n283), .B2(G107), .ZN(new_n629));
  AOI22_X1  g0429(.A1(G107), .A2(new_n493), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n601), .A2(new_n608), .B1(new_n625), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(new_n630), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n614), .A2(new_n621), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n623), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n614), .A2(new_n609), .A3(new_n621), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n632), .B1(new_n636), .B2(new_n280), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n606), .A2(new_n607), .A3(new_n475), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n365), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n602), .A2(new_n603), .A3(new_n321), .A4(new_n475), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT83), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n631), .B1(new_n637), .B2(new_n642), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n557), .A2(new_n593), .A3(new_n643), .ZN(new_n644));
  NOR4_X1   g0444(.A1(new_n335), .A2(new_n405), .A3(new_n456), .A4(new_n644), .ZN(G372));
  NOR3_X1   g0445(.A1(new_n335), .A2(new_n405), .A3(new_n456), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n541), .B1(G169), .B2(new_n542), .ZN(new_n647));
  INV_X1    g0447(.A(new_n530), .ZN(new_n648));
  AND2_X1   g0448(.A1(new_n542), .A2(G190), .ZN(new_n649));
  OAI22_X1  g0449(.A1(new_n647), .A2(new_n648), .B1(new_n553), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT84), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI211_X1 g0452(.A(new_n543), .B(KEYINPUT84), .C1(new_n553), .C2(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AND3_X1   g0454(.A1(new_n602), .A2(KEYINPUT82), .A3(new_n603), .ZN(new_n655));
  AOI21_X1  g0455(.A(KEYINPUT82), .B1(new_n602), .B2(new_n603), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g0457(.A(G200), .B1(new_n657), .B2(new_n475), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT83), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n640), .B(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n637), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n654), .A2(new_n661), .A3(new_n518), .A4(new_n511), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n608), .A2(new_n601), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n625), .A2(new_n630), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n665), .A2(new_n584), .A3(new_n589), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n543), .B1(new_n662), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n668));
  AOI21_X1  g0468(.A(KEYINPUT26), .B1(new_n654), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n555), .A2(new_n543), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT26), .ZN(new_n671));
  NOR3_X1   g0471(.A1(new_n670), .A2(new_n518), .A3(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  OR2_X1    g0473(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n646), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n328), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n455), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n452), .A2(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n390), .A2(new_n404), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT85), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n398), .B2(new_n399), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n393), .A2(new_n397), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT18), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(KEYINPUT85), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n680), .A2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n303), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n675), .A2(new_n333), .A3(new_n689), .ZN(G369));
  NAND3_X1  g0490(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(G213), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n696), .B1(new_n584), .B2(new_n589), .ZN(new_n697));
  INV_X1    g0497(.A(new_n696), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n643), .A2(new_n697), .B1(new_n631), .B2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(G330), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n584), .A2(new_n589), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n588), .A2(new_n696), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n584), .A2(new_n589), .A3(new_n591), .A4(new_n702), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n700), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT86), .ZN(new_n707));
  XNOR2_X1  g0507(.A(new_n706), .B(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n643), .B1(new_n637), .B2(new_n698), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n665), .B2(new_n698), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT87), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n705), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n707), .B1(new_n712), .B2(G330), .ZN(new_n713));
  AOI211_X1 g0513(.A(KEYINPUT86), .B(new_n700), .C1(new_n704), .C2(new_n705), .ZN(new_n714));
  OAI211_X1 g0514(.A(KEYINPUT87), .B(new_n710), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g0516(.A(new_n699), .B1(new_n711), .B2(new_n716), .ZN(G399));
  INV_X1    g0517(.A(new_n210), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(G41), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n521), .A2(G116), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n720), .A2(G1), .A3(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(new_n213), .B2(new_n720), .ZN(new_n723));
  XNOR2_X1  g0523(.A(new_n723), .B(KEYINPUT28), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n569), .A2(new_n326), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n489), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n535), .A2(new_n540), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT89), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n542), .A2(KEYINPUT89), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND4_X1  g0531(.A1(new_n726), .A2(KEYINPUT90), .A3(new_n638), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g0532(.A(G179), .B1(new_n565), .B2(new_n568), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n638), .A2(new_n515), .A3(new_n731), .A4(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT90), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(KEYINPUT91), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT88), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n567), .B1(new_n564), .B2(new_n274), .ZN(new_n741));
  NAND4_X1  g0541(.A1(new_n468), .A2(new_n480), .A3(new_n741), .A4(G179), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n606), .A2(new_n607), .A3(new_n542), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n740), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR3_X1   g0544(.A1(new_n655), .A2(new_n656), .A3(new_n727), .ZN(new_n745));
  INV_X1    g0545(.A(new_n740), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n745), .A2(new_n489), .A3(new_n587), .A4(new_n746), .ZN(new_n747));
  AND2_X1   g0547(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  AND3_X1   g0548(.A1(new_n737), .A2(new_n738), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n738), .B1(new_n737), .B2(new_n748), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n696), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(KEYINPUT31), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n557), .A2(new_n593), .A3(new_n643), .A4(new_n698), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n748), .A2(new_n734), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n698), .A2(new_n752), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  AND2_X1   g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n700), .B1(new_n753), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n668), .A2(new_n671), .A3(new_n543), .A4(new_n555), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n518), .B1(new_n652), .B2(new_n653), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n760), .B1(new_n761), .B2(new_n671), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n698), .B1(new_n667), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT29), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT29), .ZN(new_n765));
  OAI211_X1 g0565(.A(new_n765), .B(new_n698), .C1(new_n667), .C2(new_n673), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n724), .B1(new_n768), .B2(G1), .ZN(new_n769));
  XNOR2_X1  g0569(.A(new_n769), .B(KEYINPUT92), .ZN(G364));
  NOR2_X1   g0570(.A1(new_n712), .A2(G330), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(KEYINPUT93), .ZN(new_n772));
  INV_X1    g0572(.A(G13), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n206), .B1(new_n774), .B2(G45), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n719), .A2(new_n776), .ZN(new_n777));
  OR3_X1    g0577(.A1(new_n772), .A2(new_n708), .A3(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n718), .A2(new_n267), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n779), .A2(G355), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G116), .B2(new_n210), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n718), .A2(new_n270), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n783), .B1(new_n245), .B2(new_n214), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n239), .A2(new_n245), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(G13), .A2(G33), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(G20), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n215), .B1(G20), .B2(new_n323), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n791), .B(KEYINPUT94), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n777), .B1(new_n786), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n207), .A2(G179), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G190), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n270), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G283), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n794), .A2(new_n321), .A3(G200), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n798), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n321), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n326), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(G20), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(G294), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n794), .A2(G190), .A3(G200), .ZN(new_n807));
  INV_X1    g0607(.A(G303), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n801), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G311), .ZN(new_n811));
  NAND2_X1  g0611(.A1(G20), .A2(G179), .ZN(new_n812));
  XNOR2_X1  g0612(.A(new_n812), .B(KEYINPUT95), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(new_n795), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n810), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT98), .ZN(new_n816));
  AND2_X1   g0616(.A1(new_n813), .A2(new_n802), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n817), .A2(G322), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n813), .A2(G200), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n321), .ZN(new_n821));
  XOR2_X1   g0621(.A(KEYINPUT33), .B(G317), .Z(new_n822));
  OAI21_X1  g0622(.A(new_n818), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n815), .B1(new_n816), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G326), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n820), .A2(KEYINPUT97), .A3(G190), .ZN(new_n826));
  INV_X1    g0626(.A(KEYINPUT97), .ZN(new_n827));
  OAI21_X1  g0627(.A(new_n827), .B1(new_n819), .B2(new_n321), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n824), .B1(new_n816), .B2(new_n823), .C1(new_n825), .C2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(G159), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n796), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT32), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n270), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n800), .A2(new_n501), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n834), .B2(new_n833), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n837), .B1(new_n374), .B2(new_n807), .C1(new_n524), .C2(new_n805), .ZN(new_n838));
  INV_X1    g0638(.A(new_n821), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n835), .B(new_n838), .C1(G68), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n814), .ZN(new_n841));
  AOI22_X1  g0641(.A1(G77), .A2(new_n841), .B1(new_n817), .B2(G58), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT96), .ZN(new_n843));
  OAI211_X1 g0643(.A(new_n840), .B(new_n843), .C1(new_n202), .C2(new_n830), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n831), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n793), .B1(new_n845), .B2(new_n790), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n789), .B(KEYINPUT99), .Z(new_n847));
  OAI21_X1  g0647(.A(new_n846), .B1(new_n712), .B2(new_n847), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT100), .Z(new_n849));
  NAND2_X1  g0649(.A1(new_n778), .A2(new_n849), .ZN(G396));
  NAND2_X1  g0650(.A1(new_n328), .A2(KEYINPUT102), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n324), .A2(new_n852), .A3(new_n325), .A4(new_n327), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n322), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n698), .B(new_n854), .C1(new_n667), .C2(new_n673), .ZN(new_n855));
  AND2_X1   g0655(.A1(new_n674), .A2(new_n698), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n325), .A2(new_n696), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n322), .A2(new_n851), .A3(new_n857), .A4(new_n853), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n676), .A2(new_n696), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n856), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n759), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n777), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(new_n862), .B2(new_n861), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n790), .A2(new_n787), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n777), .B1(G77), .B2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n817), .ZN(new_n867));
  OAI22_X1  g0667(.A1(new_n867), .A2(new_n806), .B1(new_n220), .B2(new_n814), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n267), .B1(new_n796), .B2(new_n811), .C1(new_n805), .C2(new_n524), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n800), .A2(new_n374), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n807), .A2(new_n501), .ZN(new_n871));
  NOR4_X1   g0671(.A1(new_n868), .A2(new_n869), .A3(new_n870), .A4(new_n871), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n872), .B1(new_n799), .B2(new_n821), .C1(new_n830), .C2(new_n808), .ZN(new_n873));
  XNOR2_X1  g0673(.A(new_n873), .B(KEYINPUT101), .ZN(new_n874));
  AOI22_X1  g0674(.A1(G159), .A2(new_n841), .B1(new_n817), .B2(G143), .ZN(new_n875));
  INV_X1    g0675(.A(G150), .ZN(new_n876));
  INV_X1    g0676(.A(G137), .ZN(new_n877));
  OAI221_X1 g0677(.A(new_n875), .B1(new_n876), .B2(new_n821), .C1(new_n830), .C2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT34), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(G132), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n270), .B1(new_n796), .B2(new_n881), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n805), .A2(new_n290), .B1(new_n807), .B2(new_n202), .ZN(new_n883));
  INV_X1    g0683(.A(new_n800), .ZN(new_n884));
  AOI211_X1 g0684(.A(new_n882), .B(new_n883), .C1(G68), .C2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n878), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(KEYINPUT34), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n874), .B1(new_n880), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n866), .B1(new_n888), .B2(new_n790), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n788), .B2(new_n860), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n864), .A2(new_n890), .ZN(G384));
  NOR2_X1   g0691(.A1(new_n774), .A2(new_n206), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n364), .A2(new_n383), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n360), .A2(new_n349), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(KEYINPUT103), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n348), .B1(new_n359), .B2(G68), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT103), .ZN(new_n897));
  AOI21_X1  g0697(.A(KEYINPUT16), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g0699(.A1(new_n392), .A2(new_n304), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n339), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(new_n397), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n893), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n901), .A2(new_n694), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AND2_X1   g0705(.A1(new_n893), .A2(new_n683), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  INV_X1    g0707(.A(new_n694), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n393), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n906), .A2(new_n907), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n905), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n405), .A2(new_n904), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n913));
  AOI22_X1  g0713(.A1(new_n905), .A2(new_n910), .B1(new_n405), .B2(new_n904), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n914), .B2(KEYINPUT38), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n756), .B1(new_n749), .B2(new_n750), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n734), .B(KEYINPUT90), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n744), .A2(new_n747), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT91), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n737), .A2(new_n738), .A3(new_n748), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n698), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n754), .B(new_n916), .C1(new_n921), .C2(KEYINPUT31), .ZN(new_n922));
  INV_X1    g0722(.A(new_n860), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n451), .A2(new_n696), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n452), .A2(new_n455), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n455), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n451), .B(new_n696), .C1(new_n926), .C2(new_n437), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n923), .B1(new_n925), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n915), .A2(new_n922), .A3(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT40), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(KEYINPUT104), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n907), .B1(new_n909), .B2(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n906), .A2(new_n909), .A3(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n364), .A2(new_n694), .ZN(new_n935));
  OAI21_X1  g0735(.A(KEYINPUT37), .B1(new_n935), .B2(KEYINPUT104), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n893), .A2(new_n683), .A3(new_n909), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n934), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT105), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n384), .B2(new_n389), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n403), .A2(KEYINPUT105), .A3(new_n388), .ZN(new_n942));
  NOR3_X1   g0742(.A1(new_n398), .A2(new_n399), .A3(new_n681), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT85), .B1(new_n684), .B2(new_n685), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n939), .B1(new_n945), .B2(new_n935), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n913), .B1(new_n946), .B2(KEYINPUT38), .ZN(new_n947));
  NAND4_X1  g0747(.A1(new_n947), .A2(new_n922), .A3(KEYINPUT40), .A4(new_n928), .ZN(new_n948));
  AND2_X1   g0748(.A1(new_n931), .A2(new_n948), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n922), .A2(new_n646), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n700), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  INV_X1    g0752(.A(KEYINPUT39), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n943), .A2(new_n944), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n941), .A2(new_n942), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n935), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n939), .ZN(new_n957));
  AOI21_X1  g0757(.A(KEYINPUT38), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n911), .A2(new_n912), .A3(KEYINPUT38), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n953), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n452), .A2(new_n696), .ZN(new_n961));
  OAI211_X1 g0761(.A(new_n913), .B(KEYINPUT39), .C1(KEYINPUT38), .C2(new_n914), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g0763(.A1(new_n925), .A2(new_n927), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n851), .A2(new_n853), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n698), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n964), .B1(new_n855), .B2(new_n966), .ZN(new_n967));
  AOI22_X1  g0767(.A1(new_n967), .A2(new_n915), .B1(new_n954), .B2(new_n694), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n689), .A2(new_n333), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n767), .B2(new_n646), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n969), .B(new_n971), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n892), .B1(new_n952), .B2(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n973), .B1(new_n972), .B2(new_n952), .ZN(new_n974));
  OR2_X1    g0774(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n503), .A2(KEYINPUT35), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n975), .A2(G116), .A3(new_n216), .A4(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT36), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n345), .A2(new_n213), .A3(new_n447), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n344), .A2(G50), .ZN(new_n980));
  OAI211_X1 g0780(.A(G1), .B(new_n773), .C1(new_n979), .C2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(G367));
  OR2_X1    g0782(.A1(new_n550), .A2(new_n698), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n543), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n984), .B(KEYINPUT106), .Z(new_n985));
  NAND2_X1  g0785(.A1(new_n654), .A2(new_n983), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(KEYINPUT107), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(new_n847), .ZN(new_n990));
  INV_X1    g0790(.A(new_n792), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n991), .B1(new_n210), .B2(new_n307), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n783), .A2(new_n235), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n777), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n830), .A2(new_n811), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n839), .A2(G294), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n807), .A2(new_n220), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n997), .A2(KEYINPUT46), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n998), .B1(G283), .B2(new_n841), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n817), .A2(G303), .B1(KEYINPUT46), .B2(new_n997), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n800), .A2(new_n524), .ZN(new_n1001));
  XOR2_X1   g0801(.A(KEYINPUT109), .B(G317), .Z(new_n1002));
  OAI21_X1  g0802(.A(new_n267), .B1(new_n1002), .B2(new_n796), .ZN(new_n1003));
  AOI211_X1 g0803(.A(new_n1001), .B(new_n1003), .C1(G107), .C2(new_n804), .ZN(new_n1004));
  NAND4_X1  g0804(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .A4(new_n1004), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n270), .B1(new_n796), .B2(new_n877), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n290), .A2(new_n807), .B1(new_n800), .B2(new_n447), .ZN(new_n1007));
  AOI211_X1 g0807(.A(new_n1006), .B(new_n1007), .C1(G68), .C2(new_n804), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G50), .A2(new_n841), .B1(new_n817), .B2(G150), .ZN(new_n1009));
  OAI211_X1 g0809(.A(new_n1008), .B(new_n1009), .C1(new_n832), .C2(new_n821), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n829), .A2(G143), .ZN(new_n1011));
  OAI22_X1  g0811(.A1(new_n995), .A2(new_n1005), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT47), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n994), .B1(new_n1013), .B2(new_n790), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n990), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n701), .A2(new_n698), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n661), .A2(new_n665), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1017), .A2(new_n1018), .B1(new_n665), .B2(new_n696), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n668), .A2(new_n696), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n514), .A2(new_n696), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n511), .A2(new_n518), .A3(new_n1021), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1016), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1019), .A2(KEYINPUT44), .A3(new_n1023), .ZN(new_n1028));
  INV_X1    g0828(.A(KEYINPUT44), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n699), .B2(new_n1025), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  AND2_X1   g0831(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1032), .B1(new_n711), .B2(new_n716), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1031), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n710), .B1(new_n713), .B2(new_n714), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT87), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1034), .A2(new_n1037), .A3(new_n715), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1033), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n710), .A2(new_n697), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(new_n708), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n768), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n719), .B(KEYINPUT41), .Z(new_n1045));
  INV_X1    g0845(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n775), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1041), .A2(new_n1025), .ZN(new_n1049));
  OR2_X1    g0849(.A1(new_n1049), .A2(KEYINPUT42), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n518), .B1(new_n1022), .B2(new_n665), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n698), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(KEYINPUT42), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n987), .B(KEYINPUT107), .ZN(new_n1055));
  INV_X1    g0855(.A(KEYINPUT43), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n989), .A2(KEYINPUT43), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1054), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  AND2_X1   g0859(.A1(new_n1053), .A2(new_n1052), .ZN(new_n1060));
  NAND4_X1  g0860(.A1(new_n1060), .A2(new_n1056), .A3(new_n1055), .A4(new_n1050), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1037), .A2(new_n715), .A3(new_n1025), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1062), .B(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(KEYINPUT108), .B1(new_n1048), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n776), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT108), .ZN(new_n1068));
  NOR3_X1   g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n1064), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1015), .B1(new_n1066), .B2(new_n1069), .ZN(G387));
  OAI21_X1  g0870(.A(new_n267), .B1(new_n796), .B2(new_n825), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n841), .A2(G303), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n867), .B2(new_n1002), .C1(new_n821), .C2(new_n811), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1073), .B1(G322), .B2(new_n829), .ZN(new_n1074));
  OR2_X1    g0874(.A1(new_n1074), .A2(KEYINPUT48), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1074), .A2(KEYINPUT48), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n807), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(G294), .A2(new_n1077), .B1(new_n804), .B2(G283), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  XOR2_X1   g0879(.A(new_n1079), .B(KEYINPUT49), .Z(new_n1080));
  AOI211_X1 g0880(.A(new_n1071), .B(new_n1080), .C1(G116), .C2(new_n884), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n292), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n839), .A2(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n267), .B(new_n1001), .C1(G150), .C2(new_n797), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n805), .A2(new_n307), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(G77), .B2(new_n1077), .ZN(new_n1086));
  AOI22_X1  g0886(.A1(G68), .A2(new_n841), .B1(new_n817), .B2(G50), .ZN(new_n1087));
  NAND4_X1  g0887(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G159), .B2(new_n829), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n790), .B1(new_n1081), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n721), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n779), .A2(new_n1091), .B1(new_n501), .B2(new_n718), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n232), .A2(new_n245), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n305), .A2(new_n202), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(new_n1094), .B(KEYINPUT50), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n721), .B(new_n245), .C1(new_n344), .C2(new_n447), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n782), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1092), .B1(new_n1093), .B2(new_n1097), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n719), .B(new_n776), .C1(new_n1098), .C2(new_n991), .ZN(new_n1099));
  AND2_X1   g0899(.A1(new_n1090), .A2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n710), .A2(new_n847), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n708), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1042), .B(new_n1102), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n1100), .A2(new_n1101), .B1(new_n776), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1043), .B1(new_n759), .B2(new_n767), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1103), .A2(new_n768), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1105), .A2(new_n1106), .A3(new_n719), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1104), .A2(new_n1107), .ZN(G393));
  NAND2_X1  g0908(.A1(new_n1106), .A2(new_n1039), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1103), .A2(new_n1033), .A3(new_n768), .A4(new_n1038), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n719), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1033), .A2(new_n776), .A3(new_n1038), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n991), .B1(new_n524), .B2(new_n210), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n783), .A2(new_n242), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n777), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n829), .A2(G150), .B1(G159), .B2(new_n817), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT110), .ZN(new_n1117));
  OR2_X1    g0917(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1117), .A2(KEYINPUT51), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n267), .B(new_n870), .C1(G143), .C2(new_n797), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(G68), .A2(new_n1077), .B1(new_n804), .B2(G77), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1120), .B(new_n1121), .C1(new_n287), .C2(new_n814), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1122), .B1(G50), .B2(new_n839), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1118), .A2(new_n1119), .A3(new_n1123), .ZN(new_n1124));
  AOI22_X1  g0924(.A1(new_n829), .A2(G317), .B1(G311), .B2(new_n817), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT52), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n270), .B(new_n836), .C1(G322), .C2(new_n797), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G283), .A2(new_n1077), .B1(new_n804), .B2(G116), .ZN(new_n1128));
  AND2_X1   g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n806), .B2(new_n814), .C1(new_n808), .C2(new_n821), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1124), .B1(new_n1126), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1115), .B1(new_n1131), .B2(new_n790), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n789), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1132), .B1(new_n1133), .B2(new_n1025), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1111), .A2(new_n1112), .A3(new_n1134), .ZN(G390));
  NAND3_X1  g0935(.A1(new_n922), .A2(G330), .A3(new_n928), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n700), .B(new_n923), .C1(new_n753), .C2(new_n758), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n925), .A2(new_n927), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1136), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n855), .A2(new_n966), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n698), .B(new_n854), .C1(new_n667), .C2(new_n762), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(new_n966), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n922), .A2(G330), .A3(new_n860), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1142), .B1(new_n1143), .B2(new_n964), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n759), .A2(new_n860), .A3(new_n1138), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1139), .A2(new_n1140), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n922), .A2(G330), .A3(new_n646), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n971), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(KEYINPUT38), .B1(new_n911), .B2(new_n912), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n959), .A2(new_n1149), .A3(new_n953), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT38), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n403), .A2(KEYINPUT105), .A3(new_n388), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT105), .B1(new_n403), .B2(new_n388), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n909), .B1(new_n1154), .B2(new_n687), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1151), .B1(new_n1155), .B2(new_n939), .ZN(new_n1156));
  AOI21_X1  g0956(.A(KEYINPUT39), .B1(new_n1156), .B2(new_n913), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n1150), .A2(new_n1157), .B1(new_n961), .B2(new_n967), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1142), .A2(new_n1138), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n961), .B1(new_n1156), .B2(new_n913), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1158), .A2(new_n1145), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1136), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n1146), .A2(new_n1148), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1138), .B1(new_n759), .B2(new_n860), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n922), .A2(G330), .A3(new_n928), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1140), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1143), .A2(new_n964), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1142), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1168), .A2(new_n1145), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1158), .A2(new_n1161), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n1166), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1148), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1158), .A2(new_n1161), .A3(new_n1145), .ZN(new_n1175));
  NAND4_X1  g0975(.A1(new_n1171), .A2(new_n1173), .A3(new_n1174), .A4(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1164), .A2(new_n1176), .A3(new_n719), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n960), .A2(new_n962), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1140), .A2(new_n1138), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n961), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n1178), .A2(new_n1181), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1175), .B(new_n776), .C1(new_n1182), .C2(new_n1136), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1178), .A2(new_n787), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n777), .B1(new_n1082), .B2(new_n865), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n267), .B1(new_n797), .B2(G125), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n202), .B2(new_n800), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT111), .Z(new_n1188));
  NAND2_X1  g0988(.A1(new_n1077), .A2(G150), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT53), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n867), .A2(new_n881), .B1(new_n832), .B2(new_n805), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G137), .B2(new_n839), .ZN(new_n1192));
  XOR2_X1   g0992(.A(KEYINPUT54), .B(G143), .Z(new_n1193));
  AOI22_X1  g0993(.A1(new_n841), .A2(new_n1193), .B1(new_n1189), .B2(KEYINPUT53), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1188), .A2(new_n1190), .A3(new_n1192), .A4(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(G128), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n830), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n821), .A2(new_n501), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n867), .A2(new_n220), .B1(new_n524), .B2(new_n814), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n267), .B1(new_n796), .B2(new_n806), .C1(new_n374), .C2(new_n807), .ZN(new_n1200));
  OAI22_X1  g1000(.A1(new_n805), .A2(new_n447), .B1(new_n800), .B2(new_n344), .ZN(new_n1201));
  OR4_X1    g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .A4(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n830), .A2(new_n799), .ZN(new_n1203));
  OAI22_X1  g1003(.A1(new_n1195), .A2(new_n1197), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1185), .B1(new_n1204), .B2(new_n790), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1184), .A2(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1183), .A2(KEYINPUT112), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT112), .B1(new_n1183), .B2(new_n1206), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1177), .B1(new_n1207), .B2(new_n1208), .ZN(G378));
  NAND2_X1  g1009(.A1(new_n303), .A2(new_n333), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n295), .A2(new_n694), .ZN(new_n1211));
  OR2_X1    g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  XNOR2_X1  g1014(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1212), .A2(new_n1213), .A3(new_n1215), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n787), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n777), .B1(G50), .B2(new_n865), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n202), .B1(G33), .B2(G41), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1222), .B1(new_n267), .B2(new_n244), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n867), .A2(new_n501), .B1(new_n307), .B2(new_n814), .ZN(new_n1224));
  AOI211_X1 g1024(.A(G41), .B(new_n270), .C1(new_n797), .C2(G283), .ZN(new_n1225));
  OAI221_X1 g1025(.A(new_n1225), .B1(new_n290), .B2(new_n800), .C1(new_n447), .C2(new_n807), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1224), .B(new_n1226), .C1(G97), .C2(new_n839), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n829), .A2(G116), .B1(G68), .B2(new_n804), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT113), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n1227), .B1(new_n1230), .B2(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(KEYINPUT58), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1223), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(G33), .B(G41), .C1(new_n797), .C2(G124), .ZN(new_n1235));
  AOI22_X1  g1035(.A1(new_n841), .A2(G137), .B1(new_n1077), .B2(new_n1193), .ZN(new_n1236));
  OAI221_X1 g1036(.A(new_n1236), .B1(new_n1196), .B2(new_n867), .C1(new_n881), .C2(new_n821), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(new_n829), .A2(G125), .B1(G150), .B2(new_n804), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1238), .A2(KEYINPUT114), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(KEYINPUT114), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1237), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT59), .ZN(new_n1242));
  OAI221_X1 g1042(.A(new_n1235), .B1(new_n832), .B2(new_n800), .C1(new_n1241), .C2(new_n1242), .ZN(new_n1243));
  AND2_X1   g1043(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n1234), .B1(new_n1233), .B2(new_n1232), .C1(new_n1243), .C2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1221), .B1(new_n1245), .B2(new_n790), .ZN(new_n1246));
  AND2_X1   g1046(.A1(new_n1220), .A2(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n963), .A2(new_n968), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1138), .A2(new_n860), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n556), .A2(new_n1018), .A3(new_n592), .A4(new_n696), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n919), .A2(new_n920), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1251), .B2(new_n756), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1249), .B1(new_n1252), .B2(new_n753), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n930), .B1(new_n1156), .B2(new_n913), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n700), .B1(new_n1253), .B2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n931), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n931), .B2(new_n1255), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1248), .B1(new_n1257), .B2(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n948), .A2(G330), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT40), .B1(new_n1253), .B2(new_n915), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1219), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n931), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1262), .A2(new_n969), .A3(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1259), .A2(new_n1264), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1247), .B1(new_n1265), .B2(new_n776), .ZN(new_n1266));
  AND3_X1   g1066(.A1(new_n1262), .A2(new_n969), .A3(new_n1263), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n969), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1268));
  OAI21_X1  g1068(.A(KEYINPUT57), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1148), .B1(new_n1270), .B2(new_n1171), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n719), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1175), .B1(new_n1182), .B2(new_n1136), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1174), .B1(new_n1273), .B2(new_n1146), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT57), .B1(new_n1265), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1266), .B1(new_n1272), .B2(new_n1275), .ZN(G375));
  NAND2_X1  g1076(.A1(new_n1171), .A2(new_n776), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT115), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n964), .A2(new_n787), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n777), .B1(G68), .B2(new_n865), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n807), .A2(new_n832), .B1(new_n796), .B2(new_n1196), .ZN(new_n1281));
  OAI22_X1  g1081(.A1(new_n867), .A2(new_n877), .B1(new_n876), .B2(new_n814), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1281), .B(new_n1282), .C1(G50), .C2(new_n804), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n270), .B1(new_n800), .B2(new_n290), .ZN(new_n1284));
  XOR2_X1   g1084(.A(new_n1284), .B(KEYINPUT116), .Z(new_n1285));
  AOI21_X1  g1085(.A(new_n1285), .B1(new_n839), .B2(new_n1193), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1283), .B(new_n1286), .C1(new_n881), .C2(new_n830), .ZN(new_n1287));
  OAI22_X1  g1087(.A1(new_n867), .A2(new_n799), .B1(new_n501), .B2(new_n814), .ZN(new_n1288));
  OAI221_X1 g1088(.A(new_n267), .B1(new_n796), .B2(new_n808), .C1(new_n447), .C2(new_n800), .ZN(new_n1289));
  NOR2_X1   g1089(.A1(new_n807), .A2(new_n524), .ZN(new_n1290));
  NOR4_X1   g1090(.A1(new_n1288), .A2(new_n1085), .A3(new_n1289), .A4(new_n1290), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1291), .B1(new_n220), .B2(new_n821), .C1(new_n806), .C2(new_n830), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1287), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1280), .B1(new_n1293), .B2(new_n790), .ZN(new_n1294));
  AOI22_X1  g1094(.A1(new_n1277), .A2(new_n1278), .B1(new_n1279), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1171), .A2(KEYINPUT115), .A3(new_n776), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1171), .A2(new_n1174), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1167), .A2(new_n1148), .A3(new_n1170), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1297), .A2(new_n1046), .A3(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1295), .A2(new_n1296), .A3(new_n1299), .ZN(G381));
  XNOR2_X1  g1100(.A(G375), .B(KEYINPUT117), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1015), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1045), .B1(new_n1110), .B2(new_n768), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1065), .B(KEYINPUT108), .C1(new_n776), .C2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1068), .B1(new_n1067), .B2(new_n1064), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1303), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1177), .A2(new_n1183), .A3(new_n1206), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1107), .A2(new_n849), .A3(new_n778), .A4(new_n1104), .ZN(new_n1310));
  NOR4_X1   g1110(.A1(G381), .A2(new_n1310), .A3(G384), .A4(G390), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1302), .A2(new_n1307), .A3(new_n1309), .A4(new_n1311), .ZN(G407));
  NAND2_X1  g1112(.A1(new_n695), .A2(G213), .ZN(new_n1313));
  INV_X1    g1113(.A(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1302), .A2(new_n1309), .A3(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(G407), .A2(G213), .A3(new_n1315), .ZN(G409));
  INV_X1    g1116(.A(KEYINPUT126), .ZN(new_n1317));
  INV_X1    g1117(.A(G384), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n720), .B1(new_n1171), .B2(new_n1174), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1146), .A2(KEYINPUT60), .A3(new_n1148), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT60), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1298), .A2(new_n1321), .ZN(new_n1322));
  AND3_X1   g1122(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1278), .B1(new_n1146), .B2(new_n775), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1279), .A2(new_n1294), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1296), .A3(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1318), .B1(new_n1323), .B2(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(new_n1319), .A2(new_n1320), .A3(new_n1322), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1328), .A2(new_n1295), .A3(G384), .A4(new_n1296), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1327), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  AND4_X1   g1131(.A1(KEYINPUT118), .A2(new_n1265), .A3(new_n1274), .A4(new_n1046), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1045), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT118), .B1(new_n1333), .B2(new_n1274), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1332), .A2(new_n1334), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT119), .ZN(new_n1336));
  AOI21_X1  g1136(.A(new_n775), .B1(new_n1265), .B2(new_n1336), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1259), .A2(KEYINPUT119), .A3(new_n1264), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1247), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1339));
  AOI21_X1  g1139(.A(new_n1308), .B1(new_n1335), .B2(new_n1339), .ZN(new_n1340));
  OAI211_X1 g1140(.A(G378), .B(new_n1266), .C1(new_n1272), .C2(new_n1275), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n1341), .ZN(new_n1342));
  OAI211_X1 g1142(.A(new_n1313), .B(new_n1331), .C1(new_n1340), .C2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1343), .A2(KEYINPUT62), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1333), .A2(new_n1274), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT118), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1265), .A2(new_n1336), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1348), .A2(new_n776), .A3(new_n1338), .ZN(new_n1349));
  INV_X1    g1149(.A(new_n1247), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1333), .A2(KEYINPUT118), .A3(new_n1274), .ZN(new_n1351));
  NAND4_X1  g1151(.A1(new_n1347), .A2(new_n1349), .A3(new_n1350), .A4(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1352), .A2(new_n1309), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1341), .ZN(new_n1354));
  INV_X1    g1154(.A(KEYINPUT62), .ZN(new_n1355));
  NAND4_X1  g1155(.A1(new_n1354), .A2(new_n1355), .A3(new_n1313), .A4(new_n1331), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1344), .A2(new_n1356), .ZN(new_n1357));
  INV_X1    g1157(.A(KEYINPUT61), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT120), .ZN(new_n1359));
  INV_X1    g1159(.A(G2897), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1313), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1361), .B1(new_n1359), .B2(new_n1360), .ZN(new_n1362));
  NAND3_X1  g1162(.A1(new_n1327), .A2(new_n1329), .A3(new_n1362), .ZN(new_n1363));
  INV_X1    g1163(.A(KEYINPUT121), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1363), .A2(new_n1364), .ZN(new_n1365));
  NAND4_X1  g1165(.A1(new_n1327), .A2(KEYINPUT121), .A3(new_n1329), .A4(new_n1362), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1365), .A2(new_n1366), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1313), .A2(new_n1360), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1330), .A2(new_n1368), .ZN(new_n1369));
  NAND2_X1  g1169(.A1(new_n1367), .A2(new_n1369), .ZN(new_n1370));
  AOI21_X1  g1170(.A(new_n1314), .B1(new_n1353), .B2(new_n1341), .ZN(new_n1371));
  OAI21_X1  g1171(.A(new_n1358), .B1(new_n1370), .B2(new_n1371), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1317), .B1(new_n1357), .B2(new_n1372), .ZN(new_n1373));
  AOI22_X1  g1173(.A1(new_n1365), .A2(new_n1366), .B1(new_n1330), .B2(new_n1368), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1313), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1375));
  AOI21_X1  g1175(.A(KEYINPUT61), .B1(new_n1374), .B2(new_n1375), .ZN(new_n1376));
  NAND4_X1  g1176(.A1(new_n1376), .A2(KEYINPUT126), .A3(new_n1344), .A4(new_n1356), .ZN(new_n1377));
  NAND2_X1  g1177(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1378), .A2(new_n1015), .A3(G390), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT123), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1379), .A2(new_n1380), .ZN(new_n1381));
  INV_X1    g1181(.A(KEYINPUT124), .ZN(new_n1382));
  INV_X1    g1182(.A(G390), .ZN(new_n1383));
  NAND3_X1  g1183(.A1(G387), .A2(new_n1382), .A3(new_n1383), .ZN(new_n1384));
  OAI21_X1  g1184(.A(KEYINPUT124), .B1(new_n1307), .B2(G390), .ZN(new_n1385));
  NAND3_X1  g1185(.A1(new_n1307), .A2(KEYINPUT123), .A3(G390), .ZN(new_n1386));
  NAND4_X1  g1186(.A1(new_n1381), .A2(new_n1384), .A3(new_n1385), .A4(new_n1386), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(G393), .A2(G396), .ZN(new_n1388));
  NAND2_X1  g1188(.A1(new_n1388), .A2(new_n1310), .ZN(new_n1389));
  INV_X1    g1189(.A(new_n1389), .ZN(new_n1390));
  NAND2_X1  g1190(.A1(new_n1387), .A2(new_n1390), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT127), .ZN(new_n1392));
  INV_X1    g1192(.A(KEYINPUT125), .ZN(new_n1393));
  OAI21_X1  g1193(.A(new_n1389), .B1(new_n1307), .B2(G390), .ZN(new_n1394));
  AND3_X1   g1194(.A1(new_n1378), .A2(new_n1015), .A3(G390), .ZN(new_n1395));
  OAI21_X1  g1195(.A(new_n1393), .B1(new_n1394), .B2(new_n1395), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(G387), .A2(new_n1383), .ZN(new_n1397));
  NAND4_X1  g1197(.A1(new_n1397), .A2(KEYINPUT125), .A3(new_n1389), .A4(new_n1379), .ZN(new_n1398));
  NAND2_X1  g1198(.A1(new_n1396), .A2(new_n1398), .ZN(new_n1399));
  AND3_X1   g1199(.A1(new_n1391), .A2(new_n1392), .A3(new_n1399), .ZN(new_n1400));
  AOI21_X1  g1200(.A(new_n1392), .B1(new_n1391), .B2(new_n1399), .ZN(new_n1401));
  NOR2_X1   g1201(.A1(new_n1400), .A2(new_n1401), .ZN(new_n1402));
  NAND3_X1  g1202(.A1(new_n1373), .A2(new_n1377), .A3(new_n1402), .ZN(new_n1403));
  INV_X1    g1203(.A(KEYINPUT63), .ZN(new_n1404));
  NOR2_X1   g1204(.A1(new_n1343), .A2(new_n1404), .ZN(new_n1405));
  NOR2_X1   g1205(.A1(new_n1405), .A2(KEYINPUT61), .ZN(new_n1406));
  AOI22_X1  g1206(.A1(new_n1391), .A2(new_n1399), .B1(new_n1343), .B2(new_n1404), .ZN(new_n1407));
  AND2_X1   g1207(.A1(new_n1374), .A2(KEYINPUT122), .ZN(new_n1408));
  OAI21_X1  g1208(.A(new_n1375), .B1(new_n1374), .B2(KEYINPUT122), .ZN(new_n1409));
  OAI211_X1 g1209(.A(new_n1406), .B(new_n1407), .C1(new_n1408), .C2(new_n1409), .ZN(new_n1410));
  NAND2_X1  g1210(.A1(new_n1403), .A2(new_n1410), .ZN(G405));
  NAND2_X1  g1211(.A1(G375), .A2(new_n1309), .ZN(new_n1412));
  NAND2_X1  g1212(.A1(new_n1412), .A2(new_n1341), .ZN(new_n1413));
  XNOR2_X1  g1213(.A(new_n1413), .B(new_n1330), .ZN(new_n1414));
  NOR2_X1   g1214(.A1(new_n1402), .A2(new_n1414), .ZN(new_n1415));
  XNOR2_X1  g1215(.A(new_n1413), .B(new_n1331), .ZN(new_n1416));
  NOR3_X1   g1216(.A1(new_n1400), .A2(new_n1401), .A3(new_n1416), .ZN(new_n1417));
  NOR2_X1   g1217(.A1(new_n1415), .A2(new_n1417), .ZN(G402));
endmodule


