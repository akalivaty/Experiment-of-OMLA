

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758;

  AND2_X1 U369 ( .A1(n349), .A2(n348), .ZN(n663) );
  INV_X1 U370 ( .A(n347), .ZN(n348) );
  INV_X1 U371 ( .A(KEYINPUT77), .ZN(n351) );
  NOR2_X1 U372 ( .A1(n702), .A2(n700), .ZN(n639) );
  BUF_X1 U373 ( .A(n662), .Z(n347) );
  INV_X1 U374 ( .A(n385), .ZN(n354) );
  XNOR2_X1 U375 ( .A(n500), .B(n499), .ZN(n662) );
  XNOR2_X1 U376 ( .A(n519), .B(n352), .ZN(n534) );
  INV_X1 U377 ( .A(G478), .ZN(n352) );
  XNOR2_X1 U378 ( .A(n515), .B(n514), .ZN(n353) );
  XOR2_X1 U379 ( .A(KEYINPUT11), .B(G131), .Z(n502) );
  XOR2_X1 U380 ( .A(KEYINPUT7), .B(G134), .Z(n514) );
  INV_X1 U381 ( .A(G143), .ZN(n415) );
  XNOR2_X1 U382 ( .A(G131), .B(KEYINPUT69), .ZN(n484) );
  XNOR2_X1 U383 ( .A(G128), .B(G137), .ZN(n470) );
  NAND2_X2 U384 ( .A1(G214), .A2(n531), .ZN(n618) );
  XNOR2_X2 U385 ( .A(KEYINPUT65), .B(n678), .ZN(n390) );
  XNOR2_X2 U386 ( .A(KEYINPUT15), .B(G902), .ZN(n679) );
  XNOR2_X1 U387 ( .A(n496), .B(n433), .ZN(n683) );
  XNOR2_X1 U388 ( .A(n744), .B(n464), .ZN(n496) );
  NAND2_X1 U389 ( .A1(n346), .A2(n645), .ZN(n648) );
  XNOR2_X1 U390 ( .A(n366), .B(n643), .ZN(n346) );
  XNOR2_X2 U391 ( .A(n632), .B(KEYINPUT0), .ZN(n641) );
  XNOR2_X2 U392 ( .A(n660), .B(KEYINPUT106), .ZN(n349) );
  NAND2_X1 U393 ( .A1(n548), .A2(n652), .ZN(n368) );
  NOR2_X2 U394 ( .A1(n635), .A2(n541), .ZN(n548) );
  OR2_X2 U395 ( .A1(n716), .A2(G902), .ZN(n425) );
  XNOR2_X2 U396 ( .A(n648), .B(n647), .ZN(n756) );
  AND2_X2 U397 ( .A1(n404), .A2(KEYINPUT104), .ZN(n386) );
  NOR2_X2 U398 ( .A1(n703), .A2(KEYINPUT99), .ZN(n436) );
  NOR2_X1 U399 ( .A1(n350), .A2(n602), .ZN(n605) );
  XNOR2_X1 U400 ( .A(n592), .B(n351), .ZN(n350) );
  NAND2_X1 U401 ( .A1(n534), .A2(n599), .ZN(n533) );
  XNOR2_X2 U402 ( .A(n513), .B(n353), .ZN(n517) );
  NOR2_X2 U403 ( .A1(n377), .A2(n638), .ZN(n412) );
  XNOR2_X2 U404 ( .A(n412), .B(n411), .ZN(n703) );
  NAND2_X1 U405 ( .A1(n587), .A2(n618), .ZN(n372) );
  XNOR2_X2 U406 ( .A(n529), .B(n387), .ZN(n587) );
  OR2_X4 U407 ( .A1(n626), .A2(n354), .ZN(n632) );
  NAND2_X1 U408 ( .A1(n355), .A2(n402), .ZN(n400) );
  NAND2_X1 U409 ( .A1(n398), .A2(n386), .ZN(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT81), .B(KEYINPUT18), .ZN(n525) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(G119), .Z(n494) );
  XNOR2_X1 U412 ( .A(G122), .B(G107), .ZN(n380) );
  XNOR2_X1 U413 ( .A(G122), .B(G143), .ZN(n501) );
  XOR2_X1 U414 ( .A(KEYINPUT66), .B(G101), .Z(n381) );
  INV_X1 U415 ( .A(G119), .ZN(n374) );
  XNOR2_X2 U416 ( .A(n610), .B(n588), .ZN(n626) );
  XNOR2_X2 U417 ( .A(n359), .B(KEYINPUT80), .ZN(n526) );
  NOR2_X1 U418 ( .A1(n642), .A2(n377), .ZN(n366) );
  NAND2_X1 U419 ( .A1(n454), .A2(n389), .ZN(n453) );
  NOR2_X1 U420 ( .A1(n755), .A2(n758), .ZN(n586) );
  NOR2_X2 U421 ( .A1(n453), .A2(n452), .ZN(n690) );
  NAND2_X1 U422 ( .A1(n608), .A2(n662), .ZN(n580) );
  INV_X1 U423 ( .A(n656), .ZN(n664) );
  XNOR2_X1 U424 ( .A(n467), .B(n466), .ZN(n469) );
  XNOR2_X1 U425 ( .A(KEYINPUT16), .B(G122), .ZN(n362) );
  XNOR2_X1 U426 ( .A(KEYINPUT66), .B(G101), .ZN(n358) );
  INV_X1 U427 ( .A(G113), .ZN(n370) );
  INV_X1 U428 ( .A(KEYINPUT39), .ZN(n357) );
  INV_X1 U429 ( .A(KEYINPUT33), .ZN(n367) );
  INV_X1 U430 ( .A(G113), .ZN(n375) );
  INV_X2 U431 ( .A(G953), .ZN(n747) );
  NOR2_X1 U432 ( .A1(KEYINPUT44), .A2(n669), .ZN(n670) );
  NAND2_X1 U433 ( .A1(n664), .A2(n663), .ZN(n694) );
  AND2_X1 U434 ( .A1(n574), .A2(n700), .ZN(n576) );
  XNOR2_X1 U435 ( .A(n572), .B(n357), .ZN(n574) );
  XNOR2_X1 U436 ( .A(n368), .B(n367), .ZN(n642) );
  AND2_X1 U437 ( .A1(n656), .A2(n356), .ZN(n568) );
  XNOR2_X1 U438 ( .A(n662), .B(n432), .ZN(n652) );
  XNOR2_X1 U439 ( .A(n448), .B(n447), .ZN(n599) );
  INV_X1 U440 ( .A(n623), .ZN(n356) );
  OR2_X1 U441 ( .A1(n720), .A2(G902), .ZN(n448) );
  XNOR2_X1 U442 ( .A(n496), .B(n491), .ZN(n716) );
  XNOR2_X1 U443 ( .A(n469), .B(n468), .ZN(n512) );
  XNOR2_X1 U444 ( .A(n520), .B(n521), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n371), .B(n369), .ZN(n495) );
  XNOR2_X1 U446 ( .A(n375), .B(G104), .ZN(n520) );
  XNOR2_X1 U447 ( .A(n362), .B(n361), .ZN(n360) );
  XNOR2_X1 U448 ( .A(n374), .B(G110), .ZN(n521) );
  XNOR2_X1 U449 ( .A(n485), .B(n484), .ZN(n486) );
  INV_X1 U450 ( .A(n358), .ZN(n524) );
  XOR2_X1 U451 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n468) );
  INV_X1 U452 ( .A(KEYINPUT85), .ZN(n466) );
  NAND2_X1 U453 ( .A1(n512), .A2(G221), .ZN(n475) );
  INV_X2 U454 ( .A(KEYINPUT93), .ZN(n359) );
  XNOR2_X1 U455 ( .A(n493), .B(n492), .ZN(n363) );
  XNOR2_X2 U456 ( .A(G116), .B(KEYINPUT73), .ZN(n492) );
  XNOR2_X2 U457 ( .A(KEYINPUT72), .B(KEYINPUT3), .ZN(n493) );
  XNOR2_X1 U458 ( .A(n363), .B(n360), .ZN(n364) );
  XNOR2_X2 U459 ( .A(G107), .B(KEYINPUT75), .ZN(n361) );
  XNOR2_X1 U460 ( .A(n364), .B(n373), .ZN(n738) );
  XNOR2_X1 U461 ( .A(n527), .B(n365), .ZN(n394) );
  XNOR2_X2 U462 ( .A(n406), .B(n405), .ZN(n365) );
  XNOR2_X1 U463 ( .A(n486), .B(n365), .ZN(n744) );
  XNOR2_X1 U464 ( .A(n492), .B(n370), .ZN(n369) );
  XNOR2_X1 U465 ( .A(n494), .B(n493), .ZN(n371) );
  XNOR2_X2 U466 ( .A(n372), .B(KEYINPUT92), .ZN(n610) );
  BUF_X1 U467 ( .A(n658), .Z(n376) );
  XNOR2_X2 U468 ( .A(n632), .B(KEYINPUT0), .ZN(n377) );
  BUF_X1 U469 ( .A(n703), .Z(n378) );
  AND2_X1 U470 ( .A1(n437), .A2(n434), .ZN(n379) );
  XOR2_X2 U471 ( .A(n581), .B(KEYINPUT1), .Z(n635) );
  BUF_X1 U472 ( .A(n710), .Z(n382) );
  AND2_X1 U473 ( .A1(n422), .A2(n421), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n738), .B(n393), .ZN(n710) );
  BUF_X1 U475 ( .A(n587), .Z(n595) );
  OR2_X1 U476 ( .A1(n681), .A2(n427), .ZN(n421) );
  XNOR2_X1 U477 ( .A(n510), .B(n509), .ZN(n720) );
  NAND2_X1 U478 ( .A1(n442), .A2(KEYINPUT2), .ZN(n427) );
  XNOR2_X1 U479 ( .A(n498), .B(G472), .ZN(n499) );
  NOR2_X1 U480 ( .A1(n400), .A2(n399), .ZN(n650) );
  NAND2_X1 U481 ( .A1(n397), .A2(n396), .ZN(n399) );
  INV_X1 U482 ( .A(n746), .ZN(n442) );
  XOR2_X1 U483 ( .A(n672), .B(KEYINPUT87), .Z(n673) );
  XNOR2_X1 U484 ( .A(n495), .B(n497), .ZN(n433) );
  NAND2_X1 U485 ( .A1(n445), .A2(n443), .ZN(n746) );
  NOR2_X1 U486 ( .A1(n754), .A2(n444), .ZN(n443) );
  XNOR2_X1 U487 ( .A(n615), .B(n614), .ZN(n445) );
  INV_X1 U488 ( .A(n709), .ZN(n444) );
  INV_X1 U489 ( .A(KEYINPUT96), .ZN(n472) );
  XNOR2_X1 U490 ( .A(G140), .B(KEYINPUT10), .ZN(n446) );
  XNOR2_X1 U491 ( .A(n395), .B(n394), .ZN(n393) );
  XNOR2_X1 U492 ( .A(n430), .B(n429), .ZN(n658) );
  INV_X1 U493 ( .A(KEYINPUT22), .ZN(n429) );
  NAND2_X1 U494 ( .A1(n633), .A2(n634), .ZN(n430) );
  INV_X1 U495 ( .A(KEYINPUT6), .ZN(n432) );
  AND2_X2 U496 ( .A1(n658), .A2(n635), .ZN(n660) );
  XNOR2_X1 U497 ( .A(n683), .B(KEYINPUT62), .ZN(n684) );
  XNOR2_X1 U498 ( .A(n722), .B(n721), .ZN(n463) );
  XNOR2_X1 U499 ( .A(n720), .B(n719), .ZN(n721) );
  XOR2_X1 U500 ( .A(G104), .B(G110), .Z(n489) );
  NOR2_X1 U501 ( .A1(G952), .A2(n747), .ZN(n731) );
  XNOR2_X1 U502 ( .A(n408), .B(KEYINPUT119), .ZN(n407) );
  NAND2_X1 U503 ( .A1(n409), .A2(n383), .ZN(n408) );
  NAND2_X1 U504 ( .A1(n410), .A2(n438), .ZN(n396) );
  NAND2_X1 U505 ( .A1(n403), .A2(n438), .ZN(n402) );
  NAND2_X1 U506 ( .A1(G234), .A2(G237), .ZN(n465) );
  NOR2_X1 U507 ( .A1(G953), .A2(G237), .ZN(n504) );
  XOR2_X1 U508 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n506) );
  NAND2_X1 U509 ( .A1(n442), .A2(n441), .ZN(n680) );
  INV_X1 U510 ( .A(n679), .ZN(n441) );
  OR2_X1 U511 ( .A1(G902), .A2(G237), .ZN(n531) );
  XOR2_X1 U512 ( .A(G107), .B(G140), .Z(n488) );
  AND2_X1 U513 ( .A1(n421), .A2(n676), .ZN(n416) );
  XNOR2_X1 U514 ( .A(n562), .B(n561), .ZN(n570) );
  XNOR2_X1 U515 ( .A(n511), .B(G475), .ZN(n447) );
  INV_X1 U516 ( .A(KEYINPUT97), .ZN(n456) );
  NAND2_X1 U517 ( .A1(n458), .A2(KEYINPUT97), .ZN(n457) );
  INV_X1 U518 ( .A(n637), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n475), .B(n474), .ZN(n477) );
  XNOR2_X1 U520 ( .A(n473), .B(n472), .ZN(n474) );
  XNOR2_X1 U521 ( .A(n518), .B(n517), .ZN(n725) );
  XOR2_X1 U522 ( .A(G116), .B(KEYINPUT9), .Z(n515) );
  INV_X1 U523 ( .A(KEYINPUT31), .ZN(n411) );
  AND2_X2 U524 ( .A1(n660), .A2(n388), .ZN(n687) );
  INV_X1 U525 ( .A(KEYINPUT63), .ZN(n439) );
  INV_X1 U526 ( .A(KEYINPUT60), .ZN(n460) );
  INV_X1 U527 ( .A(n731), .ZN(n462) );
  XNOR2_X1 U528 ( .A(n716), .B(n391), .ZN(n450) );
  XNOR2_X1 U529 ( .A(n712), .B(n711), .ZN(n713) );
  INV_X1 U530 ( .A(G953), .ZN(n420) );
  XNOR2_X1 U531 ( .A(KEYINPUT118), .B(n559), .ZN(n383) );
  XOR2_X1 U532 ( .A(KEYINPUT71), .B(G469), .Z(n384) );
  OR2_X1 U533 ( .A1(n630), .A2(n629), .ZN(n385) );
  AND2_X1 U534 ( .A1(n531), .A2(G210), .ZN(n387) );
  AND2_X1 U535 ( .A1(n636), .A2(n656), .ZN(n388) );
  AND2_X1 U536 ( .A1(n459), .A2(n455), .ZN(n389) );
  INV_X1 U537 ( .A(KEYINPUT104), .ZN(n438) );
  INV_X1 U538 ( .A(KEYINPUT2), .ZN(n677) );
  XOR2_X1 U539 ( .A(n718), .B(n717), .Z(n391) );
  XOR2_X1 U540 ( .A(KEYINPUT53), .B(KEYINPUT120), .Z(n392) );
  NAND2_X1 U541 ( .A1(n710), .A2(n679), .ZN(n529) );
  XNOR2_X1 U542 ( .A(n528), .B(n523), .ZN(n395) );
  INV_X1 U543 ( .A(n687), .ZN(n397) );
  NAND2_X1 U544 ( .A1(n379), .A2(n404), .ZN(n403) );
  NOR2_X1 U545 ( .A1(n410), .A2(n426), .ZN(n398) );
  NAND2_X1 U546 ( .A1(n435), .A2(n436), .ZN(n404) );
  XNOR2_X2 U547 ( .A(KEYINPUT4), .B(KEYINPUT67), .ZN(n405) );
  XNOR2_X2 U548 ( .A(G128), .B(G143), .ZN(n406) );
  NAND2_X1 U549 ( .A1(n407), .A2(n420), .ZN(n419) );
  NAND2_X1 U550 ( .A1(n416), .A2(n424), .ZN(n409) );
  BUF_X1 U551 ( .A(n681), .Z(n735) );
  NAND2_X1 U552 ( .A1(n637), .A2(n456), .ZN(n455) );
  AND2_X1 U553 ( .A1(n690), .A2(KEYINPUT99), .ZN(n410) );
  BUF_X1 U554 ( .A(n738), .Z(n413) );
  INV_X1 U555 ( .A(n414), .ZN(n440) );
  XNOR2_X1 U556 ( .A(n524), .B(n414), .ZN(n528) );
  XNOR2_X2 U557 ( .A(G125), .B(G146), .ZN(n414) );
  AND2_X2 U558 ( .A1(n422), .A2(n421), .ZN(n723) );
  XNOR2_X1 U559 ( .A(n415), .B(G128), .ZN(n418) );
  OR2_X1 U560 ( .A1(n641), .A2(n457), .ZN(n454) );
  AND2_X1 U561 ( .A1(n377), .A2(n456), .ZN(n452) );
  XNOR2_X1 U562 ( .A(n419), .B(n392), .ZN(G75) );
  NAND2_X1 U563 ( .A1(n723), .A2(G478), .ZN(n724) );
  NAND2_X1 U564 ( .A1(n423), .A2(n390), .ZN(n422) );
  INV_X1 U565 ( .A(n682), .ZN(n423) );
  NAND2_X1 U566 ( .A1(n735), .A2(n677), .ZN(n424) );
  NOR2_X1 U567 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X2 U568 ( .A(n425), .B(n384), .ZN(n581) );
  NAND2_X1 U569 ( .A1(n437), .A2(n434), .ZN(n426) );
  XNOR2_X1 U570 ( .A(n428), .B(n439), .ZN(G57) );
  NOR2_X2 U571 ( .A1(n686), .A2(n731), .ZN(n428) );
  XNOR2_X1 U572 ( .A(n674), .B(n673), .ZN(n681) );
  XNOR2_X1 U573 ( .A(n431), .B(KEYINPUT56), .ZN(G51) );
  NOR2_X2 U574 ( .A1(n715), .A2(n731), .ZN(n431) );
  NAND2_X1 U575 ( .A1(n463), .A2(n462), .ZN(n461) );
  XNOR2_X1 U576 ( .A(n461), .B(n460), .ZN(G60) );
  INV_X1 U577 ( .A(n639), .ZN(n434) );
  INV_X1 U578 ( .A(n690), .ZN(n435) );
  NAND2_X1 U579 ( .A1(n703), .A2(KEYINPUT99), .ZN(n437) );
  XNOR2_X1 U580 ( .A(n440), .B(n446), .ZN(n743) );
  NOR2_X1 U581 ( .A1(n449), .A2(n731), .ZN(G54) );
  XNOR2_X1 U582 ( .A(n451), .B(n450), .ZN(n449) );
  NAND2_X1 U583 ( .A1(n417), .A2(G469), .ZN(n451) );
  INV_X1 U584 ( .A(n347), .ZN(n459) );
  NOR2_X2 U585 ( .A1(n726), .A2(n731), .ZN(n727) );
  XNOR2_X1 U586 ( .A(n714), .B(n713), .ZN(n715) );
  XOR2_X1 U587 ( .A(n381), .B(G146), .Z(n464) );
  INV_X1 U588 ( .A(KEYINPUT76), .ZN(n604) );
  XNOR2_X1 U589 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U590 ( .A(n522), .B(KEYINPUT17), .ZN(n523) );
  INV_X1 U591 ( .A(KEYINPUT30), .ZN(n561) );
  INV_X1 U592 ( .A(KEYINPUT98), .ZN(n498) );
  XNOR2_X1 U593 ( .A(n479), .B(KEYINPUT25), .ZN(n480) );
  XNOR2_X1 U594 ( .A(n481), .B(n480), .ZN(n656) );
  XNOR2_X1 U595 ( .A(n685), .B(n684), .ZN(n686) );
  XNOR2_X1 U596 ( .A(n465), .B(KEYINPUT14), .ZN(n564) );
  NAND2_X1 U597 ( .A1(n564), .A2(G952), .ZN(n563) );
  NAND2_X1 U598 ( .A1(G234), .A2(n747), .ZN(n467) );
  XOR2_X1 U599 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n471) );
  XNOR2_X1 U600 ( .A(n471), .B(n470), .ZN(n473) );
  XNOR2_X1 U601 ( .A(n521), .B(n743), .ZN(n476) );
  XNOR2_X1 U602 ( .A(n477), .B(n476), .ZN(n729) );
  NOR2_X1 U603 ( .A1(G902), .A2(n729), .ZN(n481) );
  NAND2_X1 U604 ( .A1(n679), .A2(G234), .ZN(n478) );
  XNOR2_X1 U605 ( .A(n478), .B(KEYINPUT20), .ZN(n482) );
  NAND2_X1 U606 ( .A1(G217), .A2(n482), .ZN(n479) );
  NAND2_X1 U607 ( .A1(G221), .A2(n482), .ZN(n483) );
  XNOR2_X1 U608 ( .A(KEYINPUT21), .B(n483), .ZN(n623) );
  INV_X1 U609 ( .A(n568), .ZN(n541) );
  XOR2_X2 U610 ( .A(G134), .B(G137), .Z(n485) );
  NAND2_X1 U611 ( .A1(G227), .A2(n747), .ZN(n487) );
  XNOR2_X1 U612 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U613 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U614 ( .A1(n504), .A2(G210), .ZN(n497) );
  NOR2_X1 U615 ( .A1(G902), .A2(n683), .ZN(n500) );
  XNOR2_X1 U616 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U617 ( .A(n743), .B(n503), .ZN(n510) );
  XNOR2_X1 U618 ( .A(n520), .B(KEYINPUT12), .ZN(n508) );
  NAND2_X1 U619 ( .A1(n504), .A2(G214), .ZN(n505) );
  XNOR2_X1 U620 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U621 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U622 ( .A(KEYINPUT13), .B(KEYINPUT102), .ZN(n511) );
  NAND2_X1 U623 ( .A1(G217), .A2(n512), .ZN(n518) );
  XOR2_X1 U624 ( .A(n418), .B(n380), .Z(n513) );
  NOR2_X1 U625 ( .A1(G902), .A2(n725), .ZN(n519) );
  INV_X1 U626 ( .A(n534), .ZN(n598) );
  NAND2_X1 U627 ( .A1(n599), .A2(n598), .ZN(n624) );
  NAND2_X1 U628 ( .A1(G224), .A2(n747), .ZN(n522) );
  XNOR2_X1 U629 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U630 ( .A(KEYINPUT38), .B(KEYINPUT79), .Z(n530) );
  XOR2_X1 U631 ( .A(n595), .B(n530), .Z(n560) );
  NOR2_X1 U632 ( .A1(n560), .A2(n618), .ZN(n532) );
  NOR2_X1 U633 ( .A1(n624), .A2(n532), .ZN(n536) );
  XNOR2_X2 U634 ( .A(n533), .B(KEYINPUT103), .ZN(n702) );
  NOR2_X1 U635 ( .A1(n534), .A2(n599), .ZN(n700) );
  NAND2_X1 U636 ( .A1(n560), .A2(n618), .ZN(n539) );
  NOR2_X1 U637 ( .A1(n639), .A2(n539), .ZN(n535) );
  NOR2_X1 U638 ( .A1(n536), .A2(n535), .ZN(n537) );
  XOR2_X1 U639 ( .A(KEYINPUT117), .B(n537), .Z(n538) );
  NOR2_X1 U640 ( .A1(n642), .A2(n538), .ZN(n554) );
  NOR2_X1 U641 ( .A1(n624), .A2(n539), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n540), .B(KEYINPUT41), .ZN(n583) );
  XNOR2_X1 U643 ( .A(KEYINPUT116), .B(KEYINPUT51), .ZN(n551) );
  NAND2_X1 U644 ( .A1(n635), .A2(n541), .ZN(n542) );
  XNOR2_X1 U645 ( .A(n542), .B(KEYINPUT50), .ZN(n547) );
  XOR2_X1 U646 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n544) );
  AND2_X1 U647 ( .A1(n623), .A2(n664), .ZN(n543) );
  XOR2_X1 U648 ( .A(n544), .B(n543), .Z(n545) );
  NOR2_X1 U649 ( .A1(n347), .A2(n545), .ZN(n546) );
  NAND2_X1 U650 ( .A1(n547), .A2(n546), .ZN(n549) );
  NAND2_X1 U651 ( .A1(n548), .A2(n347), .ZN(n638) );
  NAND2_X1 U652 ( .A1(n549), .A2(n638), .ZN(n550) );
  XNOR2_X1 U653 ( .A(n551), .B(n550), .ZN(n552) );
  NOR2_X1 U654 ( .A1(n583), .A2(n552), .ZN(n553) );
  NOR2_X1 U655 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U656 ( .A(n555), .B(KEYINPUT52), .ZN(n556) );
  NOR2_X1 U657 ( .A1(n563), .A2(n556), .ZN(n558) );
  NOR2_X1 U658 ( .A1(n642), .A2(n583), .ZN(n557) );
  NOR2_X1 U659 ( .A1(n558), .A2(n557), .ZN(n559) );
  INV_X1 U660 ( .A(n560), .ZN(n571) );
  NAND2_X1 U661 ( .A1(n618), .A2(n662), .ZN(n562) );
  NOR2_X1 U662 ( .A1(G953), .A2(n563), .ZN(n630) );
  NAND2_X1 U663 ( .A1(n564), .A2(G902), .ZN(n565) );
  XOR2_X1 U664 ( .A(KEYINPUT94), .B(n565), .Z(n627) );
  NAND2_X1 U665 ( .A1(n627), .A2(G953), .ZN(n566) );
  NOR2_X1 U666 ( .A1(G900), .A2(n566), .ZN(n567) );
  NOR2_X1 U667 ( .A1(n630), .A2(n567), .ZN(n577) );
  NAND2_X1 U668 ( .A1(n581), .A2(n568), .ZN(n637) );
  NOR2_X1 U669 ( .A1(n577), .A2(n637), .ZN(n569) );
  NAND2_X1 U670 ( .A1(n570), .A2(n569), .ZN(n596) );
  NOR2_X1 U671 ( .A1(n571), .A2(n596), .ZN(n572) );
  NAND2_X1 U672 ( .A1(n574), .A2(n702), .ZN(n573) );
  XNOR2_X1 U673 ( .A(KEYINPUT111), .B(n573), .ZN(n754) );
  XNOR2_X1 U674 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n575) );
  XNOR2_X1 U675 ( .A(n576), .B(n575), .ZN(n755) );
  NOR2_X1 U676 ( .A1(n577), .A2(n623), .ZN(n578) );
  AND2_X1 U677 ( .A1(n664), .A2(n578), .ZN(n608) );
  XNOR2_X1 U678 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n579) );
  XNOR2_X1 U679 ( .A(n580), .B(n579), .ZN(n582) );
  NAND2_X1 U680 ( .A1(n582), .A2(n581), .ZN(n589) );
  NOR2_X1 U681 ( .A1(n583), .A2(n589), .ZN(n584) );
  XNOR2_X1 U682 ( .A(KEYINPUT42), .B(n584), .ZN(n758) );
  XNOR2_X1 U683 ( .A(KEYINPUT46), .B(KEYINPUT89), .ZN(n585) );
  XNOR2_X1 U684 ( .A(n586), .B(n585), .ZN(n607) );
  INV_X1 U685 ( .A(KEYINPUT19), .ZN(n588) );
  NOR2_X1 U686 ( .A1(n626), .A2(n589), .ZN(n698) );
  INV_X1 U687 ( .A(n698), .ZN(n593) );
  NOR2_X1 U688 ( .A1(KEYINPUT47), .A2(n639), .ZN(n590) );
  XOR2_X1 U689 ( .A(KEYINPUT78), .B(n590), .Z(n591) );
  NOR2_X1 U690 ( .A1(n593), .A2(n591), .ZN(n592) );
  OR2_X1 U691 ( .A1(n639), .A2(n593), .ZN(n594) );
  NAND2_X1 U692 ( .A1(n594), .A2(KEYINPUT47), .ZN(n601) );
  INV_X1 U693 ( .A(n595), .ZN(n621) );
  NOR2_X1 U694 ( .A1(n621), .A2(n596), .ZN(n597) );
  XNOR2_X1 U695 ( .A(KEYINPUT108), .B(n597), .ZN(n600) );
  NOR2_X1 U696 ( .A1(n599), .A2(n598), .ZN(n640) );
  NAND2_X1 U697 ( .A1(n600), .A2(n640), .ZN(n697) );
  NAND2_X1 U698 ( .A1(n601), .A2(n697), .ZN(n602) );
  NOR2_X1 U699 ( .A1(n607), .A2(n606), .ZN(n613) );
  AND2_X1 U700 ( .A1(n608), .A2(n700), .ZN(n609) );
  NAND2_X1 U701 ( .A1(n609), .A2(n652), .ZN(n616) );
  NOR2_X1 U702 ( .A1(n610), .A2(n616), .ZN(n611) );
  XNOR2_X1 U703 ( .A(n611), .B(KEYINPUT36), .ZN(n612) );
  INV_X1 U704 ( .A(n635), .ZN(n653) );
  NAND2_X1 U705 ( .A1(n612), .A2(n653), .ZN(n707) );
  NAND2_X1 U706 ( .A1(n613), .A2(n707), .ZN(n615) );
  XOR2_X1 U707 ( .A(KEYINPUT48), .B(KEYINPUT70), .Z(n614) );
  NOR2_X1 U708 ( .A1(n653), .A2(n616), .ZN(n617) );
  NAND2_X1 U709 ( .A1(n618), .A2(n617), .ZN(n620) );
  XOR2_X1 U710 ( .A(KEYINPUT43), .B(KEYINPUT107), .Z(n619) );
  XNOR2_X1 U711 ( .A(n620), .B(n619), .ZN(n622) );
  NAND2_X1 U712 ( .A1(n622), .A2(n621), .ZN(n709) );
  INV_X1 U713 ( .A(n652), .ZN(n636) );
  OR2_X1 U714 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U715 ( .A(n625), .B(KEYINPUT105), .ZN(n634) );
  NOR2_X1 U716 ( .A1(G898), .A2(n747), .ZN(n740) );
  NAND2_X1 U717 ( .A1(n740), .A2(n627), .ZN(n628) );
  XNOR2_X1 U718 ( .A(KEYINPUT95), .B(n628), .ZN(n629) );
  INV_X1 U719 ( .A(n641), .ZN(n633) );
  XOR2_X1 U720 ( .A(n640), .B(KEYINPUT83), .Z(n645) );
  XNOR2_X1 U721 ( .A(KEYINPUT74), .B(KEYINPUT34), .ZN(n643) );
  XNOR2_X1 U722 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n646) );
  XNOR2_X1 U723 ( .A(n646), .B(KEYINPUT82), .ZN(n647) );
  NAND2_X1 U724 ( .A1(n756), .A2(KEYINPUT44), .ZN(n649) );
  NAND2_X1 U725 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U726 ( .A(n651), .B(KEYINPUT91), .ZN(n666) );
  XOR2_X1 U727 ( .A(KEYINPUT84), .B(n652), .Z(n654) );
  NAND2_X1 U728 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U729 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U730 ( .A1(n376), .A2(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(n659), .B(KEYINPUT32), .ZN(n757) );
  NAND2_X1 U732 ( .A1(n757), .A2(n694), .ZN(n668) );
  NAND2_X1 U733 ( .A1(KEYINPUT44), .A2(n668), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n666), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(n667), .B(KEYINPUT90), .ZN(n671) );
  OR2_X1 U736 ( .A1(n668), .A2(n756), .ZN(n669) );
  NOR2_X1 U737 ( .A1(n671), .A2(n670), .ZN(n674) );
  XNOR2_X1 U738 ( .A(KEYINPUT45), .B(KEYINPUT64), .ZN(n672) );
  NAND2_X1 U739 ( .A1(n746), .A2(n677), .ZN(n675) );
  XNOR2_X1 U740 ( .A(n675), .B(KEYINPUT86), .ZN(n676) );
  NOR2_X1 U741 ( .A1(n677), .A2(n679), .ZN(n678) );
  NAND2_X1 U742 ( .A1(n723), .A2(G472), .ZN(n685) );
  XOR2_X1 U743 ( .A(n687), .B(G101), .Z(n688) );
  XNOR2_X1 U744 ( .A(KEYINPUT112), .B(n688), .ZN(G3) );
  NAND2_X1 U745 ( .A1(n690), .A2(n700), .ZN(n689) );
  XNOR2_X1 U746 ( .A(n689), .B(G104), .ZN(G6) );
  XOR2_X1 U747 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n692) );
  NAND2_X1 U748 ( .A1(n690), .A2(n702), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U750 ( .A(G107), .B(n693), .ZN(G9) );
  XNOR2_X1 U751 ( .A(G110), .B(n694), .ZN(G12) );
  XOR2_X1 U752 ( .A(G128), .B(KEYINPUT29), .Z(n696) );
  NAND2_X1 U753 ( .A1(n698), .A2(n702), .ZN(n695) );
  XNOR2_X1 U754 ( .A(n696), .B(n695), .ZN(G30) );
  XNOR2_X1 U755 ( .A(G143), .B(n697), .ZN(G45) );
  NAND2_X1 U756 ( .A1(n698), .A2(n700), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n699), .B(G146), .ZN(G48) );
  NAND2_X1 U758 ( .A1(n378), .A2(n700), .ZN(n701) );
  XNOR2_X1 U759 ( .A(n701), .B(G113), .ZN(G15) );
  NAND2_X1 U760 ( .A1(n378), .A2(n702), .ZN(n704) );
  XNOR2_X1 U761 ( .A(n704), .B(G116), .ZN(G18) );
  XOR2_X1 U762 ( .A(KEYINPUT113), .B(KEYINPUT114), .Z(n706) );
  XNOR2_X1 U763 ( .A(G125), .B(KEYINPUT37), .ZN(n705) );
  XNOR2_X1 U764 ( .A(n706), .B(n705), .ZN(n708) );
  XOR2_X1 U765 ( .A(n708), .B(n707), .Z(G27) );
  XNOR2_X1 U766 ( .A(G140), .B(n709), .ZN(G42) );
  NAND2_X1 U767 ( .A1(n723), .A2(G210), .ZN(n714) );
  INV_X1 U768 ( .A(n382), .ZN(n712) );
  XOR2_X1 U769 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n711) );
  XOR2_X1 U770 ( .A(KEYINPUT122), .B(KEYINPUT121), .Z(n718) );
  XNOR2_X1 U771 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n717) );
  NAND2_X1 U772 ( .A1(n417), .A2(G475), .ZN(n722) );
  XOR2_X1 U773 ( .A(KEYINPUT123), .B(KEYINPUT59), .Z(n719) );
  XNOR2_X1 U774 ( .A(n724), .B(n725), .ZN(n726) );
  XNOR2_X1 U775 ( .A(n727), .B(KEYINPUT124), .ZN(G63) );
  NAND2_X1 U776 ( .A1(G217), .A2(n417), .ZN(n728) );
  XNOR2_X1 U777 ( .A(n729), .B(n728), .ZN(n730) );
  NOR2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G66) );
  NAND2_X1 U779 ( .A1(G953), .A2(G224), .ZN(n732) );
  XNOR2_X1 U780 ( .A(KEYINPUT61), .B(n732), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n733), .A2(G898), .ZN(n734) );
  XNOR2_X1 U782 ( .A(n734), .B(KEYINPUT125), .ZN(n737) );
  NOR2_X1 U783 ( .A1(G953), .A2(n735), .ZN(n736) );
  NOR2_X1 U784 ( .A1(n737), .A2(n736), .ZN(n742) );
  XNOR2_X1 U785 ( .A(n413), .B(G101), .ZN(n739) );
  NOR2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U787 ( .A(n742), .B(n741), .Z(G69) );
  XOR2_X1 U788 ( .A(n744), .B(n743), .Z(n745) );
  XNOR2_X1 U789 ( .A(KEYINPUT126), .B(n745), .ZN(n749) );
  XNOR2_X1 U790 ( .A(n749), .B(n746), .ZN(n748) );
  NAND2_X1 U791 ( .A1(n748), .A2(n747), .ZN(n753) );
  XNOR2_X1 U792 ( .A(G227), .B(n749), .ZN(n750) );
  NAND2_X1 U793 ( .A1(n750), .A2(G900), .ZN(n751) );
  NAND2_X1 U794 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U795 ( .A1(n753), .A2(n752), .ZN(G72) );
  XOR2_X1 U796 ( .A(G134), .B(n754), .Z(G36) );
  XOR2_X1 U797 ( .A(G131), .B(n755), .Z(G33) );
  XOR2_X1 U798 ( .A(n756), .B(G122), .Z(G24) );
  XNOR2_X1 U799 ( .A(G119), .B(n757), .ZN(G21) );
  XOR2_X1 U800 ( .A(G137), .B(n758), .Z(G39) );
endmodule

