

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744;

  NOR2_X1 U366 ( .A1(n528), .A2(n526), .ZN(n642) );
  XNOR2_X1 U367 ( .A(G113), .B(KEYINPUT68), .ZN(n449) );
  NOR2_X2 U368 ( .A1(n554), .A2(n553), .ZN(n599) );
  XNOR2_X2 U369 ( .A(n468), .B(n467), .ZN(n718) );
  XNOR2_X2 U370 ( .A(n409), .B(KEYINPUT4), .ZN(n475) );
  XNOR2_X2 U371 ( .A(n530), .B(KEYINPUT1), .ZN(n653) );
  AND2_X2 U372 ( .A1(n607), .A2(n606), .ZN(n712) );
  XNOR2_X1 U373 ( .A(n399), .B(n350), .ZN(n742) );
  NAND2_X1 U374 ( .A1(n395), .A2(n392), .ZN(n686) );
  XNOR2_X1 U375 ( .A(n516), .B(n517), .ZN(n368) );
  OR2_X1 U376 ( .A1(n534), .A2(n532), .ZN(n516) );
  XNOR2_X1 U377 ( .A(n472), .B(G134), .ZN(n488) );
  XNOR2_X1 U378 ( .A(G119), .B(G116), .ZN(n450) );
  XNOR2_X1 U379 ( .A(n484), .B(KEYINPUT39), .ZN(n548) );
  XNOR2_X2 U380 ( .A(n464), .B(n463), .ZN(n525) );
  NAND2_X1 U381 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X1 U382 ( .A1(n362), .A2(n360), .ZN(n359) );
  NAND2_X1 U383 ( .A1(n389), .A2(n387), .ZN(n542) );
  AND2_X1 U384 ( .A1(n594), .A2(n388), .ZN(n387) );
  INV_X1 U385 ( .A(n523), .ZN(n388) );
  NAND2_X1 U386 ( .A1(n525), .A2(n670), .ZN(n484) );
  NAND2_X1 U387 ( .A1(n356), .A2(n354), .ZN(n365) );
  NAND2_X1 U388 ( .A1(n355), .A2(n348), .ZN(n354) );
  AND2_X1 U389 ( .A1(n364), .A2(n357), .ZN(n356) );
  NAND2_X1 U390 ( .A1(n371), .A2(n370), .ZN(n369) );
  AND2_X1 U391 ( .A1(n742), .A2(n519), .ZN(n373) );
  NOR2_X1 U392 ( .A1(G953), .A2(G237), .ZN(n446) );
  INV_X1 U393 ( .A(KEYINPUT48), .ZN(n375) );
  INV_X1 U394 ( .A(KEYINPUT41), .ZN(n398) );
  XNOR2_X1 U395 ( .A(n488), .B(n384), .ZN(n730) );
  XNOR2_X1 U396 ( .A(n475), .B(n385), .ZN(n384) );
  XNOR2_X1 U397 ( .A(n386), .B(G131), .ZN(n385) );
  INV_X1 U398 ( .A(G137), .ZN(n386) );
  XNOR2_X1 U399 ( .A(G143), .B(G131), .ZN(n502) );
  XOR2_X1 U400 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n498) );
  XNOR2_X1 U401 ( .A(G104), .B(G122), .ZN(n495) );
  XOR2_X1 U402 ( .A(KEYINPUT11), .B(KEYINPUT98), .Z(n496) );
  NAND2_X1 U403 ( .A1(n403), .A2(n597), .ZN(n598) );
  XNOR2_X1 U404 ( .A(n405), .B(n404), .ZN(n403) );
  NOR2_X1 U405 ( .A1(n672), .A2(n398), .ZN(n397) );
  INV_X1 U406 ( .A(KEYINPUT38), .ZN(n390) );
  INV_X1 U407 ( .A(KEYINPUT23), .ZN(n421) );
  XNOR2_X1 U408 ( .A(n557), .B(n556), .ZN(n687) );
  XNOR2_X1 U409 ( .A(KEYINPUT87), .B(KEYINPUT33), .ZN(n556) );
  NOR2_X1 U410 ( .A1(n592), .A2(n687), .ZN(n400) );
  INV_X1 U411 ( .A(KEYINPUT76), .ZN(n463) );
  INV_X1 U412 ( .A(n532), .ZN(n663) );
  NOR2_X1 U413 ( .A1(G902), .A2(n713), .ZN(n433) );
  INV_X1 U414 ( .A(KEYINPUT47), .ZN(n360) );
  INV_X1 U415 ( .A(KEYINPUT81), .ZN(n362) );
  INV_X1 U416 ( .A(n542), .ZN(n355) );
  NAND2_X1 U417 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U418 ( .A(KEYINPUT44), .ZN(n404) );
  NAND2_X1 U419 ( .A1(G234), .A2(G237), .ZN(n438) );
  INV_X1 U420 ( .A(G237), .ZN(n458) );
  XNOR2_X1 U421 ( .A(n376), .B(n375), .ZN(n551) );
  XNOR2_X1 U422 ( .A(n730), .B(n383), .ZN(n455) );
  INV_X1 U423 ( .A(G146), .ZN(n383) );
  NOR2_X1 U424 ( .A1(n591), .A2(n513), .ZN(n380) );
  XNOR2_X1 U425 ( .A(n431), .B(n430), .ZN(n434) );
  XNOR2_X1 U426 ( .A(KEYINPUT20), .B(KEYINPUT94), .ZN(n430) );
  BUF_X1 U427 ( .A(n604), .Z(n734) );
  XOR2_X1 U428 ( .A(KEYINPUT9), .B(G122), .Z(n486) );
  XNOR2_X1 U429 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U430 ( .A(n503), .B(n502), .ZN(n504) );
  INV_X1 U431 ( .A(KEYINPUT66), .ZN(n409) );
  NAND2_X1 U432 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U433 ( .A(n367), .B(n366), .ZN(n524) );
  INV_X1 U434 ( .A(KEYINPUT109), .ZN(n366) );
  NAND2_X1 U435 ( .A1(n368), .A2(n518), .ZN(n367) );
  INV_X1 U436 ( .A(n353), .ZN(n657) );
  NAND2_X1 U437 ( .A1(n382), .A2(n381), .ZN(n591) );
  INV_X1 U438 ( .A(n530), .ZN(n382) );
  INV_X1 U439 ( .A(n555), .ZN(n381) );
  INV_X1 U440 ( .A(KEYINPUT0), .ZN(n401) );
  AND2_X1 U441 ( .A1(n563), .A2(n562), .ZN(n402) );
  XNOR2_X1 U442 ( .A(n663), .B(n533), .ZN(n584) );
  XNOR2_X1 U443 ( .A(KEYINPUT16), .B(G122), .ZN(n465) );
  XNOR2_X1 U444 ( .A(n428), .B(n427), .ZN(n713) );
  XNOR2_X1 U445 ( .A(n729), .B(n420), .ZN(n428) );
  XNOR2_X1 U446 ( .A(G128), .B(G137), .ZN(n425) );
  INV_X1 U447 ( .A(n696), .ZN(n606) );
  AND2_X1 U448 ( .A1(n611), .A2(G953), .ZN(n717) );
  INV_X1 U449 ( .A(G953), .ZN(n736) );
  AND2_X1 U450 ( .A1(n548), .A2(n642), .ZN(n511) );
  XNOR2_X1 U451 ( .A(n540), .B(n539), .ZN(n541) );
  NOR2_X1 U452 ( .A1(n543), .A2(n391), .ZN(n540) );
  NOR2_X1 U453 ( .A1(n565), .A2(n391), .ZN(n529) );
  NOR2_X1 U454 ( .A1(n593), .A2(n592), .ZN(n344) );
  XOR2_X1 U455 ( .A(n482), .B(n481), .Z(n345) );
  XNOR2_X1 U456 ( .A(G146), .B(G125), .ZN(n469) );
  XNOR2_X1 U457 ( .A(n432), .B(KEYINPUT25), .ZN(n346) );
  OR2_X1 U458 ( .A1(KEYINPUT47), .A2(n542), .ZN(n347) );
  AND2_X1 U459 ( .A1(n639), .A2(n362), .ZN(n348) );
  NOR2_X1 U460 ( .A1(n578), .A2(n353), .ZN(n349) );
  XNOR2_X1 U461 ( .A(KEYINPUT110), .B(KEYINPUT42), .ZN(n350) );
  AND2_X1 U462 ( .A1(KEYINPUT81), .A2(KEYINPUT47), .ZN(n351) );
  XNOR2_X2 U463 ( .A(n352), .B(n469), .ZN(n729) );
  XNOR2_X1 U464 ( .A(n408), .B(G140), .ZN(n352) );
  NAND2_X1 U465 ( .A1(n353), .A2(n569), .ZN(n555) );
  XNOR2_X2 U466 ( .A(n433), .B(n346), .ZN(n353) );
  NAND2_X1 U467 ( .A1(n653), .A2(n353), .ZN(n583) );
  NAND2_X1 U468 ( .A1(n361), .A2(n358), .ZN(n357) );
  NAND2_X1 U469 ( .A1(n639), .A2(n359), .ZN(n358) );
  INV_X1 U470 ( .A(n639), .ZN(n363) );
  NAND2_X1 U471 ( .A1(n542), .A2(n351), .ZN(n364) );
  NAND2_X1 U472 ( .A1(n347), .A2(n365), .ZN(n378) );
  INV_X1 U473 ( .A(n524), .ZN(n389) );
  NAND2_X1 U474 ( .A1(n372), .A2(n369), .ZN(n379) );
  NOR2_X1 U475 ( .A1(n742), .A2(n519), .ZN(n370) );
  INV_X1 U476 ( .A(n743), .ZN(n371) );
  NOR2_X1 U477 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X1 U478 ( .A1(n743), .A2(n519), .ZN(n374) );
  NAND2_X1 U479 ( .A1(n379), .A2(n377), .ZN(n376) );
  NOR2_X1 U480 ( .A1(n647), .A2(n378), .ZN(n377) );
  NAND2_X1 U481 ( .A1(n462), .A2(n380), .ZN(n464) );
  XNOR2_X2 U482 ( .A(G143), .B(G128), .ZN(n472) );
  NOR2_X1 U483 ( .A1(n524), .A2(n523), .ZN(n640) );
  NAND2_X1 U484 ( .A1(n546), .A2(n669), .ZN(n522) );
  XNOR2_X2 U485 ( .A(n546), .B(n390), .ZN(n670) );
  INV_X1 U486 ( .A(n546), .ZN(n391) );
  XNOR2_X2 U487 ( .A(n483), .B(n345), .ZN(n546) );
  AND2_X1 U488 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U489 ( .A1(n672), .A2(n398), .ZN(n393) );
  NAND2_X1 U490 ( .A1(n673), .A2(n398), .ZN(n394) );
  INV_X1 U491 ( .A(n673), .ZN(n396) );
  NOR2_X2 U492 ( .A1(n524), .A2(n686), .ZN(n399) );
  XNOR2_X1 U493 ( .A(n400), .B(n564), .ZN(n567) );
  XNOR2_X2 U494 ( .A(n402), .B(n401), .ZN(n592) );
  NOR2_X1 U495 ( .A1(n741), .A2(n622), .ZN(n406) );
  INV_X1 U496 ( .A(n625), .ZN(n407) );
  XNOR2_X2 U497 ( .A(n582), .B(n581), .ZN(n625) );
  OR2_X2 U498 ( .A1(n617), .A2(n601), .ZN(n483) );
  XNOR2_X2 U499 ( .A(n417), .B(G469), .ZN(n530) );
  XNOR2_X1 U500 ( .A(KEYINPUT67), .B(KEYINPUT10), .ZN(n408) );
  INV_X1 U501 ( .A(KEYINPUT74), .ZN(n552) );
  XNOR2_X1 U502 ( .A(n604), .B(n552), .ZN(n554) );
  INV_X1 U503 ( .A(n649), .ZN(n549) );
  BUF_X1 U504 ( .A(n555), .Z(n652) );
  NOR2_X1 U505 ( .A1(n650), .A2(n549), .ZN(n550) );
  XNOR2_X1 U506 ( .A(n422), .B(n421), .ZN(n424) );
  XNOR2_X1 U507 ( .A(n436), .B(n435), .ZN(n658) );
  XNOR2_X1 U508 ( .A(n424), .B(n423), .ZN(n426) );
  INV_X1 U509 ( .A(KEYINPUT36), .ZN(n539) );
  XNOR2_X1 U510 ( .A(G107), .B(G104), .ZN(n411) );
  INV_X1 U511 ( .A(G110), .ZN(n410) );
  XNOR2_X1 U512 ( .A(n411), .B(n410), .ZN(n413) );
  XNOR2_X1 U513 ( .A(G101), .B(KEYINPUT73), .ZN(n412) );
  XNOR2_X1 U514 ( .A(n413), .B(n412), .ZN(n467) );
  NAND2_X1 U515 ( .A1(G227), .A2(n736), .ZN(n414) );
  XNOR2_X1 U516 ( .A(n414), .B(G140), .ZN(n415) );
  XNOR2_X1 U517 ( .A(n467), .B(n415), .ZN(n416) );
  XNOR2_X1 U518 ( .A(n455), .B(n416), .ZN(n703) );
  NOR2_X1 U519 ( .A1(G902), .A2(n703), .ZN(n417) );
  XOR2_X1 U520 ( .A(KEYINPUT82), .B(KEYINPUT8), .Z(n419) );
  NAND2_X1 U521 ( .A1(G234), .A2(n736), .ZN(n418) );
  XNOR2_X1 U522 ( .A(n419), .B(n418), .ZN(n489) );
  NAND2_X1 U523 ( .A1(n489), .A2(G221), .ZN(n420) );
  XNOR2_X1 U524 ( .A(G119), .B(G110), .ZN(n422) );
  XOR2_X1 U525 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U526 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U527 ( .A(G902), .B(KEYINPUT90), .ZN(n429) );
  XNOR2_X1 U528 ( .A(n429), .B(KEYINPUT15), .ZN(n553) );
  NAND2_X1 U529 ( .A1(G234), .A2(n553), .ZN(n431) );
  NAND2_X1 U530 ( .A1(G217), .A2(n434), .ZN(n432) );
  XOR2_X1 U531 ( .A(KEYINPUT95), .B(KEYINPUT21), .Z(n436) );
  NAND2_X1 U532 ( .A1(G221), .A2(n434), .ZN(n435) );
  INV_X1 U533 ( .A(KEYINPUT96), .ZN(n437) );
  XNOR2_X1 U534 ( .A(n658), .B(n437), .ZN(n569) );
  XOR2_X1 U535 ( .A(KEYINPUT14), .B(KEYINPUT91), .Z(n439) );
  XNOR2_X1 U536 ( .A(n439), .B(n438), .ZN(n440) );
  NAND2_X1 U537 ( .A1(G952), .A2(n440), .ZN(n684) );
  NOR2_X1 U538 ( .A1(G953), .A2(n684), .ZN(n560) );
  NAND2_X1 U539 ( .A1(G902), .A2(n440), .ZN(n558) );
  OR2_X1 U540 ( .A1(n736), .A2(n558), .ZN(n441) );
  NOR2_X1 U541 ( .A1(G900), .A2(n441), .ZN(n442) );
  NOR2_X1 U542 ( .A1(n560), .A2(n442), .ZN(n443) );
  XNOR2_X1 U543 ( .A(KEYINPUT80), .B(n443), .ZN(n513) );
  XOR2_X1 U544 ( .A(KEYINPUT30), .B(KEYINPUT106), .Z(n461) );
  XOR2_X1 U545 ( .A(KEYINPUT97), .B(KEYINPUT5), .Z(n445) );
  XNOR2_X1 U546 ( .A(G101), .B(KEYINPUT72), .ZN(n444) );
  XNOR2_X1 U547 ( .A(n445), .B(n444), .ZN(n448) );
  XOR2_X1 U548 ( .A(KEYINPUT75), .B(n446), .Z(n501) );
  NAND2_X1 U549 ( .A1(n501), .A2(G210), .ZN(n447) );
  XNOR2_X1 U550 ( .A(n448), .B(n447), .ZN(n453) );
  XNOR2_X1 U551 ( .A(n450), .B(n449), .ZN(n452) );
  XNOR2_X1 U552 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n452), .B(n451), .ZN(n466) );
  XNOR2_X1 U554 ( .A(n453), .B(n466), .ZN(n454) );
  XNOR2_X1 U555 ( .A(n455), .B(n454), .ZN(n608) );
  NOR2_X1 U556 ( .A1(n608), .A2(G902), .ZN(n457) );
  INV_X1 U557 ( .A(G472), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n457), .B(n456), .ZN(n515) );
  INV_X1 U559 ( .A(G902), .ZN(n459) );
  NAND2_X1 U560 ( .A1(n459), .A2(n458), .ZN(n480) );
  NAND2_X1 U561 ( .A1(n480), .A2(G214), .ZN(n669) );
  NAND2_X1 U562 ( .A1(n515), .A2(n669), .ZN(n460) );
  XNOR2_X1 U563 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U564 ( .A(n466), .B(n465), .ZN(n468) );
  NAND2_X1 U565 ( .A1(n736), .A2(G224), .ZN(n470) );
  XNOR2_X1 U566 ( .A(n469), .B(n470), .ZN(n471) );
  XNOR2_X1 U567 ( .A(n472), .B(n471), .ZN(n478) );
  XOR2_X1 U568 ( .A(KEYINPUT88), .B(KEYINPUT17), .Z(n474) );
  XNOR2_X1 U569 ( .A(KEYINPUT77), .B(KEYINPUT18), .ZN(n473) );
  XNOR2_X1 U570 ( .A(n474), .B(n473), .ZN(n476) );
  XNOR2_X1 U571 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U573 ( .A(n718), .B(n479), .ZN(n617) );
  INV_X1 U574 ( .A(n553), .ZN(n601) );
  NAND2_X1 U575 ( .A1(n480), .A2(G210), .ZN(n482) );
  INV_X1 U576 ( .A(KEYINPUT79), .ZN(n481) );
  XNOR2_X1 U577 ( .A(G116), .B(G107), .ZN(n485) );
  XNOR2_X1 U578 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U579 ( .A(n488), .B(n487), .Z(n491) );
  NAND2_X1 U580 ( .A1(G217), .A2(n489), .ZN(n490) );
  XNOR2_X1 U581 ( .A(n491), .B(n490), .ZN(n493) );
  XOR2_X1 U582 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n492) );
  XNOR2_X1 U583 ( .A(n493), .B(n492), .ZN(n709) );
  NOR2_X1 U584 ( .A1(G902), .A2(n709), .ZN(n494) );
  XOR2_X1 U585 ( .A(G478), .B(n494), .Z(n528) );
  XNOR2_X1 U586 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U587 ( .A(G113), .B(KEYINPUT12), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U589 ( .A(n500), .B(n499), .Z(n505) );
  NAND2_X1 U590 ( .A1(G214), .A2(n501), .ZN(n503) );
  XNOR2_X1 U591 ( .A(n506), .B(n729), .ZN(n626) );
  NOR2_X1 U592 ( .A1(n626), .A2(G902), .ZN(n510) );
  XOR2_X1 U593 ( .A(KEYINPUT13), .B(KEYINPUT101), .Z(n508) );
  XNOR2_X1 U594 ( .A(KEYINPUT102), .B(G475), .ZN(n507) );
  XNOR2_X1 U595 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U596 ( .A(n510), .B(n509), .Z(n526) );
  XNOR2_X1 U597 ( .A(n511), .B(KEYINPUT40), .ZN(n743) );
  INV_X1 U598 ( .A(n528), .ZN(n512) );
  AND2_X1 U599 ( .A1(n512), .A2(n526), .ZN(n570) );
  INV_X1 U600 ( .A(n570), .ZN(n672) );
  NAND2_X1 U601 ( .A1(n670), .A2(n669), .ZN(n673) );
  XNOR2_X1 U602 ( .A(KEYINPUT107), .B(n530), .ZN(n518) );
  XOR2_X1 U603 ( .A(KEYINPUT108), .B(KEYINPUT28), .Z(n517) );
  NOR2_X1 U604 ( .A1(n658), .A2(n513), .ZN(n514) );
  NAND2_X1 U605 ( .A1(n657), .A2(n514), .ZN(n534) );
  INV_X1 U606 ( .A(n515), .ZN(n532) );
  XNOR2_X1 U607 ( .A(KEYINPUT46), .B(KEYINPUT85), .ZN(n519) );
  INV_X1 U608 ( .A(KEYINPUT65), .ZN(n520) );
  XNOR2_X1 U609 ( .A(n520), .B(KEYINPUT19), .ZN(n521) );
  XNOR2_X1 U610 ( .A(n522), .B(n521), .ZN(n563) );
  INV_X1 U611 ( .A(n563), .ZN(n523) );
  AND2_X1 U612 ( .A1(n528), .A2(n526), .ZN(n644) );
  NOR2_X1 U613 ( .A1(n644), .A2(n642), .ZN(n674) );
  INV_X1 U614 ( .A(n674), .ZN(n594) );
  INV_X1 U615 ( .A(n526), .ZN(n527) );
  NAND2_X1 U616 ( .A1(n528), .A2(n527), .ZN(n565) );
  NAND2_X1 U617 ( .A1(n525), .A2(n529), .ZN(n639) );
  INV_X1 U618 ( .A(KEYINPUT89), .ZN(n531) );
  XNOR2_X1 U619 ( .A(n653), .B(n531), .ZN(n578) );
  INV_X1 U620 ( .A(KEYINPUT6), .ZN(n533) );
  INV_X1 U621 ( .A(n642), .ZN(n535) );
  NOR2_X1 U622 ( .A1(n535), .A2(n534), .ZN(n536) );
  NAND2_X1 U623 ( .A1(n584), .A2(n536), .ZN(n537) );
  XNOR2_X1 U624 ( .A(n537), .B(KEYINPUT105), .ZN(n538) );
  NAND2_X1 U625 ( .A1(n538), .A2(n669), .ZN(n543) );
  NOR2_X1 U626 ( .A1(n578), .A2(n541), .ZN(n647) );
  INV_X1 U627 ( .A(n653), .ZN(n544) );
  NOR2_X1 U628 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U629 ( .A(n545), .B(KEYINPUT43), .ZN(n547) );
  NOR2_X1 U630 ( .A1(n547), .A2(n546), .ZN(n650) );
  NAND2_X1 U631 ( .A1(n548), .A2(n644), .ZN(n649) );
  AND2_X2 U632 ( .A1(n551), .A2(n550), .ZN(n604) );
  NOR2_X1 U633 ( .A1(n653), .A2(n652), .ZN(n588) );
  NAND2_X1 U634 ( .A1(n588), .A2(n584), .ZN(n557) );
  INV_X1 U635 ( .A(G898), .ZN(n724) );
  NAND2_X1 U636 ( .A1(G953), .A2(n724), .ZN(n719) );
  NOR2_X1 U637 ( .A1(n558), .A2(n719), .ZN(n559) );
  OR2_X1 U638 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U639 ( .A(n561), .B(KEYINPUT92), .ZN(n562) );
  XNOR2_X1 U640 ( .A(KEYINPUT70), .B(KEYINPUT34), .ZN(n564) );
  INV_X1 U641 ( .A(n565), .ZN(n566) );
  NAND2_X1 U642 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U643 ( .A(n568), .B(KEYINPUT35), .ZN(n741) );
  NAND2_X1 U644 ( .A1(n570), .A2(n569), .ZN(n571) );
  OR2_X1 U645 ( .A1(n592), .A2(n571), .ZN(n574) );
  XNOR2_X1 U646 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n572) );
  XNOR2_X1 U647 ( .A(n572), .B(KEYINPUT64), .ZN(n573) );
  XNOR2_X1 U648 ( .A(n574), .B(n573), .ZN(n586) );
  NAND2_X1 U649 ( .A1(n653), .A2(n657), .ZN(n575) );
  NOR2_X1 U650 ( .A1(n575), .A2(n663), .ZN(n576) );
  AND2_X1 U651 ( .A1(n586), .A2(n576), .ZN(n622) );
  INV_X1 U652 ( .A(KEYINPUT78), .ZN(n577) );
  XNOR2_X1 U653 ( .A(n584), .B(n577), .ZN(n579) );
  AND2_X1 U654 ( .A1(n579), .A2(n349), .ZN(n580) );
  NAND2_X1 U655 ( .A1(n580), .A2(n586), .ZN(n582) );
  INV_X1 U656 ( .A(KEYINPUT32), .ZN(n581) );
  NOR2_X1 U657 ( .A1(n584), .A2(n583), .ZN(n585) );
  NAND2_X1 U658 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U659 ( .A(n587), .B(KEYINPUT104), .ZN(n624) );
  AND2_X1 U660 ( .A1(n663), .A2(n588), .ZN(n666) );
  INV_X1 U661 ( .A(n666), .ZN(n589) );
  OR2_X1 U662 ( .A1(n589), .A2(n592), .ZN(n590) );
  XNOR2_X1 U663 ( .A(n590), .B(KEYINPUT31), .ZN(n645) );
  OR2_X1 U664 ( .A1(n663), .A2(n591), .ZN(n593) );
  OR2_X1 U665 ( .A1(n645), .A2(n344), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n596) );
  AND2_X1 U667 ( .A1(n624), .A2(n596), .ZN(n597) );
  XNOR2_X2 U668 ( .A(n598), .B(KEYINPUT45), .ZN(n690) );
  NAND2_X1 U669 ( .A1(n599), .A2(n690), .ZN(n600) );
  XNOR2_X1 U670 ( .A(n600), .B(KEYINPUT84), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n601), .A2(KEYINPUT2), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n607) );
  AND2_X1 U673 ( .A1(n734), .A2(KEYINPUT2), .ZN(n605) );
  AND2_X1 U674 ( .A1(n690), .A2(n605), .ZN(n696) );
  NAND2_X1 U675 ( .A1(n712), .A2(G472), .ZN(n610) );
  XNOR2_X1 U676 ( .A(n608), .B(KEYINPUT62), .ZN(n609) );
  XNOR2_X1 U677 ( .A(n610), .B(n609), .ZN(n612) );
  INV_X1 U678 ( .A(G952), .ZN(n611) );
  NOR2_X2 U679 ( .A1(n612), .A2(n717), .ZN(n614) );
  INV_X1 U680 ( .A(KEYINPUT63), .ZN(n613) );
  XNOR2_X1 U681 ( .A(n614), .B(n613), .ZN(G57) );
  NAND2_X1 U682 ( .A1(n712), .A2(G210), .ZN(n619) );
  XOR2_X1 U683 ( .A(KEYINPUT86), .B(KEYINPUT55), .Z(n615) );
  XNOR2_X1 U684 ( .A(n615), .B(KEYINPUT54), .ZN(n616) );
  XNOR2_X1 U685 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U686 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U687 ( .A1(n620), .A2(n717), .ZN(n621) );
  XNOR2_X1 U688 ( .A(n621), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U689 ( .A(G110), .B(KEYINPUT112), .ZN(n623) );
  XOR2_X1 U690 ( .A(n623), .B(n622), .Z(G12) );
  XNOR2_X1 U691 ( .A(n624), .B(G101), .ZN(G3) );
  XOR2_X1 U692 ( .A(G119), .B(n625), .Z(G21) );
  NAND2_X1 U693 ( .A1(n712), .A2(G475), .ZN(n628) );
  XOR2_X1 U694 ( .A(KEYINPUT59), .B(n626), .Z(n627) );
  XNOR2_X1 U695 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X2 U696 ( .A1(n629), .A2(n717), .ZN(n631) );
  XOR2_X1 U697 ( .A(KEYINPUT123), .B(KEYINPUT60), .Z(n630) );
  XNOR2_X1 U698 ( .A(n631), .B(n630), .ZN(G60) );
  NAND2_X1 U699 ( .A1(n344), .A2(n642), .ZN(n632) );
  XNOR2_X1 U700 ( .A(n632), .B(G104), .ZN(G6) );
  XOR2_X1 U701 ( .A(KEYINPUT27), .B(KEYINPUT111), .Z(n634) );
  NAND2_X1 U702 ( .A1(n344), .A2(n644), .ZN(n633) );
  XNOR2_X1 U703 ( .A(n634), .B(n633), .ZN(n636) );
  XOR2_X1 U704 ( .A(G107), .B(KEYINPUT26), .Z(n635) );
  XNOR2_X1 U705 ( .A(n636), .B(n635), .ZN(G9) );
  XOR2_X1 U706 ( .A(G128), .B(KEYINPUT29), .Z(n638) );
  NAND2_X1 U707 ( .A1(n640), .A2(n644), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(G30) );
  XNOR2_X1 U709 ( .A(G143), .B(n639), .ZN(G45) );
  NAND2_X1 U710 ( .A1(n640), .A2(n642), .ZN(n641) );
  XNOR2_X1 U711 ( .A(n641), .B(G146), .ZN(G48) );
  NAND2_X1 U712 ( .A1(n642), .A2(n645), .ZN(n643) );
  XNOR2_X1 U713 ( .A(G113), .B(n643), .ZN(G15) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n646), .B(G116), .ZN(G18) );
  XNOR2_X1 U716 ( .A(G125), .B(n647), .ZN(n648) );
  XNOR2_X1 U717 ( .A(n648), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U718 ( .A(G134), .B(n649), .ZN(G36) );
  XNOR2_X1 U719 ( .A(n650), .B(G140), .ZN(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT113), .ZN(G42) );
  XOR2_X1 U721 ( .A(KEYINPUT121), .B(KEYINPUT53), .Z(n701) );
  XOR2_X1 U722 ( .A(KEYINPUT115), .B(KEYINPUT50), .Z(n655) );
  NAND2_X1 U723 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(n656) );
  XNOR2_X1 U725 ( .A(KEYINPUT114), .B(n656), .ZN(n661) );
  NAND2_X1 U726 ( .A1(n658), .A2(n657), .ZN(n659) );
  XOR2_X1 U727 ( .A(KEYINPUT49), .B(n659), .Z(n660) );
  NAND2_X1 U728 ( .A1(n661), .A2(n660), .ZN(n662) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U730 ( .A(n664), .B(KEYINPUT116), .ZN(n665) );
  NOR2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n667) );
  XOR2_X1 U732 ( .A(KEYINPUT51), .B(n667), .Z(n668) );
  NOR2_X1 U733 ( .A1(n686), .A2(n668), .ZN(n681) );
  NOR2_X1 U734 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n672), .A2(n671), .ZN(n677) );
  NOR2_X1 U736 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U737 ( .A(KEYINPUT117), .B(n675), .Z(n676) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U739 ( .A(n678), .B(KEYINPUT118), .ZN(n679) );
  NOR2_X1 U740 ( .A1(n687), .A2(n679), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U742 ( .A(n682), .B(KEYINPUT52), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n684), .A2(n683), .ZN(n685) );
  XNOR2_X1 U744 ( .A(n685), .B(KEYINPUT119), .ZN(n689) );
  OR2_X1 U745 ( .A1(n687), .A2(n686), .ZN(n688) );
  NAND2_X1 U746 ( .A1(n689), .A2(n688), .ZN(n698) );
  INV_X1 U747 ( .A(n690), .ZN(n721) );
  INV_X1 U748 ( .A(KEYINPUT2), .ZN(n691) );
  NAND2_X1 U749 ( .A1(n721), .A2(n691), .ZN(n694) );
  NOR2_X1 U750 ( .A1(KEYINPUT2), .A2(n734), .ZN(n692) );
  XNOR2_X1 U751 ( .A(n692), .B(KEYINPUT83), .ZN(n693) );
  NAND2_X1 U752 ( .A1(n694), .A2(n693), .ZN(n695) );
  NOR2_X1 U753 ( .A1(n696), .A2(n695), .ZN(n697) );
  NOR2_X1 U754 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U755 ( .A1(n699), .A2(n736), .ZN(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  XOR2_X1 U757 ( .A(KEYINPUT120), .B(n702), .Z(G75) );
  XNOR2_X1 U758 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n705) );
  XNOR2_X1 U759 ( .A(n703), .B(KEYINPUT57), .ZN(n704) );
  XNOR2_X1 U760 ( .A(n705), .B(n704), .ZN(n707) );
  NAND2_X1 U761 ( .A1(n712), .A2(G469), .ZN(n706) );
  XOR2_X1 U762 ( .A(n707), .B(n706), .Z(n708) );
  NOR2_X1 U763 ( .A1(n717), .A2(n708), .ZN(G54) );
  NAND2_X1 U764 ( .A1(n712), .A2(G478), .ZN(n710) );
  XNOR2_X1 U765 ( .A(n710), .B(n709), .ZN(n711) );
  NOR2_X1 U766 ( .A1(n717), .A2(n711), .ZN(G63) );
  NAND2_X1 U767 ( .A1(n712), .A2(G217), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n713), .B(KEYINPUT124), .ZN(n714) );
  XNOR2_X1 U769 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U770 ( .A1(n717), .A2(n716), .ZN(G66) );
  XOR2_X1 U771 ( .A(KEYINPUT125), .B(n718), .Z(n720) );
  NAND2_X1 U772 ( .A1(n720), .A2(n719), .ZN(n728) );
  NOR2_X1 U773 ( .A1(n721), .A2(G953), .ZN(n726) );
  NAND2_X1 U774 ( .A1(G953), .A2(G224), .ZN(n722) );
  XOR2_X1 U775 ( .A(KEYINPUT61), .B(n722), .Z(n723) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U777 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U778 ( .A(n728), .B(n727), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n730), .B(n729), .ZN(n735) );
  XNOR2_X1 U780 ( .A(G227), .B(n735), .ZN(n731) );
  NAND2_X1 U781 ( .A1(n731), .A2(G900), .ZN(n732) );
  XOR2_X1 U782 ( .A(KEYINPUT126), .B(n732), .Z(n733) );
  NAND2_X1 U783 ( .A1(G953), .A2(n733), .ZN(n739) );
  XNOR2_X1 U784 ( .A(n735), .B(n734), .ZN(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U786 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U787 ( .A(n740), .B(KEYINPUT127), .ZN(G72) );
  XOR2_X1 U788 ( .A(G122), .B(n741), .Z(G24) );
  XOR2_X1 U789 ( .A(n742), .B(G137), .Z(G39) );
  BUF_X1 U790 ( .A(n743), .Z(n744) );
  XOR2_X1 U791 ( .A(G131), .B(n744), .Z(G33) );
endmodule

