//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:22 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n547, new_n548, new_n549,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n563, new_n564, new_n565, new_n566, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n617, new_n618, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203, new_n1204;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT65), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(G567), .B2(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(KEYINPUT67), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n464));
  OR2_X1    g039(.A1(new_n463), .A2(KEYINPUT68), .ZN(new_n465));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n464), .B(new_n465), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(G101), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n468), .A2(G2105), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n471), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g053(.A(new_n478), .B(KEYINPUT69), .Z(G160));
  NOR2_X1   g054(.A1(new_n468), .A2(new_n472), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(G136), .B2(new_n476), .ZN(G162));
  INV_X1    g060(.A(KEYINPUT72), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  AND2_X1   g062(.A1(G126), .A2(G2105), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(KEYINPUT70), .B(new_n488), .C1(new_n466), .C2(new_n467), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  AND2_X1   g069(.A1(KEYINPUT71), .A2(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n494), .B(new_n495), .C1(new_n467), .C2(new_n466), .ZN(new_n496));
  OR2_X1    g071(.A1(G102), .A2(G2105), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n497), .B(G2104), .C1(G114), .C2(new_n472), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n472), .A2(G138), .ZN(new_n499));
  OR2_X1    g074(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n500));
  NAND2_X1  g075(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g077(.A(KEYINPUT71), .B(KEYINPUT4), .ZN(new_n503));
  OAI211_X1 g078(.A(new_n496), .B(new_n498), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n486), .B1(new_n492), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n496), .A2(new_n498), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n488), .B1(new_n466), .B2(new_n467), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT70), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(new_n490), .ZN(new_n511));
  INV_X1    g086(.A(new_n503), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n512), .B1(new_n468), .B2(new_n499), .ZN(new_n513));
  NAND4_X1  g088(.A1(new_n507), .A2(new_n511), .A3(KEYINPUT72), .A4(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n505), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(G164));
  INV_X1    g091(.A(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(G651), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n519), .B2(KEYINPUT73), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT73), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .A3(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n517), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G50), .ZN(new_n524));
  INV_X1    g099(.A(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n520), .A2(new_n522), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT5), .A2(G543), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT5), .A2(G543), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n524), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n519), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n531), .A2(new_n533), .ZN(G303));
  INV_X1    g109(.A(G303), .ZN(G166));
  XNOR2_X1  g110(.A(KEYINPUT74), .B(G51), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n523), .A2(new_n536), .ZN(new_n537));
  AND2_X1   g112(.A1(G63), .A2(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT7), .ZN(new_n540));
  INV_X1    g115(.A(KEYINPUT7), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n541), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n529), .A2(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(G89), .ZN(new_n544));
  OAI211_X1 g119(.A(new_n537), .B(new_n543), .C1(new_n544), .C2(new_n530), .ZN(G286));
  INV_X1    g120(.A(G286), .ZN(G168));
  NAND2_X1  g121(.A1(new_n523), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n526), .A2(G90), .A3(new_n529), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n529), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n549));
  OAI211_X1 g124(.A(new_n547), .B(new_n548), .C1(new_n549), .C2(new_n519), .ZN(G301));
  INV_X1    g125(.A(G301), .ZN(G171));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  AND2_X1   g127(.A1(new_n527), .A2(new_n528), .ZN(new_n553));
  INV_X1    g128(.A(G56), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  AND2_X1   g130(.A1(new_n526), .A2(new_n529), .ZN(new_n556));
  AOI22_X1  g131(.A1(G651), .A2(new_n555), .B1(new_n556), .B2(G81), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n523), .A2(G43), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G860), .ZN(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g137(.A(KEYINPUT75), .B(KEYINPUT8), .Z(new_n563));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n563), .B(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT76), .ZN(G188));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n568), .B1(new_n523), .B2(G53), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT9), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n556), .A2(G91), .ZN(new_n572));
  NAND2_X1  g147(.A1(G78), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(G65), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n553), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G651), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n569), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n523), .A2(new_n568), .A3(G53), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n578), .A2(KEYINPUT9), .A3(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n556), .A2(G87), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n523), .A2(G49), .ZN(new_n583));
  OAI21_X1  g158(.A(G651), .B1(new_n529), .B2(G74), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(G288));
  AOI22_X1  g160(.A1(new_n556), .A2(G86), .B1(G48), .B2(new_n523), .ZN(new_n586));
  INV_X1    g161(.A(G61), .ZN(new_n587));
  AOI21_X1  g162(.A(new_n587), .B1(new_n527), .B2(new_n528), .ZN(new_n588));
  AND2_X1   g163(.A1(G73), .A2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(G651), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(KEYINPUT78), .ZN(new_n591));
  INV_X1    g166(.A(KEYINPUT78), .ZN(new_n592));
  OAI211_X1 g167(.A(new_n592), .B(G651), .C1(new_n588), .C2(new_n589), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n586), .A2(new_n591), .A3(new_n593), .ZN(G305));
  NAND2_X1  g169(.A1(new_n523), .A2(G47), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n529), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  OAI221_X1 g172(.A(new_n595), .B1(new_n530), .B2(new_n596), .C1(new_n519), .C2(new_n597), .ZN(G290));
  NAND2_X1  g173(.A1(G301), .A2(G868), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT79), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n526), .A2(G92), .A3(new_n529), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(new_n603));
  INV_X1    g178(.A(G66), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n604), .B1(new_n527), .B2(new_n528), .ZN(new_n605));
  AND2_X1   g180(.A1(G79), .A2(G543), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI21_X1  g184(.A(KEYINPUT80), .B1(new_n605), .B2(new_n606), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n609), .A2(G651), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n523), .A2(G54), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n603), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n600), .B1(G868), .B2(new_n614), .ZN(G284));
  OAI21_X1  g190(.A(new_n600), .B1(G868), .B2(new_n614), .ZN(G321));
  NAND2_X1  g191(.A1(G286), .A2(G868), .ZN(new_n617));
  AND3_X1   g192(.A1(new_n578), .A2(KEYINPUT9), .A3(new_n579), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n571), .A2(new_n572), .A3(new_n576), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n617), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n614), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n626), .B1(G868), .B2(new_n560), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NOR2_X1   g203(.A1(new_n468), .A2(new_n473), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT12), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  AOI22_X1  g209(.A1(G123), .A2(new_n480), .B1(new_n476), .B2(G135), .ZN(new_n635));
  NOR3_X1   g210(.A1(new_n472), .A2(KEYINPUT81), .A3(G111), .ZN(new_n636));
  OAI21_X1  g211(.A(KEYINPUT81), .B1(new_n472), .B2(G111), .ZN(new_n637));
  OAI211_X1 g212(.A(new_n637), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(G2096), .Z(new_n640));
  NAND3_X1  g215(.A1(new_n633), .A2(new_n634), .A3(new_n640), .ZN(G156));
  XNOR2_X1  g216(.A(G2427), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2430), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT15), .B(G2435), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g224(.A(G1341), .B(G1348), .Z(new_n650));
  XNOR2_X1  g225(.A(new_n649), .B(new_n650), .ZN(new_n651));
  XOR2_X1   g226(.A(G2451), .B(G2454), .Z(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT82), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n651), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(G14), .A3(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT83), .ZN(new_n658));
  INV_X1    g233(.A(KEYINPUT83), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n655), .A2(new_n659), .A3(G14), .A4(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n665), .A2(KEYINPUT18), .ZN(new_n666));
  XNOR2_X1  g241(.A(G2072), .B(G2078), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2096), .B(G2100), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT84), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n668), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n665), .A2(KEYINPUT17), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n663), .A2(new_n664), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n672), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n671), .B(new_n675), .Z(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT85), .B(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1956), .B(G2474), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1961), .B(G1966), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n679), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT20), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n679), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  OR2_X1    g262(.A1(new_n679), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n685), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(G1981), .B(G1986), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n692), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n691), .B(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(new_n694), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(G229));
  INV_X1    g276(.A(G16), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G22), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G166), .B2(new_n702), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(KEYINPUT90), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(KEYINPUT90), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(G1971), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n702), .A2(G23), .ZN(new_n710));
  INV_X1    g285(.A(G288), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n702), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT33), .B(G1976), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT89), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n712), .B(new_n714), .ZN(new_n715));
  MUX2_X1   g290(.A(G6), .B(G305), .S(G16), .Z(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT32), .B(G1981), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT88), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n716), .B(new_n718), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n705), .A2(G1971), .A3(new_n706), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n709), .A2(new_n715), .A3(new_n719), .A4(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G25), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n726));
  INV_X1    g301(.A(G107), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n726), .B1(new_n727), .B2(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT86), .Z(new_n729));
  AOI22_X1  g304(.A1(G119), .A2(new_n480), .B1(new_n476), .B2(G131), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n725), .B1(new_n731), .B2(new_n724), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XOR2_X1   g308(.A(new_n732), .B(new_n733), .Z(new_n734));
  NOR2_X1   g309(.A1(G16), .A2(G24), .ZN(new_n735));
  XOR2_X1   g310(.A(G290), .B(KEYINPUT87), .Z(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(G16), .ZN(new_n737));
  INV_X1    g312(.A(G1986), .ZN(new_n738));
  OR2_X1    g313(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n738), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n721), .B2(KEYINPUT34), .ZN(new_n742));
  OAI21_X1  g317(.A(KEYINPUT36), .B1(new_n723), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n721), .A2(KEYINPUT34), .ZN(new_n744));
  INV_X1    g319(.A(KEYINPUT36), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n744), .A2(new_n745), .A3(new_n722), .A4(new_n741), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n724), .A2(G32), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT98), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  NAND2_X1  g327(.A1(new_n476), .A2(G141), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n480), .A2(G129), .ZN(new_n754));
  INV_X1    g329(.A(G105), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n753), .B(new_n754), .C1(new_n755), .C2(new_n473), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n749), .B1(new_n757), .B2(new_n724), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT27), .B(G1996), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(KEYINPUT99), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n702), .A2(G21), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G168), .B2(new_n702), .ZN(new_n763));
  INV_X1    g338(.A(G1961), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n702), .A2(G5), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G301), .B2(G16), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n763), .A2(G1966), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n763), .A2(G1966), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT101), .Z(new_n770));
  NAND2_X1  g345(.A1(G160), .A2(G29), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(KEYINPUT24), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G34), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n773), .A2(new_n724), .ZN(new_n774));
  AOI21_X1  g349(.A(G2084), .B1(new_n771), .B2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT100), .ZN(new_n777));
  INV_X1    g352(.A(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n777), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n781), .B1(new_n639), .B2(new_n724), .C1(new_n766), .C2(new_n764), .ZN(new_n782));
  NOR4_X1   g357(.A1(new_n768), .A2(new_n770), .A3(new_n775), .A4(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n724), .A2(G27), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(KEYINPUT102), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G164), .B2(new_n724), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(G2078), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n771), .A2(G2084), .A3(new_n774), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT97), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n788), .A2(new_n789), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n787), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n783), .A2(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT103), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT92), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT25), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n476), .A2(G139), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT93), .ZN(new_n800));
  NAND2_X1  g375(.A1(G115), .A2(G2104), .ZN(new_n801));
  INV_X1    g376(.A(G127), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n801), .B1(new_n468), .B2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT94), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n472), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n804), .B2(new_n803), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n800), .A2(KEYINPUT95), .A3(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  AOI21_X1  g383(.A(KEYINPUT95), .B1(new_n800), .B2(new_n806), .ZN(new_n809));
  OAI21_X1  g384(.A(G29), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(G2072), .ZN(new_n811));
  INV_X1    g386(.A(G33), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n810), .B(new_n811), .C1(G29), .C2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n809), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n724), .B1(new_n814), .B2(new_n807), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n812), .A2(G29), .ZN(new_n816));
  OAI21_X1  g391(.A(G2072), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n793), .A2(new_n794), .A3(new_n813), .A4(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n817), .A2(new_n813), .A3(new_n783), .A4(new_n792), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT103), .ZN(new_n820));
  NOR2_X1   g395(.A1(G29), .A2(G35), .ZN(new_n821));
  AOI21_X1  g396(.A(new_n821), .B1(G162), .B2(G29), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT29), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2090), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n724), .A2(G26), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT28), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n476), .A2(G140), .ZN(new_n827));
  XOR2_X1   g402(.A(new_n827), .B(KEYINPUT91), .Z(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n829));
  INV_X1    g404(.A(G116), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(G2105), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n480), .B2(G128), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n826), .B1(new_n833), .B2(G29), .ZN(new_n834));
  INV_X1    g409(.A(G2067), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n834), .B(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n702), .A2(G19), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n560), .B2(new_n702), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(G1341), .ZN(new_n839));
  NOR3_X1   g414(.A1(new_n824), .A2(new_n836), .A3(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n702), .A2(G20), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT23), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n620), .B2(new_n702), .ZN(new_n843));
  INV_X1    g418(.A(G1956), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n702), .A2(G4), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(new_n614), .B2(new_n702), .ZN(new_n847));
  XOR2_X1   g422(.A(new_n847), .B(G1348), .Z(new_n848));
  AND3_X1   g423(.A1(new_n840), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n818), .A2(new_n820), .A3(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(KEYINPUT104), .B1(new_n748), .B2(new_n850), .ZN(new_n851));
  AND2_X1   g426(.A1(new_n818), .A2(new_n849), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT104), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n852), .A2(new_n747), .A3(new_n853), .A4(new_n820), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(G311));
  NAND3_X1  g430(.A1(new_n852), .A2(new_n747), .A3(new_n820), .ZN(G150));
  NAND2_X1  g431(.A1(new_n614), .A2(G559), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT38), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n523), .A2(G55), .ZN(new_n859));
  INV_X1    g434(.A(G93), .ZN(new_n860));
  AOI22_X1  g435(.A1(new_n529), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n861));
  OAI221_X1 g436(.A(new_n859), .B1(new_n530), .B2(new_n860), .C1(new_n861), .C2(new_n519), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n559), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n519), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n530), .A2(new_n860), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n866), .A2(new_n557), .A3(new_n558), .A4(new_n859), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n858), .B(new_n869), .ZN(new_n870));
  AND2_X1   g445(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n870), .A2(KEYINPUT39), .ZN(new_n872));
  NOR3_X1   g447(.A1(new_n871), .A2(new_n872), .A3(G860), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n862), .A2(G860), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  OR2_X1    g450(.A1(new_n873), .A2(new_n875), .ZN(G145));
  INV_X1    g451(.A(KEYINPUT40), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n731), .B(new_n630), .Z(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n757), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n880), .B1(new_n808), .B2(new_n809), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n814), .A2(new_n807), .A3(new_n757), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n504), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(new_n511), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n833), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n480), .A2(G130), .ZN(new_n888));
  NOR2_X1   g463(.A1(new_n472), .A2(G118), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT106), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n476), .A2(new_n891), .A3(G142), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n891), .B1(new_n476), .B2(G142), .ZN(new_n893));
  OAI221_X1 g468(.A(new_n888), .B1(new_n889), .B2(new_n890), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n887), .B(new_n894), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n881), .A2(new_n882), .A3(new_n879), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n884), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n895), .ZN(new_n898));
  INV_X1    g473(.A(new_n896), .ZN(new_n899));
  OAI21_X1  g474(.A(new_n898), .B1(new_n899), .B2(new_n883), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n639), .B(KEYINPUT105), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n901), .B(G160), .Z(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(G162), .ZN(new_n903));
  INV_X1    g478(.A(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n897), .A2(new_n900), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(G37), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n897), .B2(new_n900), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n877), .B1(new_n907), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n908), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n910), .A2(KEYINPUT40), .A3(new_n906), .A4(new_n905), .ZN(new_n911));
  AND2_X1   g486(.A1(new_n909), .A2(new_n911), .ZN(G395));
  XNOR2_X1  g487(.A(new_n869), .B(new_n625), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n613), .A2(new_n914), .A3(new_n577), .A4(new_n580), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n519), .B1(new_n607), .B2(new_n608), .ZN(new_n916));
  AOI22_X1  g491(.A1(new_n916), .A2(new_n610), .B1(G54), .B2(new_n523), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n603), .B(new_n917), .C1(new_n618), .C2(new_n619), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n914), .B1(new_n620), .B2(new_n613), .ZN(new_n920));
  NOR2_X1   g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g496(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(KEYINPUT41), .B1(new_n919), .B2(new_n920), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT107), .B1(new_n614), .B2(G299), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT41), .ZN(new_n925));
  NAND4_X1  g500(.A1(new_n924), .A2(new_n925), .A3(new_n918), .A4(new_n915), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n913), .A2(new_n923), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n922), .A2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n711), .B(G303), .ZN(new_n929));
  XNOR2_X1  g504(.A(G305), .B(G290), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n929), .B(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT42), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n931), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n931), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(KEYINPUT108), .B2(KEYINPUT42), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(new_n922), .A3(new_n927), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(KEYINPUT108), .A3(KEYINPUT42), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n935), .B(new_n938), .C1(new_n932), .C2(new_n933), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(G868), .A3(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT109), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G868), .ZN(new_n945));
  AOI21_X1  g520(.A(KEYINPUT109), .B1(new_n862), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n942), .B2(new_n946), .ZN(G295));
  AOI21_X1  g522(.A(new_n944), .B1(new_n942), .B2(new_n946), .ZN(G331));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n923), .A2(new_n926), .ZN(new_n950));
  NAND2_X1  g525(.A1(G77), .A2(G543), .ZN(new_n951));
  INV_X1    g526(.A(G64), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n951), .B1(new_n553), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(G651), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n954), .A2(KEYINPUT110), .A3(new_n547), .A4(new_n548), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT110), .ZN(new_n956));
  NAND2_X1  g531(.A1(G301), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n957), .A3(G286), .ZN(new_n958));
  NAND3_X1  g533(.A1(G168), .A2(G171), .A3(KEYINPUT110), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n868), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT111), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n863), .A2(new_n958), .A3(new_n867), .A4(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n869), .A2(KEYINPUT111), .A3(new_n959), .A4(new_n958), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n961), .A2(new_n963), .ZN(new_n967));
  OAI22_X1  g542(.A1(new_n950), .A2(new_n966), .B1(new_n921), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n931), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n924), .A2(new_n918), .A3(new_n915), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n966), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n923), .A2(new_n926), .A3(new_n967), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(new_n936), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n969), .A2(new_n906), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n949), .B1(new_n974), .B2(KEYINPUT43), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n936), .B1(new_n971), .B2(new_n972), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT112), .B1(new_n976), .B2(G37), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n923), .A2(new_n926), .A3(new_n967), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n921), .B1(new_n964), .B2(new_n965), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n931), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT112), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n980), .A2(new_n981), .A3(new_n906), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n977), .A2(new_n973), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n975), .B1(new_n983), .B2(KEYINPUT43), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT113), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(KEYINPUT43), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT43), .ZN(new_n987));
  AND4_X1   g562(.A1(new_n987), .A2(new_n969), .A3(new_n906), .A4(new_n973), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n985), .B1(new_n990), .B2(new_n949), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n988), .B1(new_n983), .B2(KEYINPUT43), .ZN(new_n992));
  NOR3_X1   g567(.A1(new_n992), .A2(KEYINPUT113), .A3(KEYINPUT44), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n984), .B1(new_n991), .B2(new_n993), .ZN(G397));
  NOR2_X1   g569(.A1(G290), .A2(G1986), .ZN(new_n995));
  XNOR2_X1  g570(.A(new_n995), .B(KEYINPUT115), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT114), .B(G1384), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(new_n492), .B2(new_n504), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n471), .A2(new_n477), .A3(G40), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n996), .A2(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(G1986), .A3(G290), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XOR2_X1   g580(.A(new_n1005), .B(KEYINPUT116), .Z(new_n1006));
  INV_X1    g581(.A(new_n1002), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n833), .B(new_n835), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n757), .B(G1996), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(new_n731), .B(new_n733), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n1011), .B(KEYINPUT117), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1007), .B1(new_n1010), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1006), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(G1976), .ZN(new_n1015));
  INV_X1    g590(.A(G1384), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(new_n492), .B2(new_n504), .ZN(new_n1017));
  OAI221_X1 g592(.A(G8), .B1(G288), .B2(new_n1015), .C1(new_n1001), .C2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n711), .A2(G1976), .ZN(new_n1019));
  OR3_X1    g594(.A1(new_n1018), .A2(KEYINPUT52), .A3(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(G305), .A2(G1981), .ZN(new_n1021));
  INV_X1    g596(.A(G1981), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n586), .A2(new_n1022), .A3(new_n591), .A4(new_n593), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1017), .A2(new_n1001), .ZN(new_n1027));
  INV_X1    g602(.A(G8), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1021), .A2(KEYINPUT49), .A3(new_n1023), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT120), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1032), .B1(new_n1018), .B2(KEYINPUT52), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1018), .A2(new_n1032), .A3(KEYINPUT52), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1020), .B(new_n1031), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT45), .B1(new_n515), .B2(new_n1016), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n471), .A2(new_n477), .A3(G40), .ZN(new_n1037));
  OAI211_X1 g612(.A(KEYINPUT45), .B(new_n997), .C1(new_n492), .C2(new_n504), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT118), .B1(new_n1036), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1041));
  INV_X1    g616(.A(KEYINPUT118), .ZN(new_n1042));
  AOI21_X1  g617(.A(G1384), .B1(new_n505), .B2(new_n514), .ZN(new_n1043));
  OAI211_X1 g618(.A(new_n1041), .B(new_n1042), .C1(KEYINPUT45), .C2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1040), .A2(new_n708), .A3(new_n1044), .ZN(new_n1045));
  AOI211_X1 g620(.A(KEYINPUT50), .B(G1384), .C1(new_n505), .C2(new_n514), .ZN(new_n1046));
  AOI21_X1  g621(.A(G1384), .B1(new_n885), .B2(new_n511), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1037), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(G2090), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1045), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(G8), .ZN(new_n1054));
  NAND2_X1  g629(.A1(G303), .A2(G8), .ZN(new_n1055));
  XNOR2_X1  g630(.A(new_n1055), .B(KEYINPUT55), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1035), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI211_X1 g632(.A(new_n999), .B(G1384), .C1(new_n505), .C2(new_n514), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1037), .B1(new_n1047), .B2(KEYINPUT45), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1061), .A2(G2078), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1001), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1063), .B1(new_n1043), .B2(new_n1048), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1060), .A2(new_n1062), .B1(new_n1064), .B2(new_n764), .ZN(new_n1065));
  AOI21_X1  g640(.A(G2078), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1065), .B1(new_n1066), .B2(KEYINPUT53), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(G171), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1068), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1037), .B1(KEYINPUT50), .B2(new_n1017), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n515), .A2(new_n1016), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1071), .B2(KEYINPUT50), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n1051), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1028), .B1(new_n1045), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  INV_X1    g650(.A(new_n1056), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1075), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1078));
  OAI211_X1 g653(.A(new_n1057), .B(new_n1069), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(G1966), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1081));
  INV_X1    g656(.A(G2084), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1063), .B(new_n1082), .C1(new_n1048), .C2(new_n1043), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  NOR2_X1   g659(.A1(G168), .A2(new_n1028), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1028), .B1(new_n1081), .B2(new_n1083), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1089), .B2(new_n1085), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1088), .B(KEYINPUT51), .C1(new_n1089), .C2(new_n1085), .ZN(new_n1093));
  AOI211_X1 g668(.A(KEYINPUT62), .B(new_n1087), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT125), .B1(new_n1079), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1020), .A2(new_n1031), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1034), .A2(new_n1033), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1028), .B1(new_n1045), .B2(new_n1052), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1098), .B1(new_n1076), .B2(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT119), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1100), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT62), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1086), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT125), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1104), .A2(new_n1107), .A3(new_n1108), .A4(new_n1069), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1086), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1110), .A2(KEYINPUT62), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n1095), .A2(new_n1109), .A3(new_n1111), .ZN(new_n1112));
  AND2_X1   g687(.A1(new_n1089), .A2(G168), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1057), .B(new_n1113), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT63), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1098), .A2(KEYINPUT63), .A3(new_n1113), .ZN(new_n1117));
  OR2_X1    g692(.A1(new_n1074), .A2(new_n1076), .ZN(new_n1118));
  OAI211_X1 g693(.A(new_n1117), .B(new_n1118), .C1(new_n1078), .C2(new_n1077), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1116), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT54), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n471), .A2(G40), .A3(new_n1062), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT123), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n477), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n477), .A2(new_n1123), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1125), .A2(new_n1000), .A3(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1064), .A2(new_n764), .B1(new_n1127), .B2(new_n1038), .ZN(new_n1128));
  OAI211_X1 g703(.A(G301), .B(new_n1128), .C1(new_n1066), .C2(KEYINPUT53), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1129), .A2(KEYINPUT124), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n1068), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1129), .A2(KEYINPUT124), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1121), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1128), .B1(new_n1066), .B2(KEYINPUT53), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1121), .B1(new_n1134), .B2(G171), .ZN(new_n1135));
  OAI211_X1 g710(.A(G301), .B(new_n1065), .C1(new_n1066), .C2(KEYINPUT53), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1105), .A2(new_n1086), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n844), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT57), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n577), .A2(new_n1139), .A3(new_n580), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT57), .B1(new_n618), .B2(new_n619), .ZN(new_n1141));
  AND2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g717(.A(KEYINPUT56), .B(G2072), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1041), .B(new_n1143), .C1(KEYINPUT45), .C2(new_n1043), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1138), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1027), .A2(new_n835), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1146), .B1(new_n1072), .B2(G1348), .ZN(new_n1147));
  AND2_X1   g722(.A1(new_n1147), .A2(new_n614), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1142), .B1(new_n1138), .B2(new_n1144), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1145), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT60), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n613), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  OAI211_X1 g727(.A(KEYINPUT60), .B(new_n1146), .C1(new_n1072), .C2(G1348), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1138), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1155), .B1(new_n1156), .B2(new_n1149), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1138), .A2(new_n1144), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1142), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(new_n1145), .A3(KEYINPUT61), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1154), .A2(new_n1157), .A3(new_n1161), .ZN(new_n1162));
  XOR2_X1   g737(.A(KEYINPUT121), .B(KEYINPUT59), .Z(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1036), .A2(new_n1039), .ZN(new_n1165));
  INV_X1    g740(.A(G1996), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1027), .ZN(new_n1167));
  XOR2_X1   g742(.A(KEYINPUT58), .B(G1341), .Z(new_n1168));
  AOI22_X1  g743(.A1(new_n1165), .A2(new_n1166), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1164), .B1(new_n1169), .B2(new_n559), .ZN(new_n1170));
  NOR3_X1   g745(.A1(new_n1036), .A2(G1996), .A3(new_n1039), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1172));
  OAI211_X1 g747(.A(new_n560), .B(new_n1163), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  OAI211_X1 g748(.A(new_n1170), .B(new_n1173), .C1(new_n1153), .C2(new_n1152), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1150), .B1(new_n1162), .B2(new_n1174), .ZN(new_n1175));
  NAND4_X1  g750(.A1(new_n1133), .A2(new_n1137), .A3(new_n1104), .A4(new_n1175), .ZN(new_n1176));
  NOR3_X1   g751(.A1(new_n1077), .A2(new_n1078), .A3(new_n1035), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1031), .A2(new_n1015), .A3(new_n711), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1023), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1177), .B1(new_n1029), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1120), .A2(new_n1176), .A3(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1014), .B1(new_n1112), .B2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1010), .A2(new_n733), .A3(new_n731), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n828), .A2(new_n835), .A3(new_n832), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1007), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(KEYINPUT48), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1013), .B1(new_n1186), .B2(new_n1003), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n996), .A2(KEYINPUT48), .A3(new_n1002), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1185), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1007), .B1(new_n1008), .B2(new_n757), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT46), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1002), .A2(new_n1166), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1190), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1192), .A2(new_n1191), .ZN(new_n1194));
  XNOR2_X1  g769(.A(new_n1194), .B(KEYINPUT126), .ZN(new_n1195));
  NAND2_X1  g770(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NOR2_X1   g771(.A1(new_n1196), .A2(KEYINPUT47), .ZN(new_n1197));
  AND2_X1   g772(.A1(new_n1196), .A2(KEYINPUT47), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1189), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT127), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1182), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g776(.A1(new_n461), .A2(G227), .ZN(new_n1203));
  AND3_X1   g777(.A1(new_n700), .A2(new_n661), .A3(new_n1203), .ZN(new_n1204));
  OAI211_X1 g778(.A(new_n1204), .B(new_n990), .C1(new_n907), .C2(new_n908), .ZN(G225));
  INV_X1    g779(.A(G225), .ZN(G308));
endmodule


