

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751;

  NOR2_X1 U368 ( .A1(n676), .A2(n722), .ZN(n679) );
  NOR2_X1 U369 ( .A1(n669), .A2(n722), .ZN(n671) );
  NOR2_X1 U370 ( .A1(G902), .A2(n673), .ZN(n534) );
  NOR2_X1 U371 ( .A1(G953), .A2(G237), .ZN(n524) );
  INV_X2 U372 ( .A(G953), .ZN(n739) );
  XNOR2_X2 U373 ( .A(n620), .B(KEYINPUT108), .ZN(n582) );
  XNOR2_X2 U374 ( .A(n534), .B(G472), .ZN(n620) );
  AND2_X2 U375 ( .A1(n379), .A2(n693), .ZN(n449) );
  NAND2_X1 U376 ( .A1(n366), .A2(n347), .ZN(n370) );
  INV_X1 U377 ( .A(n348), .ZN(n347) );
  NOR2_X1 U378 ( .A1(n374), .A2(n373), .ZN(n348) );
  XNOR2_X2 U379 ( .A(n478), .B(n425), .ZN(n424) );
  AND2_X1 U380 ( .A1(n535), .A2(n431), .ZN(n353) );
  XNOR2_X2 U381 ( .A(n523), .B(n360), .ZN(n535) );
  AND2_X1 U382 ( .A1(n616), .A2(n617), .ZN(n622) );
  NOR2_X2 U383 ( .A1(G902), .A2(n706), .ZN(n472) );
  INV_X1 U384 ( .A(KEYINPUT0), .ZN(n349) );
  XNOR2_X1 U385 ( .A(n388), .B(KEYINPUT39), .ZN(n379) );
  XNOR2_X1 U386 ( .A(n424), .B(n483), .ZN(n423) );
  BUF_X1 U387 ( .A(n656), .Z(n434) );
  OR2_X1 U388 ( .A1(n657), .A2(n658), .ZN(n408) );
  INV_X1 U389 ( .A(n751), .ZN(n402) );
  NOR2_X1 U390 ( .A1(n573), .A2(n572), .ZN(n700) );
  NOR2_X1 U391 ( .A1(n641), .A2(n555), .ZN(n540) );
  NAND2_X1 U392 ( .A1(n574), .A2(KEYINPUT70), .ZN(n403) );
  XNOR2_X1 U393 ( .A(n423), .B(n422), .ZN(n664) );
  XNOR2_X1 U394 ( .A(n518), .B(n414), .ZN(n549) );
  XNOR2_X1 U395 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U396 ( .A(n477), .B(n466), .ZN(n533) );
  XOR2_X1 U397 ( .A(G146), .B(G125), .Z(n476) );
  XNOR2_X1 U398 ( .A(KEYINPUT65), .B(G101), .ZN(n527) );
  XNOR2_X1 U399 ( .A(G137), .B(KEYINPUT66), .ZN(n467) );
  NOR2_X2 U400 ( .A1(n368), .A2(n375), .ZN(n390) );
  XNOR2_X1 U401 ( .A(n349), .B(n536), .ZN(n555) );
  NOR2_X2 U402 ( .A1(n712), .A2(n722), .ZN(n713) );
  INV_X1 U403 ( .A(KEYINPUT4), .ZN(n465) );
  INV_X1 U404 ( .A(n631), .ZN(n377) );
  INV_X1 U405 ( .A(KEYINPUT30), .ZN(n376) );
  XNOR2_X1 U406 ( .A(G131), .B(G134), .ZN(n466) );
  INV_X1 U407 ( .A(n656), .ZN(n412) );
  NOR2_X1 U408 ( .A1(n654), .A2(n386), .ZN(n662) );
  XNOR2_X1 U409 ( .A(n608), .B(n387), .ZN(n386) );
  INV_X1 U410 ( .A(KEYINPUT83), .ZN(n387) );
  XNOR2_X1 U411 ( .A(G110), .B(G104), .ZN(n462) );
  XNOR2_X1 U412 ( .A(n533), .B(n467), .ZN(n737) );
  NAND2_X1 U413 ( .A1(n402), .A2(KEYINPUT46), .ZN(n395) );
  NAND2_X1 U414 ( .A1(n751), .A2(n417), .ZN(n391) );
  XOR2_X1 U415 ( .A(G116), .B(KEYINPUT5), .Z(n526) );
  XNOR2_X1 U416 ( .A(n476), .B(n358), .ZN(n425) );
  INV_X1 U417 ( .A(KEYINPUT79), .ZN(n384) );
  NAND2_X1 U418 ( .A1(n621), .A2(n622), .ZN(n552) );
  OR2_X1 U419 ( .A1(G237), .A2(G902), .ZN(n485) );
  INV_X1 U420 ( .A(n403), .ZN(n373) );
  NAND2_X1 U421 ( .A1(n403), .A2(n356), .ZN(n371) );
  INV_X1 U422 ( .A(KEYINPUT70), .ZN(n404) );
  OR2_X1 U423 ( .A1(n720), .A2(G902), .ZN(n447) );
  XNOR2_X1 U424 ( .A(n460), .B(n461), .ZN(n446) );
  XNOR2_X1 U425 ( .A(n475), .B(n530), .ZN(n724) );
  XNOR2_X1 U426 ( .A(n453), .B(n467), .ZN(n441) );
  XNOR2_X1 U427 ( .A(n439), .B(n438), .ZN(n437) );
  XNOR2_X1 U428 ( .A(KEYINPUT78), .B(KEYINPUT23), .ZN(n438) );
  XNOR2_X1 U429 ( .A(n440), .B(G128), .ZN(n439) );
  INV_X1 U430 ( .A(G119), .ZN(n440) );
  NOR2_X2 U431 ( .A1(n663), .A2(n662), .ZN(n714) );
  NAND2_X1 U432 ( .A1(n411), .A2(n363), .ZN(n410) );
  XOR2_X1 U433 ( .A(KEYINPUT87), .B(n542), .Z(n573) );
  XNOR2_X1 U434 ( .A(n443), .B(n442), .ZN(n570) );
  INV_X1 U435 ( .A(KEYINPUT109), .ZN(n442) );
  INV_X1 U436 ( .A(n581), .ZN(n444) );
  XNOR2_X1 U437 ( .A(n620), .B(n385), .ZN(n569) );
  INV_X1 U438 ( .A(KEYINPUT6), .ZN(n385) );
  INV_X1 U439 ( .A(n569), .ZN(n429) );
  INV_X1 U440 ( .A(n542), .ZN(n430) );
  XNOR2_X1 U441 ( .A(n737), .B(n451), .ZN(n706) );
  XOR2_X1 U442 ( .A(G146), .B(G140), .Z(n469) );
  NOR2_X1 U443 ( .A1(G952), .A2(n739), .ZN(n722) );
  INV_X1 U444 ( .A(KEYINPUT104), .ZN(n381) );
  INV_X1 U445 ( .A(KEYINPUT48), .ZN(n400) );
  NAND2_X1 U446 ( .A1(n403), .A2(n357), .ZN(n372) );
  NAND2_X1 U447 ( .A1(G234), .A2(G237), .ZN(n488) );
  XNOR2_X1 U448 ( .A(n604), .B(KEYINPUT38), .ZN(n632) );
  NOR2_X1 U449 ( .A1(n593), .A2(n569), .ZN(n445) );
  INV_X1 U450 ( .A(KEYINPUT89), .ZN(n435) );
  XNOR2_X1 U451 ( .A(KEYINPUT15), .B(G902), .ZN(n436) );
  XNOR2_X1 U452 ( .A(n528), .B(n527), .ZN(n416) );
  XOR2_X1 U453 ( .A(G116), .B(G122), .Z(n502) );
  XNOR2_X1 U454 ( .A(KEYINPUT102), .B(KEYINPUT100), .ZN(n496) );
  XOR2_X1 U455 ( .A(KEYINPUT101), .B(KEYINPUT7), .Z(n497) );
  XNOR2_X1 U456 ( .A(n482), .B(n724), .ZN(n422) );
  XNOR2_X1 U457 ( .A(n609), .B(n384), .ZN(n383) );
  INV_X1 U458 ( .A(n570), .ZN(n598) );
  XNOR2_X1 U459 ( .A(n539), .B(n538), .ZN(n641) );
  NOR2_X1 U460 ( .A1(n552), .A2(n569), .ZN(n539) );
  AND2_X1 U461 ( .A1(n575), .A2(KEYINPUT70), .ZN(n375) );
  XNOR2_X1 U462 ( .A(n571), .B(n487), .ZN(n586) );
  XNOR2_X1 U463 ( .A(n486), .B(KEYINPUT71), .ZN(n487) );
  XNOR2_X1 U464 ( .A(n517), .B(G475), .ZN(n414) );
  XNOR2_X1 U465 ( .A(n441), .B(n437), .ZN(n456) );
  INV_X1 U466 ( .A(n597), .ZN(n378) );
  XNOR2_X1 U467 ( .A(n421), .B(n420), .ZN(n572) );
  INV_X1 U468 ( .A(KEYINPUT36), .ZN(n420) );
  XNOR2_X1 U469 ( .A(n364), .B(KEYINPUT32), .ZN(n749) );
  NOR2_X1 U470 ( .A1(n586), .A2(n595), .ZN(n690) );
  NOR2_X1 U471 ( .A1(n430), .A2(n429), .ZN(n428) );
  XNOR2_X1 U472 ( .A(n704), .B(n419), .ZN(n707) );
  XNOR2_X1 U473 ( .A(n415), .B(n554), .ZN(n575) );
  AND2_X1 U474 ( .A1(n606), .A2(KEYINPUT2), .ZN(n350) );
  XNOR2_X1 U475 ( .A(n436), .B(n435), .ZN(n659) );
  XNOR2_X1 U476 ( .A(n584), .B(KEYINPUT1), .ZN(n621) );
  AND2_X1 U477 ( .A1(G210), .A2(n485), .ZN(n351) );
  AND2_X1 U478 ( .A1(n380), .A2(n748), .ZN(n352) );
  OR2_X1 U479 ( .A1(KEYINPUT47), .A2(n591), .ZN(n354) );
  AND2_X1 U480 ( .A1(n377), .A2(n376), .ZN(n356) );
  NOR2_X1 U481 ( .A1(n377), .A2(n376), .ZN(n357) );
  AND2_X1 U482 ( .A1(G224), .A2(n739), .ZN(n358) );
  AND2_X1 U483 ( .A1(n405), .A2(n404), .ZN(n359) );
  XOR2_X1 U484 ( .A(n522), .B(KEYINPUT69), .Z(n360) );
  XNOR2_X1 U485 ( .A(KEYINPUT82), .B(KEYINPUT45), .ZN(n361) );
  OR2_X1 U486 ( .A1(n661), .A2(n660), .ZN(n362) );
  AND2_X1 U487 ( .A1(n362), .A2(KEYINPUT80), .ZN(n363) );
  INV_X1 U488 ( .A(KEYINPUT46), .ZN(n417) );
  INV_X1 U489 ( .A(n659), .ZN(n655) );
  NAND2_X1 U490 ( .A1(n370), .A2(n369), .ZN(n368) );
  AND2_X1 U491 ( .A1(n367), .A2(n371), .ZN(n366) );
  NAND2_X1 U492 ( .A1(n353), .A2(n562), .ZN(n364) );
  AND2_X1 U493 ( .A1(n432), .A2(n569), .ZN(n431) );
  NAND2_X1 U494 ( .A1(n365), .A2(n359), .ZN(n369) );
  INV_X1 U495 ( .A(n575), .ZN(n365) );
  OR2_X1 U496 ( .A1(n582), .A2(n372), .ZN(n367) );
  NAND2_X1 U497 ( .A1(n582), .A2(n376), .ZN(n374) );
  AND2_X1 U498 ( .A1(n379), .A2(n378), .ZN(n702) );
  XNOR2_X1 U499 ( .A(n559), .B(n381), .ZN(n380) );
  NAND2_X1 U500 ( .A1(n382), .A2(n362), .ZN(n409) );
  NAND2_X1 U501 ( .A1(n407), .A2(n408), .ZN(n382) );
  AND2_X1 U502 ( .A1(n547), .A2(n749), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n536), .B(KEYINPUT0), .ZN(n551) );
  NOR2_X2 U504 ( .A1(n586), .A2(n493), .ZN(n536) );
  INV_X1 U505 ( .A(n535), .ZN(n544) );
  NOR2_X1 U506 ( .A1(n650), .A2(n649), .ZN(n653) );
  NAND2_X1 U507 ( .A1(n383), .A2(n610), .ZN(n611) );
  NOR2_X1 U508 ( .A1(G953), .A2(n612), .ZN(n615) );
  NAND2_X2 U509 ( .A1(n607), .A2(n606), .ZN(n656) );
  NOR2_X1 U510 ( .A1(n397), .A2(n592), .ZN(n389) );
  NAND2_X1 U511 ( .A1(n607), .A2(n350), .ZN(n608) );
  XNOR2_X2 U512 ( .A(n401), .B(n400), .ZN(n607) );
  NAND2_X1 U513 ( .A1(n390), .A2(n632), .ZN(n388) );
  XNOR2_X2 U514 ( .A(n449), .B(KEYINPUT40), .ZN(n750) );
  NAND2_X1 U515 ( .A1(n399), .A2(n389), .ZN(n401) );
  NAND2_X1 U516 ( .A1(n577), .A2(n631), .ZN(n571) );
  NAND2_X1 U517 ( .A1(n390), .A2(n578), .ZN(n579) );
  NAND2_X1 U518 ( .A1(n392), .A2(n391), .ZN(n399) );
  NAND2_X1 U519 ( .A1(n394), .A2(n393), .ZN(n392) );
  NAND2_X1 U520 ( .A1(n750), .A2(KEYINPUT46), .ZN(n393) );
  NAND2_X1 U521 ( .A1(n396), .A2(n395), .ZN(n394) );
  INV_X1 U522 ( .A(n750), .ZN(n396) );
  XNOR2_X1 U523 ( .A(n700), .B(KEYINPUT85), .ZN(n398) );
  NAND2_X1 U524 ( .A1(n354), .A2(n398), .ZN(n397) );
  INV_X1 U525 ( .A(n574), .ZN(n405) );
  NAND2_X1 U526 ( .A1(n406), .A2(n657), .ZN(n407) );
  NOR2_X1 U527 ( .A1(n656), .A2(n413), .ZN(n406) );
  NAND2_X1 U528 ( .A1(n409), .A2(n410), .ZN(n663) );
  NAND2_X1 U529 ( .A1(n412), .A2(n655), .ZN(n411) );
  OR2_X1 U530 ( .A1(n659), .A2(KEYINPUT80), .ZN(n413) );
  NAND2_X1 U531 ( .A1(n584), .A2(n622), .ZN(n415) );
  XNOR2_X2 U532 ( .A(n472), .B(n471), .ZN(n584) );
  XNOR2_X1 U533 ( .A(n529), .B(n416), .ZN(n531) );
  NAND2_X1 U534 ( .A1(n445), .A2(n444), .ZN(n443) );
  NOR2_X1 U535 ( .A1(n570), .A2(n571), .ZN(n421) );
  XNOR2_X1 U536 ( .A(n450), .B(KEYINPUT44), .ZN(n427) );
  NAND2_X1 U537 ( .A1(n418), .A2(n576), .ZN(n541) );
  XNOR2_X1 U538 ( .A(n540), .B(KEYINPUT34), .ZN(n418) );
  XNOR2_X2 U539 ( .A(n463), .B(n462), .ZN(n723) );
  XOR2_X2 U540 ( .A(n723), .B(n464), .Z(n483) );
  XNOR2_X1 U541 ( .A(n706), .B(n705), .ZN(n419) );
  INV_X1 U542 ( .A(n577), .ZN(n604) );
  XNOR2_X2 U543 ( .A(n484), .B(n351), .ZN(n577) );
  INV_X1 U544 ( .A(n657), .ZN(n654) );
  XNOR2_X2 U545 ( .A(n426), .B(n361), .ZN(n657) );
  NAND2_X1 U546 ( .A1(n427), .A2(n352), .ZN(n426) );
  NAND2_X1 U547 ( .A1(n535), .A2(n428), .ZN(n560) );
  INV_X1 U548 ( .A(n573), .ZN(n432) );
  XNOR2_X1 U549 ( .A(n433), .B(G143), .ZN(G45) );
  XNOR2_X1 U550 ( .A(n433), .B(n580), .ZN(n589) );
  XNOR2_X2 U551 ( .A(n579), .B(KEYINPUT112), .ZN(n433) );
  XNOR2_X1 U552 ( .A(n434), .B(n741), .ZN(n740) );
  INV_X1 U553 ( .A(n617), .ZN(n562) );
  XNOR2_X2 U554 ( .A(n447), .B(n446), .ZN(n617) );
  XNOR2_X2 U555 ( .A(n448), .B(G143), .ZN(n499) );
  XNOR2_X2 U556 ( .A(G128), .B(KEYINPUT73), .ZN(n448) );
  XNOR2_X1 U557 ( .A(n483), .B(n470), .ZN(n451) );
  BUF_X1 U558 ( .A(n714), .Z(n718) );
  NOR2_X2 U559 ( .A1(n550), .A2(n549), .ZN(n693) );
  INV_X1 U560 ( .A(KEYINPUT77), .ZN(n580) );
  XNOR2_X1 U561 ( .A(n502), .B(KEYINPUT16), .ZN(n475) );
  INV_X1 U562 ( .A(KEYINPUT80), .ZN(n658) );
  INV_X1 U563 ( .A(KEYINPUT97), .ZN(n554) );
  INV_X1 U564 ( .A(n477), .ZN(n478) );
  XNOR2_X1 U565 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U566 ( .A(n703), .ZN(n605) );
  INV_X1 U567 ( .A(KEYINPUT22), .ZN(n522) );
  XNOR2_X1 U568 ( .A(n533), .B(n532), .ZN(n673) );
  NOR2_X1 U569 ( .A1(n702), .A2(n605), .ZN(n606) );
  INV_X1 U570 ( .A(KEYINPUT59), .ZN(n708) );
  XNOR2_X1 U571 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U572 ( .A(n675), .B(n674), .ZN(n676) );
  INV_X1 U573 ( .A(KEYINPUT53), .ZN(n651) );
  XNOR2_X1 U574 ( .A(n677), .B(KEYINPUT88), .ZN(n678) );
  XNOR2_X1 U575 ( .A(n653), .B(n652), .ZN(G75) );
  XNOR2_X1 U576 ( .A(n476), .B(KEYINPUT10), .ZN(n452) );
  XNOR2_X1 U577 ( .A(n452), .B(G140), .ZN(n736) );
  XNOR2_X1 U578 ( .A(G110), .B(KEYINPUT24), .ZN(n453) );
  NAND2_X1 U579 ( .A1(G234), .A2(n739), .ZN(n454) );
  XOR2_X1 U580 ( .A(KEYINPUT8), .B(n454), .Z(n503) );
  NAND2_X1 U581 ( .A1(G221), .A2(n503), .ZN(n455) );
  XNOR2_X1 U582 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U583 ( .A(n736), .B(n457), .ZN(n720) );
  NAND2_X1 U584 ( .A1(n659), .A2(G234), .ZN(n459) );
  XNOR2_X1 U585 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n458) );
  XNOR2_X1 U586 ( .A(n459), .B(n458), .ZN(n494) );
  NAND2_X1 U587 ( .A1(G217), .A2(n494), .ZN(n460) );
  XOR2_X1 U588 ( .A(KEYINPUT25), .B(KEYINPUT72), .Z(n461) );
  XOR2_X1 U589 ( .A(KEYINPUT90), .B(G107), .Z(n463) );
  INV_X1 U590 ( .A(n527), .ZN(n464) );
  XNOR2_X2 U591 ( .A(n499), .B(n465), .ZN(n477) );
  NAND2_X1 U592 ( .A1(G227), .A2(n739), .ZN(n468) );
  XNOR2_X1 U593 ( .A(n469), .B(n468), .ZN(n470) );
  XNOR2_X1 U594 ( .A(KEYINPUT67), .B(G469), .ZN(n471) );
  INV_X1 U595 ( .A(n621), .ZN(n542) );
  XOR2_X1 U596 ( .A(G119), .B(KEYINPUT91), .Z(n474) );
  XNOR2_X1 U597 ( .A(G113), .B(KEYINPUT3), .ZN(n473) );
  XNOR2_X1 U598 ( .A(n474), .B(n473), .ZN(n530) );
  XOR2_X1 U599 ( .A(KEYINPUT93), .B(KEYINPUT92), .Z(n480) );
  XNOR2_X1 U600 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n479) );
  XNOR2_X1 U601 ( .A(n480), .B(n479), .ZN(n481) );
  XOR2_X1 U602 ( .A(KEYINPUT86), .B(n481), .Z(n482) );
  NAND2_X1 U603 ( .A1(n664), .A2(n659), .ZN(n484) );
  NAND2_X1 U604 ( .A1(G214), .A2(n485), .ZN(n631) );
  XNOR2_X1 U605 ( .A(KEYINPUT19), .B(KEYINPUT64), .ZN(n486) );
  XNOR2_X1 U606 ( .A(n488), .B(KEYINPUT94), .ZN(n489) );
  XNOR2_X1 U607 ( .A(KEYINPUT14), .B(n489), .ZN(n490) );
  NAND2_X1 U608 ( .A1(G952), .A2(n490), .ZN(n647) );
  NOR2_X1 U609 ( .A1(G953), .A2(n647), .ZN(n566) );
  NAND2_X1 U610 ( .A1(G902), .A2(n490), .ZN(n563) );
  NOR2_X1 U611 ( .A1(G898), .A2(n739), .ZN(n491) );
  XNOR2_X1 U612 ( .A(KEYINPUT95), .B(n491), .ZN(n727) );
  NOR2_X1 U613 ( .A1(n563), .A2(n727), .ZN(n492) );
  NOR2_X1 U614 ( .A1(n566), .A2(n492), .ZN(n493) );
  NAND2_X1 U615 ( .A1(G221), .A2(n494), .ZN(n495) );
  XOR2_X1 U616 ( .A(KEYINPUT21), .B(n495), .Z(n616) );
  INV_X1 U617 ( .A(n616), .ZN(n537) );
  XNOR2_X1 U618 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U619 ( .A(KEYINPUT9), .B(n498), .Z(n501) );
  XNOR2_X1 U620 ( .A(n499), .B(G107), .ZN(n500) );
  XNOR2_X1 U621 ( .A(n501), .B(n500), .ZN(n507) );
  XOR2_X1 U622 ( .A(G134), .B(n502), .Z(n505) );
  NAND2_X1 U623 ( .A1(G217), .A2(n503), .ZN(n504) );
  XNOR2_X1 U624 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U625 ( .A(n507), .B(n506), .ZN(n716) );
  NOR2_X1 U626 ( .A1(G902), .A2(n716), .ZN(n508) );
  XNOR2_X1 U627 ( .A(G478), .B(n508), .ZN(n548) );
  XNOR2_X1 U628 ( .A(G113), .B(KEYINPUT12), .ZN(n509) );
  XNOR2_X1 U629 ( .A(n509), .B(KEYINPUT11), .ZN(n513) );
  XOR2_X1 U630 ( .A(G104), .B(G122), .Z(n511) );
  XNOR2_X1 U631 ( .A(G131), .B(G143), .ZN(n510) );
  XNOR2_X1 U632 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U633 ( .A(n512), .B(n513), .Z(n515) );
  NAND2_X1 U634 ( .A1(G214), .A2(n524), .ZN(n514) );
  XNOR2_X1 U635 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U636 ( .A(n736), .B(n516), .ZN(n709) );
  NOR2_X1 U637 ( .A1(G902), .A2(n709), .ZN(n518) );
  XNOR2_X1 U638 ( .A(KEYINPUT99), .B(KEYINPUT13), .ZN(n517) );
  AND2_X1 U639 ( .A1(n548), .A2(n549), .ZN(n519) );
  XNOR2_X1 U640 ( .A(n519), .B(KEYINPUT105), .ZN(n634) );
  NOR2_X1 U641 ( .A1(n537), .A2(n634), .ZN(n520) );
  XNOR2_X1 U642 ( .A(KEYINPUT106), .B(n520), .ZN(n521) );
  NAND2_X1 U643 ( .A1(n551), .A2(n521), .ZN(n523) );
  NAND2_X1 U644 ( .A1(n524), .A2(G210), .ZN(n525) );
  XNOR2_X1 U645 ( .A(n526), .B(n525), .ZN(n529) );
  XNOR2_X1 U646 ( .A(G137), .B(G146), .ZN(n528) );
  XNOR2_X1 U647 ( .A(KEYINPUT33), .B(KEYINPUT68), .ZN(n538) );
  NOR2_X1 U648 ( .A1(n549), .A2(n548), .ZN(n576) );
  XNOR2_X1 U649 ( .A(n541), .B(KEYINPUT35), .ZN(n747) );
  NAND2_X1 U650 ( .A1(n542), .A2(n582), .ZN(n543) );
  NOR2_X1 U651 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U652 ( .A1(n545), .A2(n562), .ZN(n687) );
  INV_X1 U653 ( .A(n687), .ZN(n546) );
  NOR2_X1 U654 ( .A1(n747), .A2(n546), .ZN(n547) );
  INV_X1 U655 ( .A(n548), .ZN(n550) );
  INV_X1 U656 ( .A(n693), .ZN(n593) );
  AND2_X1 U657 ( .A1(n550), .A2(n549), .ZN(n696) );
  XNOR2_X1 U658 ( .A(KEYINPUT103), .B(n696), .ZN(n597) );
  NAND2_X1 U659 ( .A1(n593), .A2(n597), .ZN(n587) );
  INV_X1 U660 ( .A(n587), .ZN(n636) );
  NOR2_X1 U661 ( .A1(n620), .A2(n552), .ZN(n627) );
  NAND2_X1 U662 ( .A1(n551), .A2(n627), .ZN(n553) );
  XNOR2_X1 U663 ( .A(n553), .B(KEYINPUT31), .ZN(n697) );
  NAND2_X1 U664 ( .A1(n365), .A2(n620), .ZN(n556) );
  NOR2_X1 U665 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U666 ( .A(n557), .B(KEYINPUT98), .ZN(n681) );
  NOR2_X1 U667 ( .A1(n697), .A2(n681), .ZN(n558) );
  NOR2_X1 U668 ( .A1(n636), .A2(n558), .ZN(n559) );
  NOR2_X1 U669 ( .A1(n560), .A2(n562), .ZN(n561) );
  XNOR2_X1 U670 ( .A(n561), .B(KEYINPUT107), .ZN(n748) );
  OR2_X1 U671 ( .A1(n739), .A2(n563), .ZN(n564) );
  NOR2_X1 U672 ( .A1(G900), .A2(n564), .ZN(n565) );
  NOR2_X1 U673 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U674 ( .A(KEYINPUT74), .B(n567), .ZN(n574) );
  NOR2_X1 U675 ( .A1(n617), .A2(n574), .ZN(n568) );
  NAND2_X1 U676 ( .A1(n568), .A2(n616), .ZN(n581) );
  AND2_X1 U677 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U678 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U679 ( .A(KEYINPUT28), .B(n583), .ZN(n585) );
  NAND2_X1 U680 ( .A1(n585), .A2(n584), .ZN(n595) );
  NAND2_X1 U681 ( .A1(n690), .A2(n587), .ZN(n591) );
  NAND2_X1 U682 ( .A1(n591), .A2(KEYINPUT47), .ZN(n588) );
  NAND2_X1 U683 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U684 ( .A(n590), .B(KEYINPUT76), .ZN(n592) );
  NAND2_X1 U685 ( .A1(n632), .A2(n631), .ZN(n635) );
  NOR2_X1 U686 ( .A1(n635), .A2(n634), .ZN(n594) );
  XNOR2_X1 U687 ( .A(n594), .B(KEYINPUT41), .ZN(n630) );
  NOR2_X1 U688 ( .A1(n630), .A2(n595), .ZN(n596) );
  XNOR2_X1 U689 ( .A(n596), .B(KEYINPUT42), .ZN(n751) );
  NAND2_X1 U690 ( .A1(n598), .A2(n631), .ZN(n599) );
  NOR2_X1 U691 ( .A1(n430), .A2(n599), .ZN(n602) );
  XNOR2_X1 U692 ( .A(KEYINPUT43), .B(KEYINPUT110), .ZN(n600) );
  XNOR2_X1 U693 ( .A(n600), .B(KEYINPUT111), .ZN(n601) );
  XNOR2_X1 U694 ( .A(n602), .B(n601), .ZN(n603) );
  NAND2_X1 U695 ( .A1(n604), .A2(n603), .ZN(n703) );
  INV_X1 U696 ( .A(KEYINPUT2), .ZN(n661) );
  NAND2_X1 U697 ( .A1(n434), .A2(n661), .ZN(n609) );
  NAND2_X1 U698 ( .A1(n654), .A2(n661), .ZN(n610) );
  NOR2_X1 U699 ( .A1(n662), .A2(n611), .ZN(n612) );
  NOR2_X1 U700 ( .A1(n630), .A2(n641), .ZN(n613) );
  XOR2_X1 U701 ( .A(KEYINPUT122), .B(n613), .Z(n614) );
  NAND2_X1 U702 ( .A1(n615), .A2(n614), .ZN(n650) );
  NOR2_X1 U703 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U704 ( .A(n618), .B(KEYINPUT49), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n620), .A2(n619), .ZN(n625) );
  NOR2_X1 U706 ( .A1(n622), .A2(n430), .ZN(n623) );
  XNOR2_X1 U707 ( .A(n623), .B(KEYINPUT50), .ZN(n624) );
  NOR2_X1 U708 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U709 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U710 ( .A(KEYINPUT51), .B(n628), .Z(n629) );
  NOR2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n643) );
  NOR2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U713 ( .A1(n634), .A2(n633), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT119), .B(n637), .Z(n638) );
  NOR2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n640) );
  NOR2_X1 U717 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  XNOR2_X1 U719 ( .A(n644), .B(KEYINPUT120), .ZN(n645) );
  XNOR2_X1 U720 ( .A(KEYINPUT52), .B(n645), .ZN(n646) );
  NOR2_X1 U721 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X1 U722 ( .A(n648), .B(KEYINPUT121), .Z(n649) );
  XNOR2_X1 U723 ( .A(n651), .B(KEYINPUT123), .ZN(n652) );
  XOR2_X1 U724 ( .A(KEYINPUT81), .B(n659), .Z(n660) );
  NAND2_X1 U725 ( .A1(n714), .A2(G210), .ZN(n668) );
  XOR2_X1 U726 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n666) );
  XNOR2_X1 U727 ( .A(n664), .B(KEYINPUT75), .ZN(n665) );
  XNOR2_X1 U728 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U729 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U730 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n670) );
  XNOR2_X1 U731 ( .A(n671), .B(n670), .ZN(G51) );
  NAND2_X1 U732 ( .A1(n714), .A2(G472), .ZN(n675) );
  XOR2_X1 U733 ( .A(KEYINPUT113), .B(KEYINPUT62), .Z(n672) );
  INV_X1 U734 ( .A(KEYINPUT63), .ZN(n677) );
  XNOR2_X1 U735 ( .A(n679), .B(n678), .ZN(G57) );
  NAND2_X1 U736 ( .A1(n681), .A2(n693), .ZN(n680) );
  XNOR2_X1 U737 ( .A(n680), .B(G104), .ZN(G6) );
  XOR2_X1 U738 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n683) );
  NAND2_X1 U739 ( .A1(n696), .A2(n681), .ZN(n682) );
  XNOR2_X1 U740 ( .A(n683), .B(n682), .ZN(n684) );
  XOR2_X1 U741 ( .A(n684), .B(KEYINPUT26), .Z(n686) );
  XNOR2_X1 U742 ( .A(G107), .B(KEYINPUT114), .ZN(n685) );
  XNOR2_X1 U743 ( .A(n686), .B(n685), .ZN(G9) );
  XNOR2_X1 U744 ( .A(G110), .B(n687), .ZN(G12) );
  XOR2_X1 U745 ( .A(G128), .B(KEYINPUT29), .Z(n689) );
  NAND2_X1 U746 ( .A1(n690), .A2(n696), .ZN(n688) );
  XNOR2_X1 U747 ( .A(n689), .B(n688), .ZN(G30) );
  NAND2_X1 U748 ( .A1(n690), .A2(n693), .ZN(n691) );
  XNOR2_X1 U749 ( .A(n691), .B(KEYINPUT116), .ZN(n692) );
  XNOR2_X1 U750 ( .A(G146), .B(n692), .ZN(G48) );
  XOR2_X1 U751 ( .A(G113), .B(KEYINPUT117), .Z(n695) );
  NAND2_X1 U752 ( .A1(n697), .A2(n693), .ZN(n694) );
  XNOR2_X1 U753 ( .A(n695), .B(n694), .ZN(G15) );
  NAND2_X1 U754 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U755 ( .A(n698), .B(KEYINPUT118), .ZN(n699) );
  XNOR2_X1 U756 ( .A(G116), .B(n699), .ZN(G18) );
  XNOR2_X1 U757 ( .A(G125), .B(n700), .ZN(n701) );
  XNOR2_X1 U758 ( .A(n701), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U759 ( .A(G134), .B(n702), .Z(G36) );
  XNOR2_X1 U760 ( .A(G140), .B(n703), .ZN(G42) );
  XOR2_X1 U761 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n705) );
  NAND2_X1 U762 ( .A1(n718), .A2(G469), .ZN(n704) );
  NOR2_X1 U763 ( .A1(n722), .A2(n707), .ZN(G54) );
  NAND2_X1 U764 ( .A1(n714), .A2(G475), .ZN(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(n710), .ZN(n712) );
  XNOR2_X1 U766 ( .A(KEYINPUT60), .B(n713), .ZN(G60) );
  NAND2_X1 U767 ( .A1(G478), .A2(n718), .ZN(n715) );
  XNOR2_X1 U768 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U769 ( .A1(n722), .A2(n717), .ZN(G63) );
  NAND2_X1 U770 ( .A1(G217), .A2(n718), .ZN(n719) );
  XNOR2_X1 U771 ( .A(n720), .B(n719), .ZN(n721) );
  NOR2_X1 U772 ( .A1(n722), .A2(n721), .ZN(G66) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(n725) );
  XNOR2_X1 U774 ( .A(n725), .B(KEYINPUT125), .ZN(n726) );
  XNOR2_X1 U775 ( .A(G101), .B(n726), .ZN(n728) );
  NAND2_X1 U776 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U777 ( .A(n729), .B(KEYINPUT124), .ZN(n735) );
  NAND2_X1 U778 ( .A1(G953), .A2(G224), .ZN(n730) );
  XNOR2_X1 U779 ( .A(KEYINPUT61), .B(n730), .ZN(n731) );
  NAND2_X1 U780 ( .A1(n731), .A2(G898), .ZN(n733) );
  OR2_X1 U781 ( .A1(n654), .A2(G953), .ZN(n732) );
  NAND2_X1 U782 ( .A1(n733), .A2(n732), .ZN(n734) );
  XOR2_X1 U783 ( .A(n735), .B(n734), .Z(G69) );
  XOR2_X1 U784 ( .A(n737), .B(n736), .Z(n738) );
  XOR2_X1 U785 ( .A(KEYINPUT126), .B(n738), .Z(n741) );
  NAND2_X1 U786 ( .A1(n740), .A2(n739), .ZN(n746) );
  XNOR2_X1 U787 ( .A(G227), .B(n741), .ZN(n742) );
  NAND2_X1 U788 ( .A1(n742), .A2(G900), .ZN(n743) );
  XOR2_X1 U789 ( .A(KEYINPUT127), .B(n743), .Z(n744) );
  NAND2_X1 U790 ( .A1(G953), .A2(n744), .ZN(n745) );
  NAND2_X1 U791 ( .A1(n746), .A2(n745), .ZN(G72) );
  XOR2_X1 U792 ( .A(G122), .B(n747), .Z(G24) );
  XNOR2_X1 U793 ( .A(G101), .B(n748), .ZN(G3) );
  XNOR2_X1 U794 ( .A(n749), .B(G119), .ZN(G21) );
  XOR2_X1 U795 ( .A(n750), .B(G131), .Z(G33) );
  XOR2_X1 U796 ( .A(G137), .B(n751), .Z(G39) );
endmodule

