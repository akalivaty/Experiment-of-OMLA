//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 1 0 1 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1 1 1 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:22 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1016, new_n1017;
  XNOR2_X1  g000(.A(G1gat), .B(G29gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT0), .ZN(new_n203));
  XNOR2_X1  g002(.A(G57gat), .B(G85gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G225gat), .A2(G233gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(G113gat), .B(G120gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  XNOR2_X1  g008(.A(G127gat), .B(G134gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT1), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT67), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g013(.A(new_n210), .B(new_n212), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G155gat), .A2(G162gat), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  INV_X1    g017(.A(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n220), .B2(KEYINPUT2), .ZN(new_n221));
  INV_X1    g020(.A(G148gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  INV_X1    g022(.A(G141gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G148gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT76), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n222), .A2(KEYINPUT76), .A3(G141gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n221), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G141gat), .B(G148gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n217), .B(new_n220), .C1(new_n230), .C2(KEYINPUT2), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n232), .ZN(new_n233));
  AND2_X1   g032(.A1(new_n229), .A2(new_n231), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n214), .A2(new_n215), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n207), .B1(new_n233), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT5), .ZN(new_n238));
  OAI21_X1  g037(.A(KEYINPUT79), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT79), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n235), .B(new_n232), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n240), .B(KEYINPUT5), .C1(new_n241), .C2(new_n207), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT4), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n234), .A2(new_n244), .A3(new_n235), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n244), .B1(new_n234), .B2(new_n235), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n207), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n229), .A2(new_n231), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n248), .B1(new_n229), .B2(new_n231), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n216), .B(new_n249), .C1(new_n250), .C2(KEYINPUT77), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(KEYINPUT77), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g052(.A(KEYINPUT78), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n250), .A2(KEYINPUT77), .ZN(new_n255));
  INV_X1    g054(.A(new_n249), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n256), .A2(new_n235), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT78), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n255), .A2(new_n257), .A3(new_n258), .A4(new_n252), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n247), .B1(new_n254), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n243), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n254), .A2(new_n259), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n246), .B1(new_n245), .B2(KEYINPUT80), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT80), .ZN(new_n264));
  OAI21_X1  g063(.A(new_n264), .B1(new_n236), .B2(KEYINPUT4), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n207), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(KEYINPUT5), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n262), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n206), .B1(new_n261), .B2(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n254), .A2(new_n259), .B1(new_n263), .B2(new_n265), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n271), .A2(new_n268), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n272), .B(new_n205), .C1(new_n260), .C2(new_n243), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT81), .B(KEYINPUT6), .Z(new_n274));
  NAND3_X1  g073(.A1(new_n270), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n274), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n206), .B(new_n276), .C1(new_n261), .C2(new_n269), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n272), .B1(new_n260), .B2(new_n243), .ZN(new_n280));
  NAND4_X1  g079(.A1(new_n280), .A2(KEYINPUT82), .A3(new_n206), .A4(new_n276), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n283));
  NAND2_X1  g082(.A1(G226gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(G169gat), .ZN(new_n288));
  INV_X1    g087(.A(G176gat), .ZN(new_n289));
  OAI22_X1  g088(.A1(new_n288), .A2(new_n289), .B1(KEYINPUT64), .B2(KEYINPUT23), .ZN(new_n290));
  AND2_X1   g089(.A1(KEYINPUT64), .A2(KEYINPUT23), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n287), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT65), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n294), .A2(KEYINPUT23), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n298), .A2(KEYINPUT66), .ZN(new_n299));
  OR2_X1    g098(.A1(G183gat), .A2(G190gat), .ZN(new_n300));
  NAND3_X1  g099(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT66), .ZN(new_n302));
  OAI211_X1 g101(.A(new_n300), .B(new_n301), .C1(new_n297), .C2(new_n302), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n292), .B(new_n296), .C1(new_n299), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT25), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT27), .B(G183gat), .ZN(new_n306));
  INV_X1    g105(.A(G190gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n308), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n288), .A2(new_n289), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n310), .B1(KEYINPUT26), .B2(new_n287), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n295), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n311), .B1(KEYINPUT26), .B2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n306), .A2(new_n314), .A3(new_n307), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n309), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT25), .B1(new_n286), .B2(KEYINPUT23), .ZN(new_n317));
  AND2_X1   g116(.A1(new_n292), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n298), .A2(new_n300), .A3(new_n301), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n305), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT29), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n285), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(KEYINPUT25), .A2(new_n304), .B1(new_n318), .B2(new_n319), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n284), .B1(new_n324), .B2(new_n316), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(G197gat), .ZN(new_n327));
  INV_X1    g126(.A(G204gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(G197gat), .A2(G204gat), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT22), .ZN(new_n331));
  NAND2_X1  g130(.A1(G211gat), .A2(G218gat), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n329), .A2(new_n330), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT72), .ZN(new_n334));
  XNOR2_X1  g133(.A(G211gat), .B(G218gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n334), .B1(new_n333), .B2(new_n335), .ZN(new_n338));
  OAI22_X1  g137(.A1(new_n337), .A2(new_n338), .B1(new_n335), .B2(new_n333), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT73), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n333), .A2(new_n335), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n333), .A2(new_n335), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT72), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n343), .B2(new_n336), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n283), .B1(new_n326), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n321), .A2(new_n322), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n284), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n321), .A2(new_n351), .A3(new_n285), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n351), .B1(new_n321), .B2(new_n285), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n350), .B(new_n339), .C1(new_n352), .C2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n347), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n355), .B(KEYINPUT74), .C1(new_n323), .C2(new_n325), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n348), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(G8gat), .B(G36gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(G64gat), .B(G92gat), .ZN(new_n359));
  XOR2_X1   g158(.A(new_n358), .B(new_n359), .Z(new_n360));
  INV_X1    g159(.A(new_n360), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n357), .A2(KEYINPUT30), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(new_n356), .ZN(new_n363));
  INV_X1    g162(.A(new_n325), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n350), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g164(.A(KEYINPUT74), .B1(new_n365), .B2(new_n355), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n361), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n348), .A2(new_n354), .A3(new_n356), .A4(new_n360), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT30), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n362), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n282), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT86), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n282), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT35), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(G228gat), .A2(G233gat), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n337), .A2(new_n338), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n341), .A2(KEYINPUT84), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT84), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n333), .B2(new_n335), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n322), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n234), .B1(new_n384), .B2(new_n248), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n249), .A2(new_n322), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n344), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n378), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n248), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(new_n232), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n340), .A2(new_n346), .A3(new_n386), .ZN(new_n392));
  INV_X1    g191(.A(new_n378), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(G22gat), .ZN(new_n395));
  AND3_X1   g194(.A1(new_n389), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n395), .B1(new_n389), .B2(new_n394), .ZN(new_n397));
  XNOR2_X1  g196(.A(G78gat), .B(G106gat), .ZN(new_n398));
  INV_X1    g197(.A(G50gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n396), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n400), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n380), .A2(new_n382), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n343), .A2(new_n336), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT29), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n232), .B1(new_n405), .B2(KEYINPUT3), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n393), .B1(new_n406), .B2(new_n387), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(new_n393), .ZN(new_n408));
  OAI21_X1  g207(.A(G22gat), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n394), .A3(new_n395), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n402), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n377), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n321), .A2(new_n235), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n324), .A2(new_n216), .A3(new_n316), .ZN(new_n414));
  INV_X1    g213(.A(G227gat), .ZN(new_n415));
  INV_X1    g214(.A(G233gat), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT32), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT33), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(G15gat), .B(G43gat), .Z(new_n422));
  XNOR2_X1  g221(.A(G71gat), .B(G99gat), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n419), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n424), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n418), .B(KEYINPUT32), .C1(new_n420), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n417), .B1(new_n413), .B2(new_n414), .ZN(new_n429));
  XNOR2_X1  g228(.A(KEYINPUT68), .B(KEYINPUT34), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT34), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(KEYINPUT68), .ZN(new_n433));
  AOI211_X1 g232(.A(new_n417), .B(new_n433), .C1(new_n413), .C2(new_n414), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n431), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g234(.A(new_n428), .B(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n400), .B1(new_n396), .B2(new_n397), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n409), .A2(new_n402), .A3(new_n410), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n437), .A2(new_n376), .A3(new_n438), .ZN(new_n439));
  AND4_X1   g238(.A1(new_n375), .A2(new_n412), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n372), .A2(new_n374), .A3(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT69), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n431), .A2(new_n434), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n430), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n216), .B1(new_n324), .B2(new_n316), .ZN(new_n445));
  AND4_X1   g244(.A1(new_n216), .A2(new_n305), .A3(new_n316), .A4(new_n320), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n444), .B1(new_n447), .B2(new_n417), .ZN(new_n448));
  INV_X1    g247(.A(new_n433), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(KEYINPUT69), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n428), .B1(new_n443), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(KEYINPUT70), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n442), .B1(new_n431), .B2(new_n434), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n448), .A2(new_n450), .A3(KEYINPUT69), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT70), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n456), .A2(new_n457), .A3(new_n428), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n435), .A2(new_n425), .A3(new_n427), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n459), .A2(new_n439), .A3(new_n412), .A4(new_n460), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT35), .B1(new_n461), .B2(new_n371), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n441), .A2(new_n462), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n412), .A2(new_n439), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT39), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n465), .B1(new_n241), .B2(new_n207), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n271), .B2(new_n207), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n262), .A2(new_n266), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n468), .A2(new_n465), .A3(new_n267), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n467), .A2(new_n469), .A3(new_n205), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT40), .ZN(new_n471));
  AOI22_X1  g270(.A1(new_n470), .A2(new_n471), .B1(new_n280), .B2(new_n206), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT40), .A4(new_n205), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n472), .A2(new_n362), .A3(new_n369), .A4(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(new_n344), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(KEYINPUT85), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT85), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n475), .A2(new_n478), .A3(new_n344), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n326), .A2(new_n347), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n477), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(KEYINPUT37), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT38), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n361), .A2(KEYINPUT37), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n367), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n361), .B1(new_n357), .B2(KEYINPUT37), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT38), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n275), .A2(new_n279), .A3(new_n281), .A4(new_n368), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n464), .B(new_n474), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n456), .A2(new_n457), .A3(new_n428), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n457), .B1(new_n456), .B2(new_n428), .ZN(new_n494));
  OAI211_X1 g293(.A(KEYINPUT36), .B(new_n460), .C1(new_n493), .C2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n428), .B1(new_n431), .B2(new_n434), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(new_n460), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT36), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT71), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n459), .A2(KEYINPUT71), .A3(KEYINPUT36), .A4(new_n460), .ZN(new_n501));
  AOI22_X1  g300(.A1(new_n282), .A2(new_n370), .B1(new_n412), .B2(new_n439), .ZN(new_n502));
  INV_X1    g301(.A(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n492), .A2(new_n500), .A3(new_n501), .A4(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n463), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(G15gat), .B(G22gat), .ZN(new_n506));
  INV_X1    g305(.A(G1gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT16), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n509), .B1(G1gat), .B2(new_n506), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G8gat), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n509), .B(new_n512), .C1(G1gat), .C2(new_n506), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT92), .ZN(new_n516));
  AND2_X1   g315(.A1(G57gat), .A2(G64gat), .ZN(new_n517));
  NOR2_X1   g316(.A1(G57gat), .A2(G64gat), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G57gat), .ZN(new_n520));
  INV_X1    g319(.A(G64gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G57gat), .A2(G64gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT92), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT9), .ZN(new_n525));
  INV_X1    g324(.A(G71gat), .ZN(new_n526));
  INV_X1    g325(.A(G78gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT91), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT91), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(G71gat), .B2(G78gat), .ZN(new_n530));
  AOI22_X1  g329(.A1(new_n528), .A2(new_n530), .B1(G71gat), .B2(G78gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n517), .A2(new_n518), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT9), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(new_n526), .B2(new_n527), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n525), .A2(new_n531), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n515), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT94), .ZN(new_n538));
  INV_X1    g337(.A(new_n538), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n537), .A2(KEYINPUT94), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n535), .A2(KEYINPUT21), .ZN(new_n542));
  XNOR2_X1  g341(.A(G127gat), .B(G155gat), .ZN(new_n543));
  XOR2_X1   g342(.A(new_n542), .B(new_n543), .Z(new_n544));
  OR2_X1    g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n541), .A2(new_n544), .ZN(new_n546));
  AND2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(G231gat), .A2(G233gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT93), .ZN(new_n549));
  XOR2_X1   g348(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G183gat), .B(G211gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n547), .B(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555));
  INV_X1    g354(.A(G36gat), .ZN(new_n556));
  AND2_X1   g355(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n556), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G29gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n560), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G43gat), .A2(G50gat), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g363(.A1(G43gat), .A2(G50gat), .ZN(new_n565));
  OAI21_X1  g364(.A(KEYINPUT15), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OR2_X1    g365(.A1(G43gat), .A2(G50gat), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT15), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n567), .A2(new_n568), .A3(new_n563), .ZN(new_n569));
  NAND4_X1  g368(.A1(new_n562), .A2(KEYINPUT87), .A3(new_n566), .A4(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n566), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(new_n559), .A3(new_n561), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n566), .A2(new_n569), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT87), .B1(new_n574), .B2(new_n562), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n555), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT14), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n560), .ZN(new_n578));
  NAND2_X1  g377(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n579));
  AOI21_X1  g378(.A(G36gat), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n561), .ZN(new_n581));
  OAI211_X1 g380(.A(new_n566), .B(new_n569), .C1(new_n580), .C2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT87), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n584), .A2(KEYINPUT17), .A3(new_n572), .A4(new_n570), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n576), .A2(new_n515), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G229gat), .A2(G233gat), .ZN(new_n587));
  XOR2_X1   g386(.A(new_n587), .B(KEYINPUT88), .Z(new_n588));
  INV_X1    g387(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n584), .A2(new_n572), .A3(new_n570), .ZN(new_n590));
  AND3_X1   g389(.A1(new_n590), .A2(KEYINPUT89), .A3(new_n514), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT89), .B1(new_n590), .B2(new_n514), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n586), .B(new_n589), .C1(new_n591), .C2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT18), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n590), .A2(new_n514), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT89), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n590), .A2(KEYINPUT89), .A3(new_n514), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(KEYINPUT18), .A3(new_n589), .A4(new_n586), .ZN(new_n601));
  XNOR2_X1  g400(.A(G113gat), .B(G141gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n602), .B(G197gat), .ZN(new_n603));
  XOR2_X1   g402(.A(KEYINPUT11), .B(G169gat), .Z(new_n604));
  XNOR2_X1  g403(.A(new_n603), .B(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(KEYINPUT12), .ZN(new_n606));
  OR2_X1    g405(.A1(new_n590), .A2(new_n514), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n607), .B1(new_n591), .B2(new_n592), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n588), .B(KEYINPUT13), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n595), .A2(new_n601), .A3(new_n606), .A4(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT90), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n593), .A2(new_n594), .B1(new_n608), .B2(new_n610), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n606), .B1(new_n614), .B2(new_n601), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n613), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT8), .ZN(new_n618));
  OR2_X1    g417(.A1(G85gat), .A2(G92gat), .ZN(new_n619));
  AND2_X1   g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT96), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(KEYINPUT7), .ZN(new_n624));
  AND2_X1   g423(.A1(G85gat), .A2(G92gat), .ZN(new_n625));
  AND3_X1   g424(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n625), .B1(new_n622), .B2(new_n624), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n620), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(G99gat), .A2(G106gat), .ZN(new_n629));
  NOR2_X1   g428(.A1(G99gat), .A2(G106gat), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n631), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n633), .B(new_n620), .C1(new_n626), .C2(new_n627), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n576), .A2(new_n585), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G190gat), .B(G218gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n637), .B(KEYINPUT97), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT41), .ZN(new_n639));
  NAND2_X1  g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT95), .ZN(new_n641));
  OAI22_X1  g440(.A1(new_n638), .A2(KEYINPUT98), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n635), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n642), .B1(new_n643), .B2(new_n590), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n636), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n638), .A2(KEYINPUT98), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n641), .A2(new_n639), .ZN(new_n648));
  XOR2_X1   g447(.A(G134gat), .B(G162gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  OR2_X1    g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n650), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT101), .ZN(new_n655));
  NAND2_X1  g454(.A1(G230gat), .A2(G233gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n525), .A2(new_n531), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n534), .A2(new_n532), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n634), .B(new_n632), .C1(new_n659), .C2(KEYINPUT99), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n634), .A2(KEYINPUT99), .ZN(new_n661));
  INV_X1    g460(.A(new_n625), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n623), .A2(KEYINPUT7), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n621), .A2(KEYINPUT96), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n622), .A2(new_n624), .A3(new_n625), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g466(.A(new_n633), .B1(new_n667), .B2(new_n620), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n618), .A2(new_n619), .ZN(new_n669));
  AOI211_X1 g468(.A(new_n631), .B(new_n669), .C1(new_n665), .C2(new_n666), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n661), .B(new_n535), .C1(new_n668), .C2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT10), .B1(new_n660), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT10), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n635), .A2(new_n673), .A3(new_n659), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n656), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  AND2_X1   g474(.A1(new_n660), .A2(new_n671), .ZN(new_n676));
  INV_X1    g475(.A(new_n656), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g477(.A(G120gat), .B(G148gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT100), .ZN(new_n680));
  XNOR2_X1  g479(.A(G176gat), .B(G204gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n675), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n682), .B1(new_n675), .B2(new_n678), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n655), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n675), .A2(new_n678), .ZN(new_n687));
  INV_X1    g486(.A(new_n682), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n689), .A2(KEYINPUT101), .A3(new_n683), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR4_X1   g491(.A1(new_n554), .A2(new_n616), .A3(new_n654), .A4(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n505), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g493(.A1(new_n275), .A2(new_n279), .A3(new_n281), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(G1gat), .ZN(G1324gat));
  INV_X1    g496(.A(new_n694), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT102), .B(KEYINPUT16), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G8gat), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n698), .A2(new_n370), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(new_n370), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n512), .B1(new_n694), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g502(.A(KEYINPUT42), .B1(new_n701), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(KEYINPUT42), .B2(new_n701), .ZN(G1325gat));
  OR3_X1    g504(.A1(new_n698), .A2(G15gat), .A3(new_n497), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n500), .A2(new_n501), .ZN(new_n707));
  OAI21_X1  g506(.A(G15gat), .B1(new_n698), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n706), .A2(new_n708), .ZN(G1326gat));
  NAND2_X1  g508(.A1(new_n412), .A2(new_n439), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g510(.A(KEYINPUT43), .B(G22gat), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n711), .B(new_n712), .ZN(G1327gat));
  AND2_X1   g512(.A1(new_n472), .A2(new_n473), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(new_n702), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n695), .A2(new_n368), .A3(new_n486), .A4(new_n489), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n502), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI22_X1  g516(.A1(new_n717), .A2(new_n707), .B1(new_n441), .B2(new_n462), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n718), .A2(new_n653), .ZN(new_n719));
  INV_X1    g518(.A(new_n554), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n616), .A3(new_n692), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n560), .A3(new_n695), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT45), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n726), .B1(new_n718), .B2(new_n653), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n505), .A2(KEYINPUT44), .A3(new_n654), .ZN(new_n728));
  AND2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n721), .ZN(new_n730));
  OAI21_X1  g529(.A(G29gat), .B1(new_n730), .B2(new_n282), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n725), .A2(new_n731), .ZN(G1328gat));
  NOR3_X1   g531(.A1(new_n722), .A2(G36gat), .A3(new_n370), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(KEYINPUT46), .ZN(new_n734));
  OAI21_X1  g533(.A(G36gat), .B1(new_n730), .B2(new_n370), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n734), .A2(new_n735), .ZN(G1329gat));
  INV_X1    g535(.A(new_n707), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n727), .A2(new_n728), .A3(new_n737), .A4(new_n721), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(G43gat), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n497), .A2(G43gat), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n723), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n739), .A2(new_n741), .A3(KEYINPUT47), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n739), .A2(KEYINPUT103), .B1(new_n723), .B2(new_n740), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT103), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n738), .A2(new_n744), .A3(G43gat), .ZN(new_n745));
  AOI211_X1 g544(.A(KEYINPUT104), .B(KEYINPUT47), .C1(new_n743), .C2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n739), .A2(KEYINPUT103), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n748), .A2(new_n745), .A3(new_n741), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT47), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n742), .B1(new_n746), .B2(new_n751), .ZN(G1330gat));
  OAI21_X1  g551(.A(G50gat), .B1(new_n730), .B2(new_n464), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT48), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n723), .A2(new_n399), .A3(new_n710), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n755), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n753), .B(new_n756), .C1(new_n754), .C2(KEYINPUT48), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1331gat));
  XNOR2_X1  g559(.A(new_n695), .B(KEYINPUT106), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n613), .A2(new_n615), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT90), .B(new_n606), .C1(new_n614), .C2(new_n601), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR4_X1   g563(.A1(new_n554), .A2(new_n764), .A3(new_n654), .A4(new_n691), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n505), .A2(new_n761), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g566(.A1(new_n505), .A2(new_n765), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n370), .ZN(new_n769));
  NOR2_X1   g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  AND2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n772), .B1(new_n769), .B2(new_n770), .ZN(G1333gat));
  OAI21_X1  g572(.A(G71gat), .B1(new_n768), .B2(new_n707), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n436), .A2(new_n526), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n774), .B1(new_n768), .B2(new_n775), .ZN(new_n776));
  XOR2_X1   g575(.A(new_n776), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g576(.A1(new_n768), .A2(new_n464), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n778), .B(new_n527), .ZN(G1335gat));
  INV_X1    g578(.A(KEYINPUT108), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n554), .A2(new_n616), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(KEYINPUT107), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n719), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n784), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n719), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n782), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n785), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n282), .A2(G85gat), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n788), .A2(new_n692), .A3(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n782), .A2(new_n692), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n729), .A2(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(G85gat), .B1(new_n792), .B2(new_n282), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n793), .ZN(G1336gat));
  NOR3_X1   g593(.A1(new_n370), .A2(G92gat), .A3(new_n691), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n788), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n729), .A2(new_n702), .A3(new_n791), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G92gat), .ZN(new_n798));
  XNOR2_X1  g597(.A(KEYINPUT110), .B(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n783), .B(new_n784), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n795), .B(KEYINPUT109), .Z(new_n802));
  AOI22_X1  g601(.A1(new_n801), .A2(new_n802), .B1(new_n797), .B2(G92gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n796), .A2(new_n800), .B1(new_n803), .B2(new_n804), .ZN(G1337gat));
  NOR2_X1   g604(.A1(new_n497), .A2(G99gat), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n692), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n792), .B2(new_n707), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT111), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n807), .A2(KEYINPUT111), .A3(new_n808), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(G1338gat));
  NOR3_X1   g612(.A1(new_n464), .A2(G106gat), .A3(new_n691), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n788), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n729), .A2(new_n710), .A3(new_n791), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G106gat), .ZN(new_n817));
  XNOR2_X1  g616(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n801), .A2(new_n814), .B1(new_n816), .B2(G106gat), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT53), .ZN(new_n821));
  OAI22_X1  g620(.A1(new_n815), .A2(new_n819), .B1(new_n820), .B2(new_n821), .ZN(G1339gat));
  NAND2_X1  g621(.A1(new_n464), .A2(new_n436), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n825), .B(new_n656), .C1(new_n672), .C2(new_n674), .ZN(new_n826));
  AND2_X1   g625(.A1(new_n826), .A2(new_n688), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n672), .A2(new_n656), .A3(new_n674), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT113), .ZN(new_n829));
  OAI211_X1 g628(.A(KEYINPUT54), .B(new_n675), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n674), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n677), .B(new_n831), .C1(new_n676), .C2(KEYINPUT10), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  OAI211_X1 g632(.A(KEYINPUT55), .B(new_n827), .C1(new_n830), .C2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n683), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n672), .A2(new_n674), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n837), .A2(new_n829), .A3(new_n677), .ZN(new_n838));
  NAND4_X1  g637(.A1(new_n836), .A2(KEYINPUT54), .A3(new_n838), .A4(new_n675), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT55), .B1(new_n839), .B2(new_n827), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n824), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n827), .B1(new_n830), .B2(new_n833), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT55), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n844), .A2(KEYINPUT114), .A3(new_n683), .A4(new_n834), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n764), .A3(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n608), .B2(new_n610), .ZN(new_n849));
  NAND4_X1  g648(.A1(new_n600), .A2(KEYINPUT115), .A3(new_n607), .A4(new_n609), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n588), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n849), .A2(new_n850), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(new_n605), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n612), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n691), .A2(new_n855), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n846), .A2(new_n847), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n847), .B1(new_n846), .B2(new_n856), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n857), .A2(new_n858), .A3(new_n654), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n653), .A2(new_n855), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n841), .A2(new_n860), .A3(new_n845), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n554), .B1(new_n859), .B2(new_n862), .ZN(new_n863));
  NAND4_X1  g662(.A1(new_n720), .A2(new_n616), .A3(new_n653), .A4(new_n691), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n823), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n702), .A2(new_n282), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g666(.A(G113gat), .ZN(new_n868));
  NOR3_X1   g667(.A1(new_n867), .A2(new_n868), .A3(new_n616), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n846), .A2(new_n856), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n654), .B1(new_n870), .B2(KEYINPUT116), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n846), .A2(new_n847), .A3(new_n856), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n862), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n864), .B1(new_n873), .B2(new_n720), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n874), .A2(new_n370), .A3(new_n761), .ZN(new_n875));
  INV_X1    g674(.A(new_n461), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n878), .A2(new_n764), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n869), .B1(new_n879), .B2(new_n868), .ZN(G1340gat));
  INV_X1    g679(.A(G120gat), .ZN(new_n881));
  NOR3_X1   g680(.A1(new_n867), .A2(new_n881), .A3(new_n691), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n878), .A2(new_n692), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n881), .ZN(G1341gat));
  NAND4_X1  g683(.A1(new_n865), .A2(G127gat), .A3(new_n720), .A4(new_n866), .ZN(new_n885));
  XNOR2_X1  g684(.A(new_n885), .B(KEYINPUT117), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n877), .A2(KEYINPUT118), .A3(new_n554), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n887), .A2(G127gat), .ZN(new_n888));
  OAI21_X1  g687(.A(KEYINPUT118), .B1(new_n877), .B2(new_n554), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G1342gat));
  NOR2_X1   g689(.A1(new_n653), .A2(G134gat), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n878), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g691(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  OAI21_X1  g694(.A(G134gat), .B1(new_n867), .B2(new_n653), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(G1343gat));
  NOR2_X1   g696(.A1(new_n737), .A2(new_n464), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n875), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n224), .B1(new_n899), .B2(new_n616), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n707), .A2(new_n866), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT57), .B1(new_n874), .B2(new_n710), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT57), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n464), .A2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  NOR2_X1   g704(.A1(new_n691), .A2(new_n855), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n835), .A2(new_n840), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n906), .B1(new_n907), .B2(new_n764), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n861), .B1(new_n908), .B2(new_n654), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT120), .B1(new_n909), .B2(new_n554), .ZN(new_n910));
  NOR4_X1   g709(.A1(new_n554), .A2(new_n764), .A3(new_n654), .A4(new_n692), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n909), .A2(KEYINPUT120), .A3(new_n554), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n905), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n901), .B1(new_n902), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n764), .A2(G141gat), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n900), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT58), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n900), .B(KEYINPUT58), .C1(new_n915), .C2(new_n916), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1344gat));
  AOI21_X1  g720(.A(new_n905), .B1(new_n863), .B2(new_n864), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n844), .A2(new_n683), .A3(new_n834), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n856), .B1(new_n616), .B2(new_n923), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n924), .A2(new_n653), .B1(new_n860), .B2(new_n907), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n864), .B1(new_n925), .B2(new_n720), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n464), .B1(new_n926), .B2(KEYINPUT122), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n928), .B(new_n864), .C1(new_n925), .C2(new_n720), .ZN(new_n929));
  AOI21_X1  g728(.A(KEYINPUT57), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n922), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n901), .A2(new_n692), .ZN(new_n932));
  OAI21_X1  g731(.A(G148gat), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n933), .A2(KEYINPUT59), .ZN(new_n934));
  OAI211_X1 g733(.A(new_n692), .B(new_n901), .C1(new_n902), .C2(new_n914), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n222), .A2(KEYINPUT59), .ZN(new_n936));
  AND3_X1   g735(.A1(new_n935), .A2(KEYINPUT121), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(KEYINPUT121), .B1(new_n935), .B2(new_n936), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n934), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NAND4_X1  g738(.A1(new_n875), .A2(new_n222), .A3(new_n692), .A4(new_n898), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(new_n940), .ZN(G1345gat));
  NOR3_X1   g740(.A1(new_n915), .A2(new_n218), .A3(new_n554), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n899), .A2(new_n554), .ZN(new_n943));
  OR2_X1    g742(.A1(new_n943), .A2(KEYINPUT123), .ZN(new_n944));
  AOI21_X1  g743(.A(G155gat), .B1(new_n943), .B2(KEYINPUT123), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1346gat));
  NOR3_X1   g745(.A1(new_n915), .A2(new_n219), .A3(new_n653), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n875), .A2(new_n654), .A3(new_n898), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n947), .B1(new_n219), .B2(new_n948), .ZN(G1347gat));
  OR3_X1    g748(.A1(new_n761), .A2(KEYINPUT124), .A3(new_n370), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT124), .B1(new_n761), .B2(new_n370), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n865), .A2(new_n952), .ZN(new_n953));
  NOR3_X1   g752(.A1(new_n953), .A2(new_n288), .A3(new_n616), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n702), .A2(new_n282), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n955), .B1(new_n863), .B2(new_n864), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n876), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n958), .A2(new_n764), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n954), .B1(new_n288), .B2(new_n959), .ZN(G1348gat));
  OAI21_X1  g759(.A(G176gat), .B1(new_n953), .B2(new_n691), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n692), .A2(new_n289), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n961), .B1(new_n957), .B2(new_n962), .ZN(G1349gat));
  OAI21_X1  g762(.A(G183gat), .B1(new_n953), .B2(new_n554), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n720), .A2(new_n306), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n964), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  XNOR2_X1  g765(.A(new_n966), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g766(.A1(new_n958), .A2(new_n307), .A3(new_n654), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n865), .A2(new_n654), .A3(new_n952), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n969), .A2(new_n970), .A3(G190gat), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n970), .B1(new_n969), .B2(G190gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1351gat));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n898), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G197gat), .B1(new_n975), .B2(new_n764), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n931), .A2(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n931), .A2(KEYINPUT125), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n952), .A2(new_n707), .ZN(new_n979));
  AND3_X1   g778(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(new_n616), .A2(new_n327), .ZN(new_n981));
  AOI21_X1  g780(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(G1352gat));
  NAND4_X1  g781(.A1(new_n977), .A2(new_n692), .A3(new_n978), .A4(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G204gat), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT62), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n692), .A2(new_n328), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n974), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n989));
  XNOR2_X1  g788(.A(new_n988), .B(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n984), .A2(new_n990), .ZN(G1353gat));
  INV_X1    g790(.A(G211gat), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n975), .A2(new_n992), .A3(new_n720), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n950), .A2(new_n707), .A3(new_n720), .A4(new_n951), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n922), .B2(new_n930), .ZN(new_n996));
  AOI21_X1  g795(.A(KEYINPUT63), .B1(new_n996), .B2(G211gat), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n998));
  NAND3_X1  g797(.A1(new_n998), .A2(new_n653), .A3(new_n872), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n720), .B1(new_n999), .B2(new_n861), .ZN(new_n1000));
  OAI21_X1  g799(.A(new_n904), .B1(new_n1000), .B2(new_n911), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n907), .A2(new_n860), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1002), .B1(new_n908), .B2(new_n654), .ZN(new_n1003));
  AOI21_X1  g802(.A(new_n911), .B1(new_n1003), .B2(new_n554), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n710), .B1(new_n1004), .B2(new_n928), .ZN(new_n1005));
  INV_X1    g804(.A(new_n929), .ZN(new_n1006));
  OAI21_X1  g805(.A(new_n903), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g806(.A(new_n994), .B1(new_n1001), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT63), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n1008), .A2(new_n1009), .A3(new_n992), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n993), .B1(new_n997), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n1011), .A2(KEYINPUT127), .ZN(new_n1012));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n1013));
  OAI211_X1 g812(.A(new_n993), .B(new_n1013), .C1(new_n997), .C2(new_n1010), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1012), .A2(new_n1014), .ZN(G1354gat));
  AOI21_X1  g814(.A(G218gat), .B1(new_n975), .B2(new_n654), .ZN(new_n1016));
  AND2_X1   g815(.A1(new_n654), .A2(G218gat), .ZN(new_n1017));
  AOI21_X1  g816(.A(new_n1016), .B1(new_n980), .B2(new_n1017), .ZN(G1355gat));
endmodule


