//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n650, new_n651, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n678, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n826, new_n827,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n834, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G197gat), .ZN(new_n204));
  INV_X1    g003(.A(G204gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  AND2_X1   g006(.A1(G211gat), .A2(G218gat), .ZN(new_n208));
  OAI22_X1  g007(.A1(new_n206), .A2(new_n207), .B1(KEYINPUT22), .B2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(G211gat), .A2(G218gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n209), .B(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT29), .ZN(new_n213));
  AOI21_X1  g012(.A(KEYINPUT3), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT76), .B(G162gat), .ZN(new_n215));
  INV_X1    g014(.A(G155gat), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT2), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G155gat), .B(G162gat), .ZN(new_n218));
  INV_X1    g017(.A(G141gat), .ZN(new_n219));
  INV_X1    g018(.A(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G141gat), .A2(G148gat), .ZN(new_n222));
  AND2_X1   g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n217), .A2(new_n218), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT2), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n221), .A2(new_n225), .A3(new_n222), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT75), .B1(G155gat), .B2(G162gat), .ZN(new_n227));
  XOR2_X1   g026(.A(G155gat), .B(G162gat), .Z(new_n228));
  OAI211_X1 g027(.A(new_n226), .B(new_n227), .C1(new_n228), .C2(KEYINPUT75), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n230), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n214), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n224), .A2(new_n233), .A3(new_n229), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n212), .B1(new_n234), .B2(new_n213), .ZN(new_n235));
  OAI211_X1 g034(.A(G228gat), .B(G233gat), .C1(new_n232), .C2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G228gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n235), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n230), .A2(KEYINPUT78), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT78), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n240), .B1(new_n224), .B2(new_n229), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  OAI211_X1 g041(.A(new_n237), .B(new_n238), .C1(new_n242), .C2(new_n214), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n203), .B1(new_n236), .B2(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G78gat), .B(G106gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n246), .B(G22gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n236), .A2(new_n243), .A3(new_n203), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n247), .ZN(new_n250));
  INV_X1    g049(.A(new_n248), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n250), .B1(new_n251), .B2(new_n244), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n249), .A2(new_n252), .ZN(new_n253));
  OR2_X1    g052(.A1(new_n253), .A2(KEYINPUT35), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT70), .ZN(new_n255));
  NOR2_X1   g054(.A1(G169gat), .A2(G176gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(KEYINPUT26), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT26), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(G183gat), .A2(G190gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(KEYINPUT27), .B(G183gat), .ZN(new_n264));
  INV_X1    g063(.A(G190gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT28), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G183gat), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT27), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT27), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n269), .A2(G183gat), .ZN(new_n270));
  AND4_X1   g069(.A1(KEYINPUT28), .A2(new_n268), .A3(new_n270), .A4(new_n265), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n262), .B(new_n263), .C1(new_n266), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT66), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n268), .A2(new_n270), .A3(new_n265), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n264), .A2(KEYINPUT28), .A3(new_n265), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT66), .ZN(new_n279));
  NAND4_X1  g078(.A1(new_n278), .A2(new_n279), .A3(new_n263), .A4(new_n262), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT25), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n256), .A2(KEYINPUT23), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT24), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n283), .A2(G183gat), .A3(G190gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n263), .A2(KEYINPUT24), .ZN(new_n285));
  NOR2_X1   g084(.A1(G183gat), .A2(G190gat), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n282), .B(new_n284), .C1(new_n285), .C2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n261), .B1(new_n256), .B2(KEYINPUT23), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n281), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g088(.A1(new_n282), .A2(new_n284), .ZN(new_n290));
  OR2_X1    g089(.A1(new_n285), .A2(new_n286), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n261), .B(KEYINPUT65), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT23), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n281), .B1(new_n257), .B2(new_n293), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n290), .A2(new_n291), .A3(new_n292), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n280), .A3(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  OR2_X1    g097(.A1(new_n298), .A2(KEYINPUT1), .ZN(new_n299));
  XOR2_X1   g098(.A(G127gat), .B(G134gat), .Z(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  OR2_X1    g100(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n303));
  NAND4_X1  g102(.A1(new_n302), .A2(KEYINPUT68), .A3(G113gat), .A4(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n305), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT68), .B1(new_n307), .B2(G120gat), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(KEYINPUT69), .B(new_n304), .C1(new_n308), .C2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n300), .A2(KEYINPUT1), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n302), .A2(new_n303), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n309), .B1(new_n314), .B2(new_n307), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT69), .B1(new_n315), .B2(new_n304), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n301), .B1(new_n313), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n255), .B1(new_n297), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n301), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n311), .A2(new_n312), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n315), .A2(new_n304), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT69), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n319), .B1(new_n320), .B2(new_n323), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n272), .A2(KEYINPUT66), .B1(new_n289), .B2(new_n295), .ZN(new_n325));
  NAND4_X1  g124(.A1(new_n324), .A2(KEYINPUT70), .A3(new_n280), .A4(new_n325), .ZN(new_n326));
  NAND2_X1  g125(.A1(G227gat), .A2(G233gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT64), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n297), .A2(new_n317), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n318), .A2(new_n326), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  AOI21_X1  g130(.A(KEYINPUT34), .B1(new_n331), .B2(KEYINPUT71), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT32), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n318), .A2(new_n326), .A3(new_n330), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n336), .B1(new_n337), .B2(new_n328), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT33), .B1(new_n337), .B2(new_n328), .ZN(new_n339));
  XOR2_X1   g138(.A(G15gat), .B(G43gat), .Z(new_n340));
  XNOR2_X1  g139(.A(G71gat), .B(G99gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR3_X1   g142(.A1(new_n338), .A2(new_n339), .A3(new_n343), .ZN(new_n344));
  AOI221_X4 g143(.A(new_n336), .B1(KEYINPUT33), .B2(new_n342), .C1(new_n337), .C2(new_n328), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n335), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n334), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(new_n332), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n337), .A2(new_n328), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT33), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n343), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n338), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n345), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n346), .A2(new_n355), .A3(KEYINPUT73), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n353), .A2(new_n354), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n358), .A3(new_n335), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n254), .B1(new_n356), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G226gat), .A2(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n297), .A2(new_n362), .ZN(new_n363));
  OR2_X1    g162(.A1(new_n363), .A2(KEYINPUT74), .ZN(new_n364));
  AND2_X1   g163(.A1(new_n296), .A2(new_n272), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n365), .B2(KEYINPUT29), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n366), .A2(KEYINPUT74), .A3(new_n363), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(new_n212), .ZN(new_n369));
  XNOR2_X1  g168(.A(G8gat), .B(G36gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G64gat), .B(G92gat), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(new_n371), .Z(new_n372));
  NOR2_X1   g171(.A1(new_n362), .A2(KEYINPUT29), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n297), .A2(new_n373), .B1(new_n365), .B2(new_n362), .ZN(new_n374));
  INV_X1    g173(.A(new_n212), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n369), .A2(new_n372), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n372), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n364), .B2(new_n367), .ZN(new_n379));
  INV_X1    g178(.A(new_n376), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(KEYINPUT30), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT30), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n383), .A2(new_n384), .A3(new_n372), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G1gat), .B(G29gat), .ZN(new_n387));
  XNOR2_X1  g186(.A(new_n387), .B(KEYINPUT0), .ZN(new_n388));
  XNOR2_X1  g187(.A(G57gat), .B(G85gat), .ZN(new_n389));
  XOR2_X1   g188(.A(new_n388), .B(new_n389), .Z(new_n390));
  NAND3_X1  g189(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n324), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n234), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n230), .A2(KEYINPUT3), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n230), .A2(new_n392), .A3(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n395), .A2(new_n317), .A3(new_n396), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n231), .B(new_n301), .C1(new_n316), .C2(new_n313), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT4), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n391), .A2(new_n397), .A3(new_n400), .A4(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n317), .A2(new_n230), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT79), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n398), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n401), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n317), .A2(KEYINPUT79), .A3(new_n230), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n405), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n402), .A2(new_n408), .A3(KEYINPUT5), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n242), .A2(new_n399), .A3(new_n324), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n398), .A2(KEYINPUT4), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT5), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n401), .A4(new_n397), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n390), .B1(new_n409), .B2(new_n414), .ZN(new_n415));
  AND3_X1   g214(.A1(new_n415), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n416));
  AOI21_X1  g215(.A(KEYINPUT81), .B1(new_n415), .B2(KEYINPUT6), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n409), .A2(new_n414), .ZN(new_n419));
  INV_X1    g218(.A(new_n390), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT80), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n415), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT80), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n409), .A2(new_n414), .A3(new_n424), .A4(new_n390), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n421), .A2(new_n422), .A3(new_n423), .A4(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n386), .B1(new_n418), .B2(new_n426), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n360), .A2(new_n427), .A3(KEYINPUT85), .ZN(new_n428));
  AOI21_X1  g227(.A(KEYINPUT85), .B1(new_n360), .B2(new_n427), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n344), .A2(new_n345), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n253), .B1(new_n431), .B2(new_n348), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n346), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n357), .A2(KEYINPUT72), .A3(new_n335), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n432), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(KEYINPUT86), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT86), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n432), .A2(new_n434), .A3(new_n438), .A4(new_n435), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n427), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n441));
  INV_X1    g240(.A(new_n253), .ZN(new_n442));
  INV_X1    g241(.A(new_n417), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n415), .A2(KEYINPUT81), .A3(KEYINPUT6), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n426), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n386), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n442), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n382), .A2(new_n422), .A3(new_n385), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT39), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT82), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n412), .A2(new_n397), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n406), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n324), .B1(new_n394), .B2(new_n393), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n411), .A2(new_n410), .B1(new_n453), .B2(new_n396), .ZN(new_n454));
  NOR3_X1   g253(.A1(new_n454), .A2(KEYINPUT82), .A3(new_n401), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n449), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT82), .B1(new_n454), .B2(new_n401), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n451), .A2(new_n450), .A3(new_n406), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n405), .A2(new_n407), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n449), .B1(new_n459), .B2(new_n401), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n458), .A3(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n456), .A2(new_n390), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n448), .B1(new_n462), .B2(KEYINPUT40), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n456), .A2(new_n390), .A3(new_n461), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT40), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n253), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n426), .A2(new_n443), .A3(new_n444), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT37), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n369), .A2(new_n469), .A3(new_n376), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT83), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT83), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n383), .A2(new_n472), .A3(new_n469), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT84), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n475), .B(new_n378), .C1(new_n383), .C2(new_n469), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n469), .B1(new_n369), .B2(new_n376), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n477), .B2(new_n372), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n474), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(KEYINPUT38), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n368), .A2(new_n375), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n469), .B1(new_n374), .B2(new_n212), .ZN(new_n482));
  AOI211_X1 g281(.A(KEYINPUT38), .B(new_n372), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n474), .A2(new_n483), .B1(new_n372), .B2(new_n383), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n480), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n447), .B1(new_n467), .B2(new_n485), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n434), .A2(new_n435), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT36), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n431), .B2(new_n348), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n356), .A2(new_n359), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n490), .B1(KEYINPUT36), .B2(new_n491), .ZN(new_n492));
  AOI22_X1  g291(.A1(new_n430), .A2(new_n441), .B1(new_n486), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(G43gat), .B(G50gat), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n495), .A2(KEYINPUT15), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT89), .B(G29gat), .Z(new_n497));
  XNOR2_X1  g296(.A(KEYINPUT90), .B(G36gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g298(.A1(G29gat), .A2(G36gat), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n500), .B(KEYINPUT14), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n501), .B2(KEYINPUT88), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n501), .A2(KEYINPUT88), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n496), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n496), .A2(new_n501), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n505), .B(new_n499), .C1(KEYINPUT15), .C2(new_n495), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g306(.A(G15gat), .B(G22gat), .ZN(new_n508));
  INV_X1    g307(.A(G1gat), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n508), .A2(KEYINPUT16), .A3(new_n509), .ZN(new_n510));
  OR2_X1    g309(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n510), .B(new_n511), .C1(new_n509), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g311(.A1(KEYINPUT91), .A2(G8gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT17), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n507), .B(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n514), .B(KEYINPUT92), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n494), .B(new_n515), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT93), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XOR2_X1   g320(.A(new_n494), .B(KEYINPUT13), .Z(new_n522));
  OAI21_X1  g321(.A(KEYINPUT94), .B1(new_n507), .B2(new_n514), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(new_n515), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n521), .A2(KEYINPUT18), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT18), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n519), .A2(new_n520), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G113gat), .B(G141gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g331(.A(new_n532), .B(KEYINPUT12), .Z(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n525), .A2(new_n527), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n534), .B1(new_n525), .B2(new_n527), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n493), .A2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(G71gat), .A2(G78gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g341(.A(G57gat), .B(G64gat), .Z(new_n543));
  AOI21_X1  g342(.A(new_n542), .B1(new_n543), .B2(KEYINPUT95), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n543), .B1(KEYINPUT9), .B2(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI221_X1 g345(.A(new_n543), .B1(KEYINPUT9), .B2(new_n540), .C1(new_n542), .C2(KEYINPUT95), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT96), .B(KEYINPUT21), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(G231gat), .A2(G233gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n551), .B(new_n552), .ZN(new_n553));
  XNOR2_X1  g352(.A(new_n553), .B(G127gat), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n514), .B1(KEYINPUT21), .B2(new_n548), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n555), .B(KEYINPUT97), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n554), .B(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(G155gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(G183gat), .B(G211gat), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n559), .B(new_n560), .ZN(new_n561));
  XNOR2_X1  g360(.A(new_n557), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G85gat), .A2(G92gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(new_n563), .B(KEYINPUT7), .ZN(new_n564));
  INV_X1    g363(.A(G99gat), .ZN(new_n565));
  INV_X1    g364(.A(G106gat), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT8), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(KEYINPUT98), .B(G85gat), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n564), .B(new_n567), .C1(G92gat), .C2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(G99gat), .B(G106gat), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n569), .B(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT99), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n569), .B(new_n570), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AND2_X1   g375(.A1(new_n573), .A2(new_n576), .ZN(new_n577));
  OR2_X1    g376(.A1(new_n517), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n573), .A3(new_n507), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT100), .ZN(new_n580));
  NAND2_X1  g379(.A1(G232gat), .A2(G233gat), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT41), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n580), .B1(new_n579), .B2(new_n584), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n578), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G190gat), .B(G218gat), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n578), .B(new_n590), .C1(new_n585), .C2(new_n586), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  AOI21_X1  g391(.A(KEYINPUT101), .B1(new_n587), .B2(new_n588), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n581), .A2(new_n582), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(G134gat), .Z(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(G162gat), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n592), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n589), .A2(KEYINPUT101), .A3(new_n591), .A4(new_n596), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n562), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(G230gat), .ZN(new_n602));
  INV_X1    g401(.A(G233gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n572), .A2(new_n549), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n574), .A2(new_n548), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n576), .A2(new_n573), .A3(KEYINPUT10), .A4(new_n548), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n604), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NOR3_X1   g410(.A1(new_n607), .A2(new_n602), .A3(new_n603), .ZN(new_n612));
  OR2_X1    g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G176gat), .B(G204gat), .ZN(new_n615));
  XOR2_X1   g414(.A(new_n614), .B(new_n615), .Z(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT102), .ZN(new_n619));
  OR3_X1    g418(.A1(new_n611), .A2(new_n612), .A3(new_n617), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n613), .A2(KEYINPUT102), .A3(new_n617), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n601), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n539), .A2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n626), .A2(new_n445), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(new_n509), .ZN(G1324gat));
  INV_X1    g427(.A(KEYINPUT42), .ZN(new_n629));
  OAI21_X1  g428(.A(G8gat), .B1(new_n626), .B2(new_n446), .ZN(new_n630));
  XOR2_X1   g429(.A(KEYINPUT16), .B(G8gat), .Z(new_n631));
  NAND4_X1  g430(.A1(new_n539), .A2(new_n386), .A3(new_n625), .A4(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n629), .B1(new_n630), .B2(new_n632), .ZN(new_n633));
  AND2_X1   g432(.A1(new_n632), .A2(new_n629), .ZN(new_n634));
  NOR2_X1   g433(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT103), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n633), .A2(KEYINPUT103), .A3(new_n634), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(G1325gat));
  INV_X1    g438(.A(KEYINPUT104), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n492), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n491), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n642), .A2(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(KEYINPUT104), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n641), .A2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(G15gat), .B1(new_n626), .B2(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n642), .A2(G15gat), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n646), .B1(new_n626), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT105), .Z(G1326gat));
  NOR2_X1   g448(.A1(new_n626), .A2(new_n442), .ZN(new_n650));
  XOR2_X1   g449(.A(KEYINPUT43), .B(G22gat), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(G1327gat));
  INV_X1    g451(.A(new_n600), .ZN(new_n653));
  INV_X1    g452(.A(new_n562), .ZN(new_n654));
  AND4_X1   g453(.A1(new_n539), .A2(new_n623), .A3(new_n653), .A4(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n445), .A2(new_n497), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT45), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT44), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n659), .B1(new_n493), .B2(new_n600), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n467), .A2(new_n485), .ZN(new_n661));
  INV_X1    g460(.A(new_n447), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n492), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n360), .A2(new_n427), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT85), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n360), .A2(new_n427), .A3(KEYINPUT85), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n663), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n670), .A2(KEYINPUT44), .A3(new_n653), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n660), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n623), .B(KEYINPUT106), .ZN(new_n673));
  NOR3_X1   g472(.A1(new_n673), .A2(new_n538), .A3(new_n562), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n497), .B1(new_n675), .B2(new_n445), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n658), .A2(new_n676), .ZN(G1328gat));
  NOR2_X1   g476(.A1(new_n446), .A2(new_n498), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n655), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(new_n679), .B(KEYINPUT46), .Z(new_n680));
  OAI21_X1  g479(.A(new_n498), .B1(new_n675), .B2(new_n446), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  OAI21_X1  g481(.A(G43gat), .B1(new_n675), .B2(new_n492), .ZN(new_n683));
  INV_X1    g482(.A(G43gat), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n655), .A2(new_n684), .A3(new_n491), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n683), .A2(KEYINPUT47), .A3(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(G43gat), .B1(new_n675), .B2(new_n645), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n687), .A2(new_n685), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n686), .B1(new_n688), .B2(KEYINPUT47), .ZN(G1330gat));
  INV_X1    g488(.A(G50gat), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n655), .A2(new_n690), .A3(new_n253), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n660), .A2(new_n671), .A3(new_n253), .A4(new_n674), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(G50gat), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  OAI211_X1 g495(.A(KEYINPUT48), .B(new_n691), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n692), .A2(G50gat), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n691), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n697), .B1(KEYINPUT48), .B2(new_n699), .ZN(G1331gat));
  INV_X1    g499(.A(new_n673), .ZN(new_n701));
  INV_X1    g500(.A(new_n537), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n535), .ZN(new_n703));
  NOR3_X1   g502(.A1(new_n701), .A2(new_n703), .A3(new_n601), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n670), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  XNOR2_X1  g505(.A(new_n445), .B(KEYINPUT108), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g508(.A1(new_n705), .A2(new_n446), .ZN(new_n710));
  NOR2_X1   g509(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n711));
  AND2_X1   g510(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n710), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(new_n713), .B1(new_n710), .B2(new_n711), .ZN(G1333gat));
  NOR3_X1   g513(.A1(new_n705), .A2(G71gat), .A3(new_n642), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n641), .A2(new_n644), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n706), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n715), .B1(G71gat), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g518(.A1(new_n706), .A2(new_n253), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g520(.A1(new_n562), .A2(new_n703), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n670), .A2(KEYINPUT51), .A3(new_n653), .A4(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n670), .A2(new_n653), .A3(new_n722), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT51), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n430), .A2(new_n441), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n600), .B1(new_n729), .B2(new_n663), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n730), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n722), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n725), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n445), .A2(new_n568), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n732), .A2(new_n624), .A3(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n722), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n735), .A2(new_n623), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n672), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT109), .B1(new_n737), .B2(new_n445), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n568), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n737), .A2(KEYINPUT109), .A3(new_n445), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(G1336gat));
  NOR3_X1   g540(.A1(new_n701), .A2(G92gat), .A3(new_n446), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n732), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g542(.A1(new_n660), .A2(new_n671), .A3(new_n386), .A4(new_n736), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(G92gat), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT52), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(KEYINPUT113), .ZN(new_n747));
  OR2_X1    g546(.A1(new_n746), .A2(KEYINPUT113), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n743), .A2(new_n745), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT112), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n493), .A2(new_n600), .A3(new_n735), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n727), .B1(new_n751), .B2(KEYINPUT111), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT111), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n726), .A2(new_n753), .A3(KEYINPUT51), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n754), .A3(new_n742), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n745), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n750), .B1(new_n756), .B2(KEYINPUT52), .ZN(new_n757));
  AOI211_X1 g556(.A(KEYINPUT112), .B(new_n746), .C1(new_n755), .C2(new_n745), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n749), .B1(new_n757), .B2(new_n758), .ZN(G1337gat));
  OAI21_X1  g558(.A(G99gat), .B1(new_n737), .B2(new_n645), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n732), .A2(new_n565), .A3(new_n491), .A4(new_n624), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1338gat));
  INV_X1    g561(.A(KEYINPUT114), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n701), .A2(G106gat), .A3(new_n442), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n732), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n660), .A2(new_n671), .A3(new_n253), .A4(new_n736), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT53), .B1(new_n766), .B2(G106gat), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT53), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n752), .A2(new_n754), .A3(new_n764), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(G106gat), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n763), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n765), .A2(new_n767), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n770), .A2(new_n771), .ZN(new_n775));
  OAI211_X1 g574(.A(KEYINPUT114), .B(new_n774), .C1(new_n775), .C2(new_n769), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(G1339gat));
  NOR3_X1   g576(.A1(new_n601), .A2(new_n703), .A3(new_n624), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  AND4_X1   g578(.A1(KEYINPUT10), .A2(new_n573), .A3(new_n576), .A4(new_n548), .ZN(new_n780));
  AOI21_X1  g579(.A(KEYINPUT10), .B1(new_n606), .B2(new_n605), .ZN(new_n781));
  OAI22_X1  g580(.A1(new_n780), .A2(new_n781), .B1(new_n602), .B2(new_n603), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n609), .A2(new_n604), .A3(new_n610), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n782), .A2(KEYINPUT54), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT54), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n616), .B1(new_n611), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT55), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n784), .A2(new_n786), .A3(KEYINPUT55), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n789), .A2(new_n620), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(KEYINPUT115), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n789), .A2(new_n793), .A3(new_n620), .A4(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n517), .A2(new_n518), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n494), .B1(new_n796), .B2(new_n515), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n524), .A2(new_n522), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n532), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n598), .A2(new_n535), .A3(new_n599), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n795), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n535), .A2(new_n799), .ZN(new_n802));
  OR2_X1    g601(.A1(new_n802), .A2(new_n623), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n795), .B2(new_n538), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n801), .B1(new_n804), .B2(new_n600), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n779), .B1(new_n805), .B2(new_n562), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n707), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n437), .A2(new_n439), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n446), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n538), .A2(G113gat), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n703), .A2(new_n792), .A3(new_n794), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n653), .B1(new_n816), .B2(new_n803), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n654), .B1(new_n817), .B2(new_n801), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n253), .B1(new_n818), .B2(new_n779), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n468), .A2(new_n446), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n642), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n819), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(G113gat), .B1(new_n823), .B2(new_n538), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n815), .A2(new_n824), .ZN(G1340gat));
  NOR2_X1   g624(.A1(new_n623), .A2(new_n314), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n813), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n823), .B2(new_n701), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(KEYINPUT117), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(G1341gat));
  AND3_X1   g629(.A1(new_n822), .A2(G127gat), .A3(new_n562), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n811), .A2(new_n654), .ZN(new_n832));
  OR2_X1    g631(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  AOI21_X1  g632(.A(G127gat), .B1(new_n832), .B2(KEYINPUT118), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n831), .B1(new_n833), .B2(new_n834), .ZN(G1342gat));
  NAND2_X1  g634(.A1(new_n653), .A2(new_n446), .ZN(new_n836));
  XNOR2_X1  g635(.A(new_n836), .B(KEYINPUT119), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(G134gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n810), .A2(new_n838), .ZN(new_n839));
  OR2_X1    g638(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n840));
  OAI21_X1  g639(.A(G134gat), .B1(new_n823), .B2(new_n600), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(KEYINPUT56), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(G1343gat));
  AOI21_X1  g642(.A(new_n791), .B1(new_n702), .B2(new_n535), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n802), .A2(new_n623), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n600), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n800), .B2(new_n795), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n778), .B1(new_n847), .B2(new_n654), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT57), .B1(new_n848), .B2(new_n442), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n643), .A2(new_n820), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n806), .A2(new_n253), .ZN(new_n851));
  OAI211_X1 g650(.A(new_n849), .B(new_n850), .C1(new_n851), .C2(KEYINPUT57), .ZN(new_n852));
  OAI21_X1  g651(.A(G141gat), .B1(new_n852), .B2(new_n538), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n645), .A2(new_n253), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n807), .A2(new_n446), .A3(new_n855), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n538), .A2(G141gat), .ZN(new_n857));
  XNOR2_X1  g656(.A(new_n857), .B(KEYINPUT120), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n853), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  XNOR2_X1  g658(.A(new_n859), .B(KEYINPUT58), .ZN(G1344gat));
  NAND2_X1  g659(.A1(new_n851), .A2(KEYINPUT57), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT57), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n800), .A2(new_n791), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n562), .B1(new_n846), .B2(new_n863), .ZN(new_n864));
  OAI211_X1 g663(.A(new_n862), .B(new_n253), .C1(new_n864), .C2(new_n778), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n861), .A2(new_n624), .A3(new_n850), .A4(new_n865), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g667(.A(G148gat), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT59), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n220), .A2(KEYINPUT59), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n852), .B2(new_n623), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n856), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n874), .A2(new_n220), .A3(new_n624), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n873), .A2(new_n875), .ZN(G1345gat));
  OAI21_X1  g675(.A(G155gat), .B1(new_n852), .B2(new_n654), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n562), .A2(new_n216), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n877), .B1(new_n856), .B2(new_n878), .ZN(G1346gat));
  INV_X1    g678(.A(new_n215), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n880), .B1(new_n852), .B2(new_n600), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n837), .A2(new_n880), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n807), .A2(new_n855), .A3(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1347gat));
  NAND2_X1  g683(.A1(new_n445), .A2(new_n386), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n806), .A2(new_n886), .ZN(new_n887));
  NOR4_X1   g686(.A1(new_n887), .A2(G169gat), .A3(new_n538), .A4(new_n808), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT122), .Z(new_n889));
  OR2_X1    g688(.A1(new_n707), .A2(new_n446), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n642), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n819), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(G169gat), .B1(new_n892), .B2(new_n538), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n889), .A2(new_n893), .ZN(G1348gat));
  NOR2_X1   g693(.A1(new_n887), .A2(new_n808), .ZN(new_n895));
  INV_X1    g694(.A(G176gat), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n895), .A2(new_n896), .A3(new_n624), .ZN(new_n897));
  OAI21_X1  g696(.A(G176gat), .B1(new_n892), .B2(new_n701), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(G1349gat));
  NAND3_X1  g698(.A1(new_n895), .A2(new_n264), .A3(new_n562), .ZN(new_n900));
  OAI21_X1  g699(.A(G183gat), .B1(new_n892), .B2(new_n654), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g701(.A(new_n902), .B(KEYINPUT60), .ZN(G1350gat));
  INV_X1    g702(.A(KEYINPUT123), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n819), .A2(new_n653), .A3(new_n891), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G190gat), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n904), .A3(G190gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n907), .A2(KEYINPUT61), .A3(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n895), .A2(new_n265), .A3(new_n653), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n909), .B(new_n910), .C1(KEYINPUT61), .C2(new_n907), .ZN(G1351gat));
  AOI21_X1  g710(.A(new_n890), .B1(new_n644), .B2(new_n641), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n442), .B1(new_n818), .B2(new_n779), .ZN(new_n913));
  OAI211_X1 g712(.A(new_n865), .B(new_n912), .C1(new_n913), .C2(new_n862), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n914), .A2(new_n204), .A3(new_n538), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT124), .B1(new_n887), .B2(new_n854), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT124), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n885), .B1(new_n818), .B2(new_n779), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n855), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  AND2_X1   g718(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n920), .A2(new_n703), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n915), .B1(new_n921), .B2(new_n204), .ZN(G1352gat));
  NAND4_X1  g721(.A1(new_n855), .A2(new_n205), .A3(new_n918), .A4(new_n624), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT62), .Z(new_n924));
  OAI21_X1  g723(.A(G204gat), .B1(new_n914), .B2(new_n701), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n924), .A2(new_n925), .ZN(G1353gat));
  OAI21_X1  g725(.A(G211gat), .B1(new_n914), .B2(new_n654), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT63), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OAI211_X1 g728(.A(KEYINPUT63), .B(G211gat), .C1(new_n914), .C2(new_n654), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n654), .A2(G211gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n916), .A2(new_n919), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT125), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n916), .A2(new_n919), .A3(KEYINPUT125), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n931), .A2(new_n937), .A3(KEYINPUT126), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1354gat));
  AOI21_X1  g741(.A(G218gat), .B1(new_n920), .B2(new_n653), .ZN(new_n943));
  INV_X1    g742(.A(new_n914), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n653), .A2(G218gat), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT127), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n943), .B1(new_n944), .B2(new_n946), .ZN(G1355gat));
endmodule


