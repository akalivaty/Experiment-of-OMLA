//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:40 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n549, new_n550, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n569, new_n570, new_n571, new_n573, new_n574, new_n575, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT64), .B(G44), .Z(G218));
  XOR2_X1   g009(.A(KEYINPUT65), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  OR4_X1    g027(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n466), .B2(KEYINPUT69), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI211_X1 g044(.A(KEYINPUT69), .B(G125), .C1(new_n468), .C2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g046(.A(G2105), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(G101), .ZN(new_n474));
  AOI21_X1  g049(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  AND3_X1   g051(.A1(new_n472), .A2(new_n474), .A3(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n475), .A2(G136), .ZN(new_n478));
  INV_X1    g053(.A(new_n478), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  INV_X1    g055(.A(G112), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n480), .B1(new_n481), .B2(G2105), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT70), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n464), .A2(new_n465), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(new_n486));
  AOI211_X1 g061(.A(new_n479), .B(new_n483), .C1(G124), .C2(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n468), .C2(new_n469), .ZN(new_n488));
  OR2_X1    g063(.A1(G102), .A2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(G114), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G2105), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n489), .A2(new_n491), .A3(G2104), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n494), .C1(new_n468), .C2(new_n469), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n484), .A2(new_n497), .A3(G138), .A4(new_n494), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n496), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(KEYINPUT71), .A2(KEYINPUT5), .ZN(new_n500));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(KEYINPUT71), .A2(KEYINPUT5), .A3(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(G88), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT72), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n506), .A2(new_n510), .A3(new_n507), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n504), .A2(G62), .ZN(new_n512));
  INV_X1    g087(.A(G75), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n512), .B1(new_n513), .B2(new_n501), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n509), .A2(new_n511), .B1(G651), .B2(new_n514), .ZN(G166));
  XNOR2_X1  g090(.A(KEYINPUT73), .B(G89), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n504), .A2(new_n505), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n504), .A2(G63), .A3(G651), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n505), .A2(G51), .A3(G543), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n517), .A2(new_n518), .A3(new_n520), .A4(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(new_n503), .ZN(new_n527));
  AOI21_X1  g102(.A(G543), .B1(KEYINPUT71), .B2(KEYINPUT5), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  AND2_X1   g104(.A1(KEYINPUT6), .A2(G651), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n505), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n531), .A2(new_n532), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n526), .A2(new_n535), .ZN(G171));
  INV_X1    g111(.A(new_n531), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n505), .A2(G543), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n537), .A2(G81), .B1(new_n538), .B2(G43), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n504), .A2(G56), .ZN(new_n541));
  NAND2_X1  g116(.A1(G68), .A2(G543), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n525), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n539), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g119(.A1(new_n543), .A2(new_n540), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  NAND4_X1  g122(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT8), .ZN(new_n550));
  NAND4_X1  g125(.A1(G319), .A2(G483), .A3(G661), .A4(new_n550), .ZN(G188));
  AOI22_X1  g126(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n552));
  OR2_X1    g127(.A1(new_n552), .A2(new_n525), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n531), .A2(KEYINPUT76), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n504), .A2(new_n555), .A3(new_n505), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(new_n556), .A3(G91), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n505), .A2(G53), .A3(G543), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT75), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n538), .A2(new_n560), .A3(G53), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(KEYINPUT9), .ZN(new_n565));
  AND3_X1   g140(.A1(new_n564), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n558), .B1(new_n563), .B2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  NAND2_X1  g143(.A1(new_n514), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(new_n511), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n510), .B1(new_n506), .B2(new_n507), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(G303));
  OR2_X1    g147(.A1(new_n504), .A2(G74), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n538), .B2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n554), .A2(new_n556), .A3(G87), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G288));
  OAI21_X1  g151(.A(G61), .B1(new_n527), .B2(new_n528), .ZN(new_n577));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n579), .A2(G651), .B1(new_n538), .B2(G48), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n554), .A2(new_n556), .A3(G86), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(G305));
  AOI22_X1  g158(.A1(new_n537), .A2(G85), .B1(new_n538), .B2(G47), .ZN(new_n584));
  AOI22_X1  g159(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n525), .B2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n554), .A2(new_n556), .A3(G92), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  OR2_X1    g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n589), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G54), .ZN(new_n593));
  OAI22_X1  g168(.A1(new_n592), .A2(new_n525), .B1(new_n593), .B2(new_n533), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT77), .ZN(new_n595));
  INV_X1    g170(.A(KEYINPUT77), .ZN(new_n596));
  OAI221_X1 g171(.A(new_n596), .B1(new_n593), .B2(new_n533), .C1(new_n592), .C2(new_n525), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n590), .A2(new_n591), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n587), .B1(new_n598), .B2(G868), .ZN(G284));
  OAI21_X1  g174(.A(new_n587), .B1(new_n598), .B2(G868), .ZN(G321));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT78), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n553), .A2(new_n557), .ZN(new_n603));
  INV_X1    g178(.A(new_n566), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n564), .A2(new_n565), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n605), .A2(KEYINPUT75), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n603), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n602), .B1(new_n607), .B2(G868), .ZN(G297));
  OAI21_X1  g183(.A(new_n602), .B1(new_n607), .B2(G868), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n598), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n598), .A2(new_n610), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(G868), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n486), .A2(G123), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT80), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n475), .A2(G135), .ZN(new_n618));
  NOR2_X1   g193(.A1(new_n494), .A2(G111), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  OAI211_X1 g195(.A(new_n617), .B(new_n618), .C1(new_n619), .C2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT81), .B(G2096), .Z(new_n622));
  OR2_X1    g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  XOR2_X1   g199(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n625));
  NOR3_X1   g200(.A1(new_n462), .A2(new_n463), .A3(G2105), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT13), .B(G2100), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n623), .A2(new_n624), .A3(new_n629), .ZN(G156));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2435), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT82), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(G2427), .B(G2430), .Z(new_n634));
  OR2_X1    g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n634), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n635), .A2(KEYINPUT14), .A3(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G1341), .B(G1348), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT83), .ZN(new_n645));
  OAI21_X1  g220(.A(G14), .B1(new_n642), .B2(new_n643), .ZN(new_n646));
  NOR2_X1   g221(.A1(new_n645), .A2(new_n646), .ZN(G401));
  INV_X1    g222(.A(KEYINPUT18), .ZN(new_n648));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT17), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n649), .A2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n648), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2100), .ZN(new_n655));
  XOR2_X1   g230(.A(G2072), .B(G2078), .Z(new_n656));
  AOI21_X1  g231(.A(new_n656), .B1(new_n651), .B2(KEYINPUT18), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n655), .B(new_n658), .ZN(G227));
  XOR2_X1   g234(.A(G1971), .B(G1976), .Z(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(G1956), .B(G2474), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT20), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n663), .A2(new_n664), .ZN(new_n668));
  NOR3_X1   g243(.A1(new_n661), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n669), .B1(new_n661), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  XNOR2_X1  g248(.A(G1991), .B(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G229));
  MUX2_X1   g253(.A(G23), .B(G288), .S(G16), .Z(new_n679));
  XOR2_X1   g254(.A(KEYINPUT33), .B(G1976), .Z(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G6), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n582), .B2(new_n682), .ZN(new_n684));
  XOR2_X1   g259(.A(KEYINPUT32), .B(G1981), .Z(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(G22), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT86), .Z(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(G166), .B2(new_n682), .ZN(new_n689));
  OAI21_X1  g264(.A(new_n686), .B1(G1971), .B2(new_n689), .ZN(new_n690));
  AOI211_X1 g265(.A(new_n681), .B(new_n690), .C1(G1971), .C2(new_n689), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT34), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  MUX2_X1   g269(.A(G24), .B(G290), .S(G16), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n697));
  AND2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n696), .A2(new_n697), .ZN(new_n699));
  NOR2_X1   g274(.A1(G25), .A2(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n486), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n475), .A2(G131), .ZN(new_n702));
  OR2_X1    g277(.A1(G95), .A2(G2105), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n703), .B(G2104), .C1(G107), .C2(new_n494), .ZN(new_n704));
  NAND3_X1  g279(.A1(new_n701), .A2(new_n702), .A3(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n700), .B1(new_n706), .B2(G29), .ZN(new_n707));
  XOR2_X1   g282(.A(KEYINPUT35), .B(G1991), .Z(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT84), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NOR3_X1   g285(.A1(new_n698), .A2(new_n699), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n693), .A2(new_n694), .A3(new_n711), .ZN(new_n712));
  XOR2_X1   g287(.A(new_n712), .B(KEYINPUT36), .Z(new_n713));
  INV_X1    g288(.A(G29), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n714), .A2(G33), .ZN(new_n715));
  XNOR2_X1  g290(.A(KEYINPUT88), .B(KEYINPUT25), .ZN(new_n716));
  AND3_X1   g291(.A1(new_n494), .A2(G103), .A3(G2104), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n475), .A2(G139), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n484), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n718), .B(new_n719), .C1(new_n494), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n715), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2072), .ZN(new_n725));
  NOR2_X1   g300(.A1(G286), .A2(new_n682), .ZN(new_n726));
  INV_X1    g301(.A(KEYINPUT92), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G16), .B2(G21), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n726), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n729), .B1(KEYINPUT92), .B2(new_n726), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT93), .B(G1966), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n724), .A2(new_n725), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n730), .A2(new_n731), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n732), .B(new_n733), .C1(new_n725), .C2(new_n724), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n682), .A2(G5), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(G171), .B2(new_n682), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(G1961), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n714), .A2(G27), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G164), .B2(new_n714), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n739), .B(G2078), .ZN(new_n740));
  NOR2_X1   g315(.A1(G29), .A2(G32), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(KEYINPUT91), .ZN(new_n742));
  NAND3_X1  g317(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n743));
  XOR2_X1   g318(.A(new_n743), .B(KEYINPUT26), .Z(new_n744));
  INV_X1    g319(.A(G129), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n485), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n475), .A2(G141), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n473), .A2(G105), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT90), .Z(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(new_n714), .ZN(new_n752));
  MUX2_X1   g327(.A(new_n742), .B(KEYINPUT91), .S(new_n752), .Z(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT27), .B(G1996), .ZN(new_n754));
  INV_X1    g329(.A(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n737), .B(new_n740), .C1(new_n753), .C2(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n682), .A2(G4), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(new_n598), .B2(new_n682), .ZN(new_n758));
  INV_X1    g333(.A(G1348), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n756), .B(new_n760), .C1(new_n755), .C2(new_n753), .ZN(new_n761));
  NAND2_X1  g336(.A1(G162), .A2(G29), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G29), .B2(G35), .ZN(new_n763));
  XOR2_X1   g338(.A(KEYINPUT29), .B(G2090), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n621), .A2(new_n714), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n765), .B1(KEYINPUT94), .B2(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n767), .B1(KEYINPUT94), .B2(new_n766), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n770), .A2(G28), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n714), .B1(new_n770), .B2(G28), .ZN(new_n772));
  OAI221_X1 g347(.A(new_n769), .B1(new_n771), .B2(new_n772), .C1(new_n763), .C2(new_n764), .ZN(new_n773));
  XNOR2_X1  g348(.A(KEYINPUT87), .B(KEYINPUT28), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n714), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n475), .A2(G140), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n494), .A2(G116), .ZN(new_n778));
  OAI21_X1  g353(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n779));
  INV_X1    g354(.A(G128), .ZN(new_n780));
  OAI221_X1 g355(.A(new_n777), .B1(new_n778), .B2(new_n779), .C1(new_n780), .C2(new_n485), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n776), .B1(new_n781), .B2(G29), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n773), .A2(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT24), .ZN(new_n786));
  INV_X1    g361(.A(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(G29), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n788), .B1(new_n786), .B2(new_n787), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G160), .B2(new_n714), .ZN(new_n790));
  INV_X1    g365(.A(G2084), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n768), .A2(new_n785), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n682), .A2(G20), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT23), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n607), .B2(new_n682), .ZN(new_n796));
  INV_X1    g371(.A(G1956), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n796), .B(new_n797), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n682), .A2(G19), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n546), .B2(new_n682), .ZN(new_n800));
  XOR2_X1   g375(.A(new_n800), .B(G1341), .Z(new_n801));
  NAND2_X1  g376(.A1(new_n798), .A2(new_n801), .ZN(new_n802));
  OR4_X1    g377(.A1(new_n734), .A2(new_n761), .A3(new_n793), .A4(new_n802), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n713), .A2(new_n803), .ZN(G311));
  OR2_X1    g379(.A1(new_n713), .A2(new_n803), .ZN(G150));
  AOI22_X1  g380(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(new_n525), .ZN(new_n807));
  INV_X1    g382(.A(G93), .ZN(new_n808));
  INV_X1    g383(.A(G55), .ZN(new_n809));
  OAI22_X1  g384(.A1(new_n531), .A2(new_n808), .B1(new_n533), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n807), .A2(new_n810), .ZN(new_n811));
  INV_X1    g386(.A(G860), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT37), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n598), .A2(G559), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT95), .Z(new_n816));
  INV_X1    g391(.A(KEYINPUT38), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n546), .A2(new_n811), .ZN(new_n819));
  OAI22_X1  g394(.A1(new_n544), .A2(new_n545), .B1(new_n807), .B2(new_n810), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n818), .B(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  OR2_X1    g398(.A1(new_n818), .A2(new_n821), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n818), .A2(new_n821), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n823), .A2(new_n827), .A3(new_n812), .ZN(new_n828));
  AND2_X1   g403(.A1(new_n828), .A2(KEYINPUT96), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(KEYINPUT96), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n814), .B1(new_n829), .B2(new_n830), .ZN(G145));
  MUX2_X1   g406(.A(new_n751), .B(new_n750), .S(new_n723), .Z(new_n832));
  NAND2_X1  g407(.A1(G126), .A2(G2105), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n464), .B2(new_n465), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n494), .A2(G114), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g412(.A(KEYINPUT97), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT97), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n488), .A2(new_n839), .A3(new_n492), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n497), .B1(new_n475), .B2(G138), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n842));
  OAI211_X1 g417(.A(new_n838), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(new_n781), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n832), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n475), .A2(G142), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n846), .B(KEYINPUT98), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n486), .A2(G130), .ZN(new_n848));
  NOR2_X1   g423(.A1(new_n494), .A2(G118), .ZN(new_n849));
  OAI21_X1  g424(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n847), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n706), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n627), .ZN(new_n853));
  OR2_X1    g428(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n845), .A2(new_n853), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n854), .A2(KEYINPUT99), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(G162), .B(G160), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(new_n621), .ZN(new_n858));
  AOI21_X1  g433(.A(G37), .B1(new_n856), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n858), .B2(new_n856), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g436(.A(new_n821), .B(new_n612), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n863), .B1(new_n598), .B2(G299), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n590), .A2(new_n591), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n595), .A2(new_n597), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n867), .A2(new_n607), .A3(KEYINPUT100), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n598), .A2(G299), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n862), .A2(new_n870), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT101), .Z(new_n872));
  INV_X1    g447(.A(KEYINPUT41), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g449(.A1(new_n864), .A2(new_n868), .A3(KEYINPUT41), .A4(new_n869), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(KEYINPUT102), .A3(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n862), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT102), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n870), .A2(new_n878), .A3(new_n873), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n582), .B(G288), .ZN(new_n881));
  XNOR2_X1  g456(.A(G303), .B(G290), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n881), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n872), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n872), .B2(new_n880), .ZN(new_n888));
  OAI21_X1  g463(.A(G868), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n811), .A2(G868), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(G295));
  INV_X1    g467(.A(G868), .ZN(new_n893));
  INV_X1    g468(.A(new_n888), .ZN(new_n894));
  AOI21_X1  g469(.A(new_n893), .B1(new_n894), .B2(new_n886), .ZN(new_n895));
  OAI21_X1  g470(.A(KEYINPUT103), .B1(new_n895), .B2(new_n890), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT103), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n889), .A2(new_n897), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(G331));
  AOI21_X1  g474(.A(G286), .B1(G171), .B2(KEYINPUT104), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(G171), .A2(KEYINPUT104), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n819), .A2(new_n820), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n903), .B1(new_n819), .B2(new_n820), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n901), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(new_n906), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n908), .A2(new_n900), .A3(new_n904), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n876), .A2(new_n910), .A3(new_n879), .ZN(new_n911));
  INV_X1    g486(.A(new_n883), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n907), .A2(new_n909), .A3(new_n870), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  AOI21_X1  g490(.A(G37), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n911), .A2(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(new_n883), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n911), .A2(KEYINPUT105), .A3(new_n912), .A4(new_n913), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n916), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT43), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT106), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n910), .B1(new_n923), .B2(new_n875), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n874), .A2(new_n923), .A3(new_n875), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n913), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(new_n883), .ZN(new_n927));
  AND4_X1   g502(.A1(KEYINPUT43), .A2(new_n916), .A3(new_n919), .A4(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(KEYINPUT44), .B1(new_n922), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n920), .A2(KEYINPUT43), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n916), .A2(new_n921), .A3(new_n927), .A4(new_n919), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  NAND3_X1  g510(.A1(new_n476), .A2(G40), .A3(new_n474), .ZN(new_n936));
  OAI21_X1  g511(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT69), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n939), .A2(new_n470), .A3(new_n460), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n936), .B1(new_n940), .B2(G2105), .ZN(new_n941));
  INV_X1    g516(.A(G1384), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT50), .B1(new_n843), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT50), .ZN(new_n944));
  NOR3_X1   g519(.A1(G164), .A2(new_n944), .A3(G1384), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n941), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G1961), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(KEYINPUT45), .B1(new_n843), .B2(new_n942), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n476), .A2(G40), .A3(new_n474), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n942), .A2(KEYINPUT45), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n472), .B(new_n950), .C1(G164), .C2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G2078), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT53), .ZN(new_n954));
  OR3_X1    g529(.A1(new_n949), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(KEYINPUT107), .B(G1384), .Z(new_n956));
  NAND3_X1  g531(.A1(new_n843), .A2(KEYINPUT45), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n958), .B1(G164), .B2(G1384), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n957), .A2(new_n959), .A3(new_n953), .A4(new_n941), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT53), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n948), .A2(new_n955), .A3(new_n962), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n963), .A2(G171), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n843), .A2(new_n956), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n954), .B1(new_n965), .B2(new_n958), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n966), .A2(new_n941), .A3(new_n957), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n948), .A2(new_n962), .A3(new_n967), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n968), .A2(KEYINPUT122), .A3(G171), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT122), .B1(new_n968), .B2(G171), .ZN(new_n970));
  OAI211_X1 g545(.A(KEYINPUT54), .B(new_n964), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT55), .ZN(new_n972));
  INV_X1    g547(.A(G8), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n972), .B1(G166), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT109), .ZN(new_n975));
  NAND4_X1  g550(.A1(G303), .A2(new_n975), .A3(KEYINPUT55), .A4(G8), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n509), .A2(new_n511), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n973), .B1(new_n978), .B2(new_n569), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n975), .B1(new_n979), .B2(KEYINPUT55), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n977), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n493), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n841), .B2(new_n842), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n983), .A2(new_n944), .A3(new_n942), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(new_n941), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n944), .B1(new_n843), .B2(new_n942), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(G2090), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n957), .A2(new_n941), .A3(new_n959), .ZN(new_n989));
  INV_X1    g564(.A(G1971), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n987), .A2(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n981), .B1(new_n991), .B2(new_n973), .ZN(new_n992));
  INV_X1    g567(.A(G1981), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n580), .A2(new_n581), .A3(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n580), .A2(new_n581), .A3(KEYINPUT111), .A4(new_n993), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(G86), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n580), .B1(new_n999), .B2(new_n531), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(G1981), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n998), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT49), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n998), .A2(KEYINPUT49), .A3(new_n1001), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n941), .A2(new_n942), .A3(new_n843), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(G8), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1004), .A2(new_n1005), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n989), .A2(new_n990), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1010), .B1(G2090), .B2(new_n946), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT109), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(new_n974), .A3(new_n976), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1014), .A3(G8), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n574), .A2(new_n575), .A3(G1976), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1006), .A2(G8), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT52), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(new_n1020), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(KEYINPUT52), .A2(G1976), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1017), .A2(new_n1021), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1022), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n992), .A2(new_n1009), .A3(new_n1015), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n963), .A2(G171), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n948), .A2(new_n967), .A3(new_n962), .A4(G301), .ZN(new_n1028));
  AOI21_X1  g603(.A(KEYINPUT54), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1026), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1966), .ZN(new_n1031));
  OAI21_X1  g606(.A(new_n1031), .B1(new_n949), .B2(new_n952), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n472), .A2(new_n791), .A3(new_n950), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n943), .B2(new_n945), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(G8), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n1037));
  NAND3_X1  g612(.A1(G286), .A2(new_n1037), .A3(G8), .ZN(new_n1038));
  INV_X1    g613(.A(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1037), .B1(G286), .B2(G8), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  NOR2_X1   g619(.A1(KEYINPUT120), .A2(KEYINPUT51), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1036), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(new_n1045), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n973), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n1043), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1046), .A2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1041), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1051));
  XNOR2_X1  g626(.A(new_n1051), .B(KEYINPUT119), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n1053));
  AND3_X1   g628(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1053), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n971), .B(new_n1030), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT116), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n797), .B1(new_n985), .B2(new_n986), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n957), .A2(new_n959), .A3(new_n941), .A4(new_n1060), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1059), .B1(new_n1058), .B2(new_n1061), .ZN(new_n1063));
  NOR3_X1   g638(.A1(new_n603), .A2(KEYINPUT57), .A3(new_n561), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(G299), .B2(KEYINPUT57), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n1062), .A2(new_n1063), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1065), .A2(new_n1058), .A3(new_n1061), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT61), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1057), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1065), .B1(new_n1070), .B2(KEYINPUT113), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(KEYINPUT116), .A3(KEYINPUT61), .A4(new_n1067), .ZN(new_n1074));
  AND4_X1   g649(.A1(new_n942), .A2(new_n843), .A3(new_n472), .A4(new_n950), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT58), .B(G1341), .ZN(new_n1076));
  OAI22_X1  g651(.A1(new_n989), .A2(G1996), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n546), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1078), .A2(KEYINPUT115), .A3(KEYINPUT59), .ZN(new_n1079));
  NAND2_X1  g654(.A1(KEYINPUT115), .A2(KEYINPUT59), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n546), .A3(new_n1080), .ZN(new_n1081));
  AOI22_X1  g656(.A1(new_n946), .A2(new_n759), .B1(new_n783), .B2(new_n1075), .ZN(new_n1082));
  OR2_X1    g657(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n867), .B1(new_n1082), .B2(KEYINPUT60), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n1079), .A2(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1064), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1086), .B1(new_n607), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1070), .A2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1067), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT61), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1082), .A2(KEYINPUT60), .ZN(new_n1092));
  AOI22_X1  g667(.A1(new_n1090), .A2(new_n1091), .B1(new_n1092), .B2(new_n867), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1069), .A2(new_n1074), .A3(new_n1085), .A4(new_n1093), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1082), .A2(new_n867), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1095), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1067), .ZN(new_n1097));
  OAI21_X1  g672(.A(KEYINPUT114), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT114), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1099), .B(new_n1067), .C1(new_n1066), .C2(new_n1095), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1094), .A2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1056), .B1(new_n1102), .B2(KEYINPUT117), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT117), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1094), .A2(new_n1101), .A3(new_n1104), .ZN(new_n1105));
  NOR2_X1   g680(.A1(G288), .A2(G1976), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1009), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n998), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1015), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1007), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1110));
  AOI22_X1  g685(.A1(new_n1110), .A2(new_n1005), .B1(new_n1022), .B2(new_n1024), .ZN(new_n1111));
  AOI22_X1  g686(.A1(new_n1108), .A2(new_n1008), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1014), .B1(new_n1011), .B2(G8), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT63), .ZN(new_n1114));
  NOR4_X1   g689(.A1(new_n1113), .A2(new_n1114), .A3(G286), .A4(new_n1036), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1009), .A2(new_n1025), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1109), .ZN(new_n1117));
  AND2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1036), .A2(G286), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1111), .A2(new_n992), .A3(new_n1015), .A4(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1120), .A2(new_n1114), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT112), .B(new_n1112), .C1(new_n1118), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT112), .ZN(new_n1123));
  AOI22_X1  g698(.A1(new_n1117), .A2(new_n1115), .B1(new_n1120), .B2(new_n1114), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1107), .A2(new_n998), .ZN(new_n1125));
  OAI22_X1  g700(.A1(new_n1125), .A2(new_n1007), .B1(new_n1116), .B2(new_n1015), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1123), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1127));
  AOI22_X1  g702(.A1(new_n1103), .A2(new_n1105), .B1(new_n1122), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT124), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1045), .B1(new_n1036), .B2(new_n1044), .ZN(new_n1130));
  NOR3_X1   g705(.A1(new_n1048), .A2(new_n1043), .A3(new_n1047), .ZN(new_n1131));
  NOR2_X1   g706(.A1(new_n1051), .A2(KEYINPUT119), .ZN(new_n1132));
  OR2_X1    g707(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1035), .A2(KEYINPUT119), .A3(new_n1133), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1130), .A2(new_n1131), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1135), .A2(KEYINPUT121), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT62), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1050), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1136), .A2(new_n1137), .A3(new_n1138), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1139), .A2(KEYINPUT123), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT62), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(KEYINPUT123), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1129), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT123), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1148), .A2(KEYINPUT124), .A3(new_n1142), .A4(new_n1141), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1128), .A2(new_n1145), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n965), .A2(new_n958), .ZN(new_n1151));
  INV_X1    g726(.A(new_n941), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n781), .B(new_n783), .ZN(new_n1154));
  OAI21_X1  g729(.A(G1996), .B1(new_n746), .B2(new_n749), .ZN(new_n1155));
  OAI211_X1 g730(.A(new_n1154), .B(new_n1155), .C1(new_n751), .C2(G1996), .ZN(new_n1156));
  XNOR2_X1  g731(.A(new_n705), .B(new_n708), .ZN(new_n1157));
  XNOR2_X1  g732(.A(new_n1157), .B(KEYINPUT108), .ZN(new_n1158));
  OR2_X1    g733(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g734(.A(G290), .B(G1986), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1153), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1150), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1153), .ZN(new_n1163));
  OR3_X1    g738(.A1(new_n1163), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1164));
  OAI21_X1  g739(.A(KEYINPUT46), .B1(new_n1163), .B2(G1996), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1154), .A2(new_n750), .ZN(new_n1166));
  AOI22_X1  g741(.A1(new_n1164), .A2(new_n1165), .B1(new_n1153), .B2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT47), .Z(new_n1168));
  NAND2_X1  g743(.A1(new_n706), .A2(new_n708), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1156), .A2(new_n1169), .ZN(new_n1170));
  OR2_X1    g745(.A1(new_n781), .A2(G2067), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1163), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  OR3_X1    g747(.A1(new_n1163), .A2(G1986), .A3(G290), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT125), .B(KEYINPUT48), .ZN(new_n1174));
  AOI22_X1  g749(.A1(new_n1159), .A2(new_n1153), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  OR2_X1    g750(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n1172), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  XOR2_X1   g753(.A(new_n1178), .B(KEYINPUT126), .Z(new_n1179));
  NAND2_X1  g754(.A1(new_n1162), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g755(.A1(G227), .A2(new_n458), .ZN(new_n1182));
  XNOR2_X1  g756(.A(new_n1182), .B(KEYINPUT127), .ZN(new_n1183));
  NOR3_X1   g757(.A1(G229), .A2(G401), .A3(new_n1183), .ZN(new_n1184));
  NAND3_X1  g758(.A1(new_n932), .A2(new_n860), .A3(new_n1184), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


