

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594;

  XNOR2_X1 U325 ( .A(n450), .B(KEYINPUT114), .ZN(n451) );
  XNOR2_X1 U326 ( .A(n452), .B(n451), .ZN(n453) );
  NOR2_X1 U327 ( .A1(n537), .A2(n456), .ZN(n457) );
  INV_X1 U328 ( .A(G169GAT), .ZN(n462) );
  XNOR2_X1 U329 ( .A(n368), .B(n367), .ZN(n561) );
  XNOR2_X1 U330 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U331 ( .A(n461), .B(n460), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n294) );
  XNOR2_X1 U333 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n293) );
  XNOR2_X1 U334 ( .A(n294), .B(n293), .ZN(n445) );
  XOR2_X1 U335 ( .A(KEYINPUT0), .B(G127GAT), .Z(n332) );
  XOR2_X1 U336 ( .A(n445), .B(n332), .Z(n296) );
  NAND2_X1 U337 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U339 ( .A(KEYINPUT81), .B(KEYINPUT20), .Z(n298) );
  XNOR2_X1 U340 ( .A(G15GAT), .B(G183GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U342 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U343 ( .A(G190GAT), .B(G99GAT), .Z(n302) );
  XNOR2_X1 U344 ( .A(G43GAT), .B(G134GAT), .ZN(n301) );
  XNOR2_X1 U345 ( .A(n302), .B(n301), .ZN(n306) );
  XOR2_X1 U346 ( .A(G176GAT), .B(G71GAT), .Z(n304) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G120GAT), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U350 ( .A(n308), .B(n307), .ZN(n537) );
  XOR2_X1 U351 ( .A(KEYINPUT22), .B(KEYINPUT84), .Z(n310) );
  XNOR2_X1 U352 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n322) );
  XOR2_X1 U354 ( .A(G50GAT), .B(KEYINPUT73), .Z(n347) );
  XOR2_X1 U355 ( .A(n347), .B(G204GAT), .Z(n312) );
  XOR2_X1 U356 ( .A(G106GAT), .B(G78GAT), .Z(n413) );
  XNOR2_X1 U357 ( .A(G148GAT), .B(n413), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(n313), .B(KEYINPUT83), .Z(n320) );
  XOR2_X1 U360 ( .A(KEYINPUT21), .B(G211GAT), .Z(n315) );
  XNOR2_X1 U361 ( .A(G197GAT), .B(G218GAT), .ZN(n314) );
  XNOR2_X1 U362 ( .A(n315), .B(n314), .ZN(n449) );
  XOR2_X1 U363 ( .A(n449), .B(KEYINPUT82), .Z(n317) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XNOR2_X1 U366 ( .A(G22GAT), .B(n318), .ZN(n319) );
  XNOR2_X1 U367 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U368 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U369 ( .A(KEYINPUT3), .B(G162GAT), .Z(n324) );
  XNOR2_X1 U370 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n323) );
  XNOR2_X1 U371 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U372 ( .A(G141GAT), .B(n325), .Z(n342) );
  XOR2_X1 U373 ( .A(n326), .B(n342), .Z(n473) );
  XNOR2_X1 U374 ( .A(G120GAT), .B(G57GAT), .ZN(n327) );
  XNOR2_X1 U375 ( .A(n327), .B(G148GAT), .ZN(n408) );
  XNOR2_X1 U376 ( .A(G29GAT), .B(G134GAT), .ZN(n328) );
  XNOR2_X1 U377 ( .A(n328), .B(KEYINPUT76), .ZN(n349) );
  XOR2_X1 U378 ( .A(KEYINPUT88), .B(n349), .Z(n330) );
  NAND2_X1 U379 ( .A1(G225GAT), .A2(G233GAT), .ZN(n329) );
  XNOR2_X1 U380 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U381 ( .A(n408), .B(n331), .Z(n334) );
  XOR2_X1 U382 ( .A(G113GAT), .B(G1GAT), .Z(n401) );
  XNOR2_X1 U383 ( .A(n401), .B(n332), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U385 ( .A(KEYINPUT5), .B(KEYINPUT86), .Z(n336) );
  XNOR2_X1 U386 ( .A(G85GAT), .B(KEYINPUT1), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U388 ( .A(n338), .B(n337), .Z(n344) );
  XOR2_X1 U389 ( .A(KEYINPUT87), .B(KEYINPUT6), .Z(n340) );
  XNOR2_X1 U390 ( .A(KEYINPUT4), .B(KEYINPUT85), .ZN(n339) );
  XNOR2_X1 U391 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U392 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U393 ( .A(n344), .B(n343), .Z(n471) );
  XNOR2_X1 U394 ( .A(KEYINPUT89), .B(n471), .ZN(n475) );
  INV_X1 U395 ( .A(n475), .ZN(n521) );
  INV_X1 U396 ( .A(KEYINPUT36), .ZN(n369) );
  XOR2_X1 U397 ( .A(KEYINPUT9), .B(KEYINPUT74), .Z(n346) );
  XNOR2_X1 U398 ( .A(G218GAT), .B(KEYINPUT10), .ZN(n345) );
  XNOR2_X1 U399 ( .A(n346), .B(n345), .ZN(n348) );
  XOR2_X1 U400 ( .A(n348), .B(n347), .Z(n355) );
  INV_X1 U401 ( .A(G106GAT), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n350), .B(n349), .ZN(n353) );
  XOR2_X1 U403 ( .A(G99GAT), .B(G85GAT), .Z(n414) );
  NAND2_X1 U404 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U405 ( .A(n414), .B(n351), .ZN(n352) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n354) );
  NAND2_X1 U407 ( .A1(n355), .A2(n354), .ZN(n359) );
  INV_X1 U408 ( .A(n354), .ZN(n357) );
  INV_X1 U409 ( .A(n355), .ZN(n356) );
  NAND2_X1 U410 ( .A1(n357), .A2(n356), .ZN(n358) );
  NAND2_X1 U411 ( .A1(n359), .A2(n358), .ZN(n363) );
  XOR2_X1 U412 ( .A(KEYINPUT75), .B(KEYINPUT11), .Z(n361) );
  XNOR2_X1 U413 ( .A(G162GAT), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U414 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n368) );
  XOR2_X1 U416 ( .A(G43GAT), .B(KEYINPUT8), .Z(n365) );
  XNOR2_X1 U417 ( .A(KEYINPUT7), .B(KEYINPUT67), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n402) );
  XNOR2_X1 U419 ( .A(G36GAT), .B(G190GAT), .ZN(n366) );
  XNOR2_X1 U420 ( .A(n366), .B(KEYINPUT77), .ZN(n437) );
  XOR2_X1 U421 ( .A(n402), .B(n437), .Z(n367) );
  XNOR2_X1 U422 ( .A(n369), .B(n561), .ZN(n490) );
  XOR2_X1 U423 ( .A(G8GAT), .B(G183GAT), .Z(n440) );
  XOR2_X1 U424 ( .A(G71GAT), .B(KEYINPUT13), .Z(n419) );
  XOR2_X1 U425 ( .A(n440), .B(n419), .Z(n371) );
  XNOR2_X1 U426 ( .A(G155GAT), .B(G57GAT), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U428 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n373) );
  NAND2_X1 U429 ( .A1(G231GAT), .A2(G233GAT), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U431 ( .A(n375), .B(n374), .Z(n377) );
  XOR2_X1 U432 ( .A(G22GAT), .B(G15GAT), .Z(n399) );
  XNOR2_X1 U433 ( .A(n399), .B(KEYINPUT14), .ZN(n376) );
  XNOR2_X1 U434 ( .A(n377), .B(n376), .ZN(n385) );
  XOR2_X1 U435 ( .A(G64GAT), .B(G78GAT), .Z(n379) );
  XNOR2_X1 U436 ( .A(G1GAT), .B(G127GAT), .ZN(n378) );
  XNOR2_X1 U437 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U438 ( .A(G211GAT), .B(KEYINPUT80), .Z(n381) );
  XNOR2_X1 U439 ( .A(KEYINPUT79), .B(KEYINPUT78), .ZN(n380) );
  XNOR2_X1 U440 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U441 ( .A(n383), .B(n382), .Z(n384) );
  XNOR2_X1 U442 ( .A(n385), .B(n384), .ZN(n545) );
  NOR2_X1 U443 ( .A1(n490), .A2(n545), .ZN(n387) );
  INV_X1 U444 ( .A(KEYINPUT45), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n405) );
  XOR2_X1 U446 ( .A(G197GAT), .B(KEYINPUT29), .Z(n389) );
  NAND2_X1 U447 ( .A1(G229GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n393) );
  XOR2_X1 U449 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n391) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(KEYINPUT66), .ZN(n390) );
  XNOR2_X1 U451 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U452 ( .A(n393), .B(n392), .Z(n398) );
  XOR2_X1 U453 ( .A(G141GAT), .B(G36GAT), .Z(n395) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(G50GAT), .ZN(n394) );
  XNOR2_X1 U455 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U456 ( .A(G169GAT), .B(n396), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U458 ( .A(n400), .B(n399), .Z(n404) );
  XNOR2_X1 U459 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n577) );
  NOR2_X1 U461 ( .A1(n405), .A2(n577), .ZN(n424) );
  XOR2_X1 U462 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT70), .B(KEYINPUT69), .ZN(n406) );
  XNOR2_X1 U464 ( .A(n407), .B(n406), .ZN(n412) );
  XOR2_X1 U465 ( .A(n408), .B(KEYINPUT72), .Z(n410) );
  NAND2_X1 U466 ( .A1(G230GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U467 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n423) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n417) );
  XOR2_X1 U470 ( .A(G64GAT), .B(G204GAT), .Z(n416) );
  XNOR2_X1 U471 ( .A(G176GAT), .B(G92GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n444) );
  XNOR2_X1 U473 ( .A(n417), .B(n444), .ZN(n418) );
  XOR2_X1 U474 ( .A(n418), .B(KEYINPUT33), .Z(n421) );
  XNOR2_X1 U475 ( .A(n419), .B(KEYINPUT71), .ZN(n420) );
  XNOR2_X1 U476 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U477 ( .A(n423), .B(n422), .ZN(n582) );
  NAND2_X1 U478 ( .A1(n424), .A2(n582), .ZN(n431) );
  XNOR2_X1 U479 ( .A(n582), .B(KEYINPUT41), .ZN(n555) );
  NAND2_X1 U480 ( .A1(n577), .A2(n555), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n425), .B(KEYINPUT46), .ZN(n426) );
  NAND2_X1 U482 ( .A1(n426), .A2(n545), .ZN(n427) );
  NOR2_X1 U483 ( .A1(n561), .A2(n427), .ZN(n428) );
  XNOR2_X1 U484 ( .A(n428), .B(KEYINPUT47), .ZN(n432) );
  AND2_X1 U485 ( .A1(n431), .A2(n432), .ZN(n430) );
  XNOR2_X1 U486 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n433) );
  INV_X1 U487 ( .A(n433), .ZN(n429) );
  NAND2_X1 U488 ( .A1(n430), .A2(n429), .ZN(n436) );
  NAND2_X1 U489 ( .A1(n432), .A2(n431), .ZN(n434) );
  NAND2_X1 U490 ( .A1(n434), .A2(n433), .ZN(n435) );
  NAND2_X1 U491 ( .A1(n436), .A2(n435), .ZN(n534) );
  XOR2_X1 U492 ( .A(n437), .B(KEYINPUT92), .Z(n439) );
  NAND2_X1 U493 ( .A1(G226GAT), .A2(G233GAT), .ZN(n438) );
  XNOR2_X1 U494 ( .A(n439), .B(n438), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n440), .B(KEYINPUT90), .ZN(n441) );
  XNOR2_X1 U496 ( .A(n441), .B(KEYINPUT91), .ZN(n442) );
  XOR2_X1 U497 ( .A(n443), .B(n442), .Z(n447) );
  XNOR2_X1 U498 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U500 ( .A(n449), .B(n448), .ZN(n525) );
  NAND2_X1 U501 ( .A1(n534), .A2(n525), .ZN(n452) );
  XOR2_X1 U502 ( .A(KEYINPUT115), .B(KEYINPUT54), .Z(n450) );
  NOR2_X1 U503 ( .A1(n521), .A2(n453), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n454), .B(KEYINPUT65), .ZN(n575) );
  NOR2_X1 U505 ( .A1(n473), .A2(n575), .ZN(n455) );
  XNOR2_X1 U506 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  XNOR2_X1 U507 ( .A(n457), .B(KEYINPUT116), .ZN(n570) );
  AND2_X1 U508 ( .A1(n570), .A2(n561), .ZN(n461) );
  XNOR2_X1 U509 ( .A(KEYINPUT120), .B(KEYINPUT58), .ZN(n459) );
  INV_X1 U510 ( .A(G190GAT), .ZN(n458) );
  NAND2_X1 U511 ( .A1(n570), .A2(n577), .ZN(n464) );
  XNOR2_X1 U512 ( .A(n462), .B(KEYINPUT117), .ZN(n463) );
  XNOR2_X1 U513 ( .A(n464), .B(n463), .ZN(G1348GAT) );
  XNOR2_X1 U514 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n483) );
  NAND2_X1 U515 ( .A1(n577), .A2(n582), .ZN(n494) );
  NOR2_X1 U516 ( .A1(n561), .A2(n545), .ZN(n465) );
  XNOR2_X1 U517 ( .A(n465), .B(KEYINPUT16), .ZN(n480) );
  INV_X1 U518 ( .A(n537), .ZN(n527) );
  AND2_X1 U519 ( .A1(n527), .A2(n525), .ZN(n466) );
  NOR2_X1 U520 ( .A1(n473), .A2(n466), .ZN(n467) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n467), .Z(n470) );
  NAND2_X1 U522 ( .A1(n473), .A2(n537), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(KEYINPUT26), .ZN(n576) );
  XOR2_X1 U524 ( .A(KEYINPUT27), .B(n525), .Z(n474) );
  NOR2_X1 U525 ( .A1(n576), .A2(n474), .ZN(n469) );
  NOR2_X1 U526 ( .A1(n470), .A2(n469), .ZN(n472) );
  NOR2_X1 U527 ( .A1(n472), .A2(n471), .ZN(n478) );
  XNOR2_X1 U528 ( .A(KEYINPUT28), .B(n473), .ZN(n540) );
  NOR2_X1 U529 ( .A1(n475), .A2(n474), .ZN(n535) );
  NAND2_X1 U530 ( .A1(n537), .A2(n535), .ZN(n476) );
  NOR2_X1 U531 ( .A1(n540), .A2(n476), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n478), .A2(n477), .ZN(n491) );
  INV_X1 U533 ( .A(n491), .ZN(n479) );
  NAND2_X1 U534 ( .A1(n480), .A2(n479), .ZN(n508) );
  NOR2_X1 U535 ( .A1(n494), .A2(n508), .ZN(n481) );
  XOR2_X1 U536 ( .A(KEYINPUT93), .B(n481), .Z(n488) );
  NAND2_X1 U537 ( .A1(n488), .A2(n521), .ZN(n482) );
  XNOR2_X1 U538 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U539 ( .A1(n525), .A2(n488), .ZN(n484) );
  XNOR2_X1 U540 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT94), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U542 ( .A1(n488), .A2(n527), .ZN(n485) );
  XNOR2_X1 U543 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U544 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n488), .A2(n540), .ZN(n489) );
  XNOR2_X1 U546 ( .A(n489), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT95), .B(KEYINPUT39), .Z(n498) );
  NOR2_X1 U548 ( .A1(n490), .A2(n491), .ZN(n492) );
  NAND2_X1 U549 ( .A1(n545), .A2(n492), .ZN(n493) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(n493), .Z(n518) );
  NOR2_X1 U551 ( .A1(n518), .A2(n494), .ZN(n496) );
  XNOR2_X1 U552 ( .A(KEYINPUT96), .B(KEYINPUT38), .ZN(n495) );
  XNOR2_X1 U553 ( .A(n496), .B(n495), .ZN(n505) );
  NAND2_X1 U554 ( .A1(n505), .A2(n521), .ZN(n497) );
  XNOR2_X1 U555 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U556 ( .A(G29GAT), .B(n499), .Z(G1328GAT) );
  XOR2_X1 U557 ( .A(G36GAT), .B(KEYINPUT97), .Z(n501) );
  NAND2_X1 U558 ( .A1(n505), .A2(n525), .ZN(n500) );
  XNOR2_X1 U559 ( .A(n501), .B(n500), .ZN(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT98), .B(KEYINPUT40), .Z(n503) );
  NAND2_X1 U561 ( .A1(n505), .A2(n527), .ZN(n502) );
  XNOR2_X1 U562 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U563 ( .A(G43GAT), .B(n504), .Z(G1330GAT) );
  NAND2_X1 U564 ( .A1(n505), .A2(n540), .ZN(n506) );
  XNOR2_X1 U565 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U566 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n510) );
  INV_X1 U567 ( .A(n577), .ZN(n507) );
  XOR2_X1 U568 ( .A(KEYINPUT99), .B(n555), .Z(n565) );
  NAND2_X1 U569 ( .A1(n507), .A2(n565), .ZN(n519) );
  NOR2_X1 U570 ( .A1(n519), .A2(n508), .ZN(n514) );
  NAND2_X1 U571 ( .A1(n514), .A2(n521), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U573 ( .A1(n525), .A2(n514), .ZN(n511) );
  XNOR2_X1 U574 ( .A(n511), .B(KEYINPUT100), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G64GAT), .B(n512), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n527), .A2(n514), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U579 ( .A1(n514), .A2(n540), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  XOR2_X1 U582 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n523) );
  NOR2_X1 U583 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U584 ( .A(n520), .B(KEYINPUT102), .ZN(n530) );
  NAND2_X1 U585 ( .A1(n530), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U588 ( .A1(n530), .A2(n525), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U590 ( .A(G99GAT), .B(KEYINPUT105), .Z(n529) );
  NAND2_X1 U591 ( .A1(n530), .A2(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(G1338GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n532) );
  NAND2_X1 U594 ( .A1(n540), .A2(n530), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U596 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  XOR2_X1 U597 ( .A(G113GAT), .B(KEYINPUT109), .Z(n542) );
  NAND2_X1 U598 ( .A1(n534), .A2(n535), .ZN(n536) );
  XOR2_X1 U599 ( .A(KEYINPUT107), .B(n536), .Z(n553) );
  NOR2_X1 U600 ( .A1(n537), .A2(n553), .ZN(n538) );
  XOR2_X1 U601 ( .A(KEYINPUT108), .B(n538), .Z(n539) );
  NOR2_X1 U602 ( .A1(n540), .A2(n539), .ZN(n550) );
  NAND2_X1 U603 ( .A1(n550), .A2(n577), .ZN(n541) );
  XNOR2_X1 U604 ( .A(n542), .B(n541), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U606 ( .A1(n550), .A2(n565), .ZN(n543) );
  XNOR2_X1 U607 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n549) );
  XOR2_X1 U609 ( .A(KEYINPUT111), .B(KEYINPUT110), .Z(n547) );
  INV_X1 U610 ( .A(n545), .ZN(n586) );
  NAND2_X1 U611 ( .A1(n550), .A2(n586), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .Z(n552) );
  NAND2_X1 U615 ( .A1(n550), .A2(n561), .ZN(n551) );
  XNOR2_X1 U616 ( .A(n552), .B(n551), .ZN(G1343GAT) );
  NOR2_X1 U617 ( .A1(n576), .A2(n553), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n577), .A2(n562), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT112), .ZN(n559) );
  XOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U622 ( .A1(n562), .A2(n555), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U625 ( .A1(n562), .A2(n586), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT113), .Z(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  XNOR2_X1 U630 ( .A(KEYINPUT57), .B(KEYINPUT118), .ZN(n569) );
  XOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT56), .Z(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n570), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  XOR2_X1 U635 ( .A(G183GAT), .B(KEYINPUT119), .Z(n572) );
  NAND2_X1 U636 ( .A1(n586), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT123), .B(KEYINPUT122), .Z(n574) );
  XNOR2_X1 U639 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n581) );
  XOR2_X1 U641 ( .A(G197GAT), .B(KEYINPUT121), .Z(n579) );
  NOR2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n587) );
  NAND2_X1 U643 ( .A1(n587), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XOR2_X1 U645 ( .A(n581), .B(n580), .Z(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U647 ( .A(n587), .ZN(n589) );
  OR2_X1 U648 ( .A1(n589), .A2(n582), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(n585), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n588), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n490), .A2(n589), .ZN(n591) );
  XNOR2_X1 U654 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n591), .B(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(n592), .B(KEYINPUT126), .Z(n594) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(KEYINPUT125), .ZN(n593) );
  XNOR2_X1 U658 ( .A(n594), .B(n593), .ZN(G1355GAT) );
endmodule

