//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:32 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n767, new_n769,
    new_n770, new_n771, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT32), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n188), .A2(new_n189), .ZN(new_n190));
  NOR2_X1   g004(.A1(G237), .A2(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G210), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n192), .B(KEYINPUT27), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT26), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT27), .ZN(new_n195));
  XNOR2_X1  g009(.A(new_n192), .B(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT26), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G101), .B1(new_n194), .B2(new_n198), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  INV_X1    g018(.A(G134), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G137), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(G137), .ZN(new_n207));
  INV_X1    g021(.A(G137), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n208), .A2(KEYINPUT11), .A3(G134), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n207), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G131), .ZN(new_n211));
  INV_X1    g025(.A(G131), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n206), .A2(new_n209), .A3(new_n212), .A4(new_n207), .ZN(new_n213));
  AND2_X1   g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT0), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G143), .B2(new_n215), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n223), .A2(KEYINPUT66), .A3(G146), .ZN(new_n224));
  OAI211_X1 g038(.A(new_n217), .B(new_n220), .C1(new_n222), .C2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT64), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(KEYINPUT0), .B2(G128), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n220), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n223), .A2(G146), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n215), .B2(G143), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n223), .A2(KEYINPUT65), .A3(G146), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n225), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n215), .A2(G143), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n223), .A2(KEYINPUT65), .A3(G146), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT65), .B1(new_n223), .B2(G146), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n219), .B1(new_n238), .B2(KEYINPUT1), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT66), .B1(new_n223), .B2(G146), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n221), .A2(new_n215), .A3(G143), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n216), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n247));
  AOI22_X1  g061(.A1(new_n241), .A2(new_n243), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n205), .A2(G137), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n208), .A2(G134), .ZN(new_n250));
  OAI21_X1  g064(.A(G131), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n213), .A2(new_n251), .ZN(new_n252));
  OAI22_X1  g066(.A1(new_n214), .A2(new_n237), .B1(new_n248), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G116), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT67), .B1(new_n254), .B2(G119), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  INV_X1    g070(.A(G119), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n256), .A2(new_n257), .A3(G116), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n255), .A2(new_n258), .B1(new_n254), .B2(G119), .ZN(new_n259));
  XOR2_X1   g073(.A(KEYINPUT2), .B(G113), .Z(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n259), .A2(new_n260), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(new_n264), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n253), .A2(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n217), .B(new_n247), .C1(new_n222), .C2(new_n224), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n236), .B2(new_n242), .ZN(new_n268));
  INV_X1    g082(.A(new_n252), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n220), .B1(new_n228), .B2(new_n226), .ZN(new_n271));
  AOI22_X1  g085(.A1(new_n241), .A2(new_n271), .B1(new_n246), .B2(new_n220), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n211), .A2(new_n213), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n264), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT28), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n274), .A2(new_n270), .A3(new_n264), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT28), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n203), .B1(new_n276), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT30), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n253), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n274), .A2(new_n270), .A3(KEYINPUT30), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n283), .A2(new_n265), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT31), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n285), .A2(new_n286), .A3(new_n277), .A4(new_n203), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n281), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n285), .A2(new_n277), .A3(new_n203), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n291), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT68), .B1(new_n291), .B2(KEYINPUT31), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n190), .B1(new_n290), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G472), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT29), .ZN(new_n297));
  XNOR2_X1  g111(.A(new_n199), .B(new_n200), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n276), .B2(new_n279), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n285), .A2(new_n277), .A3(new_n298), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n297), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n279), .ZN(new_n302));
  INV_X1    g116(.A(new_n275), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n277), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n304), .B2(KEYINPUT28), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n298), .A2(new_n297), .ZN(new_n306));
  AOI21_X1  g120(.A(G902), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n296), .B1(new_n301), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AND3_X1   g123(.A1(new_n274), .A2(new_n270), .A3(KEYINPUT30), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT30), .B1(new_n274), .B2(new_n270), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n266), .B1(new_n312), .B2(new_n265), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT69), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n313), .A2(new_n314), .A3(new_n286), .A4(new_n203), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n287), .A2(KEYINPUT69), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n280), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n291), .A2(KEYINPUT31), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT68), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n291), .A2(KEYINPUT68), .A3(KEYINPUT31), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n188), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n295), .B(new_n309), .C1(new_n323), .C2(KEYINPUT32), .ZN(new_n324));
  XOR2_X1   g138(.A(KEYINPUT70), .B(G217), .Z(new_n325));
  INV_X1    g139(.A(G234), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n328), .B1(new_n257), .B2(G128), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n329), .B(new_n330), .C1(G119), .C2(new_n219), .ZN(new_n331));
  XNOR2_X1  g145(.A(G119), .B(G128), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT24), .B(G110), .Z(new_n333));
  AOI22_X1  g147(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n335), .A2(G125), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n336), .A2(new_n338), .A3(KEYINPUT16), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n337), .A2(KEYINPUT16), .A3(G140), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(G146), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G146), .B1(new_n339), .B2(new_n340), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n334), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI22_X1  g158(.A1(new_n331), .A2(G110), .B1(new_n332), .B2(new_n333), .ZN(new_n345));
  XNOR2_X1  g159(.A(G125), .B(G140), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n215), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n345), .A2(new_n347), .A3(new_n341), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(G953), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(G221), .A3(G234), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT22), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(G137), .ZN(new_n354));
  XNOR2_X1  g168(.A(new_n351), .B(KEYINPUT22), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n208), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n349), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(KEYINPUT72), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT71), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n357), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n354), .A2(new_n356), .A3(KEYINPUT71), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n349), .ZN(new_n365));
  OR3_X1    g179(.A1(new_n349), .A2(KEYINPUT72), .A3(new_n357), .ZN(new_n366));
  INV_X1    g180(.A(G902), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n359), .A2(new_n365), .A3(new_n366), .A4(new_n367), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n327), .B1(new_n368), .B2(KEYINPUT25), .ZN(new_n369));
  AOI22_X1  g183(.A1(KEYINPUT72), .A2(new_n358), .B1(new_n364), .B2(new_n349), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n367), .A4(new_n366), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  AND2_X1   g187(.A1(new_n370), .A2(new_n366), .ZN(new_n374));
  AOI21_X1  g188(.A(G902), .B1(new_n325), .B2(new_n326), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n324), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT73), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n187), .B1(new_n290), .B2(new_n294), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n189), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n317), .A2(new_n322), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n308), .B1(new_n384), .B2(new_n190), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n377), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT73), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n381), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT3), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n389), .A2(new_n390), .A3(G104), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G107), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT74), .ZN(new_n395));
  OAI21_X1  g209(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n200), .A4(new_n396), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n396), .A2(new_n391), .A3(new_n200), .A4(new_n393), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n390), .A2(G104), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n200), .B1(new_n401), .B2(new_n393), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n254), .A2(G119), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n256), .B1(G116), .B2(new_n257), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n254), .A2(KEYINPUT67), .A3(G119), .ZN(new_n406));
  OAI211_X1 g220(.A(KEYINPUT5), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT5), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n257), .A3(G116), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n409), .A2(KEYINPUT77), .ZN(new_n410));
  INV_X1    g224(.A(G113), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(new_n409), .B2(KEYINPUT77), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n407), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n400), .A2(new_n403), .A3(new_n261), .A4(new_n413), .ZN(new_n414));
  XOR2_X1   g228(.A(G110), .B(G122), .Z(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n396), .A2(new_n391), .A3(new_n393), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(G101), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(KEYINPUT4), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n419), .B1(new_n397), .B2(new_n399), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT4), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n421), .A3(G101), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n422), .B1(new_n262), .B2(new_n263), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n414), .B(new_n416), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n267), .B(new_n337), .C1(new_n236), .C2(new_n242), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n425), .B1(new_n272), .B2(new_n337), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n350), .A2(G224), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n425), .B(new_n428), .C1(new_n272), .C2(new_n337), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(KEYINPUT79), .B(KEYINPUT8), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n415), .B(new_n433), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n403), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n413), .A2(new_n261), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n434), .B1(new_n439), .B2(new_n414), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n424), .B(new_n432), .C1(new_n440), .C2(KEYINPUT80), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT80), .ZN(new_n442));
  AOI211_X1 g256(.A(new_n442), .B(new_n434), .C1(new_n439), .C2(new_n414), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n367), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(KEYINPUT81), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT81), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n446), .B(new_n367), .C1(new_n441), .C2(new_n443), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n420), .A2(new_n423), .ZN(new_n448));
  INV_X1    g262(.A(new_n414), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n415), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT6), .A3(new_n424), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n427), .B(KEYINPUT78), .Z(new_n452));
  XNOR2_X1  g266(.A(new_n426), .B(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT6), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n454), .B(new_n415), .C1(new_n448), .C2(new_n449), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n451), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n445), .A2(new_n447), .A3(new_n456), .ZN(new_n457));
  OAI21_X1  g271(.A(G210), .B1(G237), .B2(G902), .ZN(new_n458));
  XOR2_X1   g272(.A(new_n458), .B(KEYINPUT82), .Z(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(G214), .B1(G237), .B2(G902), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n445), .A2(new_n459), .A3(new_n456), .A4(new_n447), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n461), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(KEYINPUT83), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT18), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n466), .A2(new_n212), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n191), .A2(G143), .A3(G214), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G143), .B1(new_n191), .B2(G214), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n336), .A2(new_n338), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(G146), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(new_n347), .ZN(new_n474));
  INV_X1    g288(.A(G237), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n350), .A3(G214), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n476), .A2(new_n223), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n477), .B(new_n468), .C1(new_n466), .C2(new_n212), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n471), .A2(new_n474), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT84), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT84), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n471), .A2(new_n474), .A3(new_n478), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n342), .A2(new_n343), .ZN(new_n484));
  OAI211_X1 g298(.A(KEYINPUT17), .B(G131), .C1(new_n469), .C2(new_n470), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT87), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(new_n343), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n487), .A2(new_n485), .A3(KEYINPUT87), .A4(new_n341), .ZN(new_n488));
  OAI21_X1  g302(.A(G131), .B1(new_n469), .B2(new_n470), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n477), .A2(new_n212), .A3(new_n468), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n483), .B1(new_n486), .B2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(G113), .B(G122), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT86), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n495), .A2(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n392), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n499), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(G104), .A3(new_n497), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n346), .A2(KEYINPUT19), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n346), .A2(KEYINPUT19), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n341), .B1(new_n507), .B2(G146), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT85), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT85), .ZN(new_n510));
  OAI211_X1 g324(.A(new_n510), .B(new_n341), .C1(new_n507), .C2(G146), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n489), .A2(new_n491), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n509), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n503), .B1(new_n480), .B2(new_n482), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n504), .A2(KEYINPUT88), .A3(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT20), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n494), .A2(new_n503), .B1(new_n513), .B2(new_n514), .ZN(new_n519));
  NOR2_X1   g333(.A1(G475), .A2(G902), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n516), .A2(new_n517), .A3(new_n519), .A4(new_n520), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(G234), .A2(G237), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n525), .A2(G952), .A3(new_n350), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(G902), .A3(G953), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n503), .A2(KEYINPUT89), .ZN(new_n532));
  AOI21_X1  g346(.A(G902), .B1(new_n494), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n533), .B1(new_n494), .B2(new_n532), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n531), .B1(new_n534), .B2(G475), .ZN(new_n535));
  XNOR2_X1  g349(.A(KEYINPUT9), .B(G234), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n325), .A3(new_n350), .ZN(new_n538));
  AND2_X1   g352(.A1(KEYINPUT90), .A2(G122), .ZN(new_n539));
  NOR2_X1   g353(.A1(KEYINPUT90), .A2(G122), .ZN(new_n540));
  OAI21_X1  g354(.A(G116), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n254), .A2(G122), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT91), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n541), .A2(new_n545), .A3(new_n542), .ZN(new_n546));
  AOI21_X1  g360(.A(G107), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(G122), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n548), .A2(G116), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n541), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT92), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n553), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n542), .A2(KEYINPUT92), .A3(KEYINPUT14), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n390), .B1(new_n552), .B2(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G128), .B(G143), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(G134), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n547), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n558), .A2(KEYINPUT13), .ZN(new_n561));
  NOR3_X1   g375(.A1(new_n219), .A2(KEYINPUT13), .A3(G143), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n562), .A2(new_n205), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n558), .A2(new_n205), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n546), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n545), .B1(new_n541), .B2(new_n542), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n390), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n544), .A2(G107), .A3(new_n546), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n566), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n538), .B1(new_n560), .B2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n566), .ZN(new_n573));
  NOR3_X1   g387(.A1(new_n567), .A2(new_n568), .A3(new_n390), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n573), .B1(new_n574), .B2(new_n547), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n552), .A2(new_n556), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n559), .B1(new_n576), .B2(G107), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n569), .ZN(new_n578));
  INV_X1    g392(.A(new_n538), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n572), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  AOI211_X1 g399(.A(G902), .B(new_n583), .C1(new_n572), .C2(new_n580), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n524), .A2(new_n535), .A3(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT83), .ZN(new_n589));
  NAND4_X1  g403(.A1(new_n461), .A2(new_n589), .A3(new_n462), .A4(new_n463), .ZN(new_n590));
  OAI21_X1  g404(.A(G221), .B1(new_n536), .B2(G902), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G140), .ZN(new_n593));
  AND2_X1   g407(.A1(new_n350), .A2(G227), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n402), .B1(new_n397), .B2(new_n399), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n267), .A2(KEYINPUT75), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT75), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n246), .A2(new_n599), .A3(new_n247), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n217), .B1(new_n222), .B2(new_n224), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n243), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n598), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  AND2_X1   g417(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(new_n597), .A2(new_n268), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n273), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT12), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n437), .A2(new_n248), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n597), .A2(new_n603), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n214), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT12), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n418), .ZN(new_n614));
  INV_X1    g428(.A(new_n422), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n237), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT10), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n241), .A2(new_n243), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n617), .B1(new_n618), .B2(new_n267), .ZN(new_n619));
  AOI22_X1  g433(.A1(new_n614), .A2(new_n616), .B1(new_n597), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n617), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n620), .A2(new_n214), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n596), .B1(new_n613), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n272), .A2(new_n422), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n268), .A2(KEYINPUT10), .ZN(new_n625));
  OAI22_X1  g439(.A1(new_n420), .A2(new_n624), .B1(new_n437), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT10), .B1(new_n597), .B2(new_n603), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n626), .A2(new_n273), .A3(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n214), .B1(new_n620), .B2(new_n621), .ZN(new_n629));
  NOR3_X1   g443(.A1(new_n628), .A2(new_n629), .A3(new_n595), .ZN(new_n630));
  OAI21_X1  g444(.A(KEYINPUT76), .B1(new_n623), .B2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n626), .A2(new_n627), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n595), .B1(new_n632), .B2(new_n214), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n273), .B1(new_n626), .B2(new_n627), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT76), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n628), .B1(new_n608), .B2(new_n612), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n635), .B(new_n636), .C1(new_n637), .C2(new_n596), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n631), .A2(G469), .A3(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G469), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n640), .A2(new_n367), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n611), .A2(KEYINPUT12), .ZN(new_n642));
  AOI211_X1 g456(.A(new_n607), .B(new_n214), .C1(new_n609), .C2(new_n610), .ZN(new_n643));
  OAI211_X1 g457(.A(new_n622), .B(new_n596), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n595), .B1(new_n628), .B2(new_n629), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n641), .B1(new_n646), .B2(new_n640), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n592), .B1(new_n639), .B2(new_n647), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n465), .A2(new_n588), .A3(new_n590), .A4(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(KEYINPUT93), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n648), .A2(new_n588), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT93), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n651), .A2(new_n465), .A3(new_n652), .A4(new_n590), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n388), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G101), .ZN(G3));
  NAND2_X1  g469(.A1(new_n464), .A2(KEYINPUT94), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT94), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n461), .A2(new_n657), .A3(new_n462), .A4(new_n463), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n572), .A2(KEYINPUT33), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT96), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n575), .A2(new_n578), .A3(new_n663), .A4(new_n579), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n660), .A2(new_n661), .A3(new_n662), .A4(new_n664), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n572), .A2(new_n664), .A3(KEYINPUT33), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n580), .A2(KEYINPUT96), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT97), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(KEYINPUT33), .B1(new_n572), .B2(new_n580), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT95), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n582), .A2(G902), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n572), .A2(new_n580), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n367), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(new_n582), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n534), .A2(G475), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n504), .A2(new_n515), .ZN(new_n679));
  INV_X1    g493(.A(new_n520), .ZN(new_n680));
  NOR4_X1   g494(.A1(new_n679), .A2(KEYINPUT88), .A3(KEYINPUT20), .A4(new_n680), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n516), .A2(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n678), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n531), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n659), .A2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n648), .ZN(new_n687));
  AOI21_X1  g501(.A(G902), .B1(new_n317), .B2(new_n322), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n382), .B1(new_n688), .B2(new_n296), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n687), .A2(new_n377), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n686), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT34), .B(G104), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G6));
  INV_X1    g507(.A(new_n587), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n519), .A2(KEYINPUT20), .A3(new_n520), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT20), .B1(new_n519), .B2(new_n520), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n694), .A2(new_n535), .A3(new_n697), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n659), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n690), .ZN(new_n700));
  XOR2_X1   g514(.A(KEYINPUT35), .B(G107), .Z(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G9));
  OAI21_X1  g516(.A(new_n349), .B1(new_n364), .B2(KEYINPUT36), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT36), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n363), .A2(new_n704), .A3(new_n344), .A4(new_n348), .ZN(new_n705));
  AND3_X1   g519(.A1(new_n703), .A2(new_n375), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n369), .B2(new_n372), .ZN(new_n707));
  INV_X1    g521(.A(new_n707), .ZN(new_n708));
  OAI211_X1 g522(.A(new_n382), .B(new_n708), .C1(new_n688), .C2(new_n296), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(KEYINPUT98), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n650), .A2(new_n653), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT37), .B(G110), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G12));
  AND3_X1   g527(.A1(new_n324), .A2(new_n648), .A3(new_n708), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n528), .A2(G900), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT99), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(KEYINPUT99), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n526), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n719), .B1(new_n534), .B2(G475), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n697), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n694), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n714), .A2(new_n659), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G128), .ZN(G30));
  XNOR2_X1  g539(.A(new_n718), .B(KEYINPUT39), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n648), .A2(KEYINPUT40), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(KEYINPUT40), .B1(new_n648), .B2(new_n726), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT101), .ZN(new_n729));
  OR3_X1    g543(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n729), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n461), .A2(new_n463), .ZN(new_n732));
  XOR2_X1   g546(.A(new_n732), .B(KEYINPUT38), .Z(new_n733));
  OAI21_X1  g547(.A(new_n367), .B1(new_n304), .B2(new_n203), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n298), .B1(new_n285), .B2(new_n277), .ZN(new_n735));
  OAI21_X1  g549(.A(G472), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT100), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n738), .B(G472), .C1(new_n734), .C2(new_n735), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n740), .B1(new_n384), .B2(new_n190), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n383), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n462), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n683), .A2(new_n694), .ZN(new_n745));
  NOR4_X1   g559(.A1(new_n743), .A2(new_n744), .A3(new_n708), .A4(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n730), .A2(new_n731), .A3(new_n733), .A4(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G143), .ZN(G45));
  AOI21_X1  g562(.A(new_n707), .B1(new_n383), .B2(new_n385), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n677), .A2(new_n683), .A3(new_n718), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n659), .A2(new_n648), .A3(new_n749), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  NAND2_X1  g567(.A1(new_n634), .A2(new_n622), .ZN(new_n754));
  AOI22_X1  g568(.A1(new_n613), .A2(new_n633), .B1(new_n754), .B2(new_n595), .ZN(new_n755));
  OAI21_X1  g569(.A(G469), .B1(new_n755), .B2(G902), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n644), .A2(new_n645), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n640), .A3(new_n367), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(KEYINPUT102), .A3(new_n758), .ZN(new_n759));
  OR3_X1    g573(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n640), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n591), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n379), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n686), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(KEYINPUT41), .B(G113), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(G15));
  NAND2_X1  g580(.A1(new_n699), .A2(new_n763), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G116), .ZN(G18));
  AOI21_X1  g582(.A(new_n762), .B1(new_n656), .B2(new_n658), .ZN(new_n769));
  AND3_X1   g583(.A1(new_n324), .A2(new_n588), .A3(new_n708), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G119), .ZN(G21));
  INV_X1    g586(.A(new_n531), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n761), .A2(new_n591), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(new_n318), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n187), .B1(new_n290), .B2(new_n775), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n378), .B(new_n776), .C1(new_n296), .C2(new_n688), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n745), .B1(new_n656), .B2(new_n658), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  OAI211_X1 g595(.A(new_n776), .B(new_n708), .C1(new_n688), .C2(new_n296), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n750), .ZN(new_n783));
  INV_X1    g597(.A(new_n762), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n659), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  XOR2_X1   g599(.A(KEYINPUT103), .B(G125), .Z(new_n786));
  XNOR2_X1  g600(.A(new_n785), .B(new_n786), .ZN(G27));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n744), .B1(new_n461), .B2(new_n463), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n635), .B(G469), .C1(new_n637), .C2(new_n596), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n592), .B1(new_n647), .B2(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n324), .A2(new_n378), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n788), .B1(new_n792), .B2(new_n750), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n789), .A2(new_n791), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(new_n751), .A3(KEYINPUT42), .A4(new_n386), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n793), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G131), .ZN(G33));
  INV_X1    g612(.A(KEYINPUT104), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n792), .B2(new_n722), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n795), .A2(KEYINPUT104), .A3(new_n386), .A4(new_n723), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  INV_X1    g617(.A(new_n683), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT43), .B1(new_n677), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT43), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n806), .B1(new_n673), .B2(new_n676), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n683), .A2(KEYINPUT106), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT106), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n524), .A2(new_n809), .A3(new_n678), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n807), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT107), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n808), .A2(new_n810), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT107), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n807), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n805), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT108), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n689), .A2(new_n708), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(KEYINPUT109), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(KEYINPUT108), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT44), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n635), .B1(new_n637), .B2(new_n596), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT45), .ZN(new_n825));
  OAI21_X1  g639(.A(G469), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n631), .A2(new_n638), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n826), .B1(new_n827), .B2(new_n825), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT46), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n828), .A2(new_n829), .A3(new_n641), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n829), .B1(new_n828), .B2(new_n641), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n830), .A2(new_n758), .A3(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n591), .A3(new_n726), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT105), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n817), .A2(new_n819), .A3(KEYINPUT44), .A4(new_n820), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n823), .A2(new_n834), .A3(new_n789), .A4(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n836), .B(G137), .ZN(G39));
  INV_X1    g651(.A(KEYINPUT47), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT110), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n832), .A2(new_n839), .A3(new_n591), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n839), .B1(new_n832), .B2(new_n591), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n832), .A2(new_n591), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(KEYINPUT110), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n832), .A2(new_n839), .A3(new_n591), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(KEYINPUT47), .A3(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n789), .ZN(new_n847));
  NOR4_X1   g661(.A1(new_n847), .A2(new_n324), .A3(new_n750), .A4(new_n378), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n842), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  XNOR2_X1  g663(.A(new_n849), .B(G140), .ZN(G42));
  AND4_X1   g664(.A1(new_n462), .A2(new_n677), .A3(new_n378), .A4(new_n591), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n851), .B(new_n813), .C1(new_n852), .C2(new_n761), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT111), .Z(new_n854));
  AOI211_X1 g668(.A(new_n742), .B(new_n733), .C1(new_n852), .C2(new_n761), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT119), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT114), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n812), .A2(new_n815), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n858), .B(new_n527), .C1(new_n859), .C2(new_n805), .ZN(new_n860));
  OAI21_X1  g674(.A(KEYINPUT114), .B1(new_n816), .B2(new_n526), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n777), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n862), .A2(new_n789), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n842), .A2(new_n846), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g679(.A(new_n761), .B(KEYINPUT116), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(new_n592), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT117), .Z(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n864), .B1(new_n842), .B2(new_n846), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n863), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n762), .A2(new_n847), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n872), .A2(new_n527), .A3(new_n378), .A4(new_n743), .ZN(new_n873));
  OR3_X1    g687(.A1(new_n873), .A2(new_n683), .A3(new_n677), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n860), .A2(new_n861), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n872), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n874), .B1(new_n876), .B2(new_n782), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT50), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n462), .B(new_n733), .C1(KEYINPUT118), .C2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n862), .A2(new_n784), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(KEYINPUT118), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n862), .A2(new_n784), .A3(new_n881), .A4(new_n879), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n871), .A2(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n857), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n862), .A2(new_n659), .A3(new_n784), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(KEYINPUT120), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT120), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n862), .A2(new_n891), .A3(new_n659), .A4(new_n784), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(G952), .B(new_n350), .C1(new_n873), .C2(new_n684), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n875), .A2(new_n386), .A3(new_n872), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(KEYINPUT48), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT48), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n875), .A2(new_n897), .A3(new_n386), .A4(new_n872), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n894), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n893), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n842), .A2(new_n846), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(new_n867), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n887), .B1(new_n902), .B2(new_n863), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n885), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n675), .A2(new_n583), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n581), .A2(new_n584), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n905), .A2(new_n906), .A3(KEYINPUT112), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT112), .ZN(new_n908));
  OAI21_X1  g722(.A(new_n908), .B1(new_n585), .B2(new_n586), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n804), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n531), .B1(new_n684), .B2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n690), .A2(new_n465), .A3(new_n590), .A4(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n654), .A2(new_n711), .A3(new_n913), .ZN(new_n914));
  NOR3_X1   g728(.A1(new_n794), .A2(new_n750), .A3(new_n782), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT113), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n324), .A2(new_n648), .A3(new_n708), .ZN(new_n917));
  INV_X1    g731(.A(new_n910), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n789), .A2(new_n721), .A3(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n916), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n697), .A2(new_n907), .A3(new_n909), .A4(new_n720), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n744), .B(new_n921), .C1(new_n463), .C2(new_n461), .ZN(new_n922));
  NAND4_X1  g736(.A1(new_n922), .A2(new_n749), .A3(KEYINPUT113), .A4(new_n648), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n915), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI22_X1  g738(.A1(new_n769), .A2(new_n770), .B1(new_n778), .B2(new_n779), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n763), .B(new_n659), .C1(new_n685), .C2(new_n698), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n797), .A2(new_n802), .ZN(new_n928));
  NOR3_X1   g742(.A1(new_n914), .A2(new_n927), .A3(new_n928), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n706), .B(new_n719), .C1(new_n369), .C2(new_n372), .ZN(new_n930));
  INV_X1    g744(.A(new_n641), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n758), .A2(new_n931), .A3(new_n790), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n930), .A2(new_n932), .A3(new_n591), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n383), .B2(new_n741), .ZN(new_n934));
  INV_X1    g748(.A(new_n745), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n659), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n724), .A2(new_n752), .A3(new_n936), .A4(new_n785), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT52), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n714), .B(new_n659), .C1(new_n723), .C2(new_n751), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n940), .A2(KEYINPUT52), .A3(new_n785), .A4(new_n936), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(KEYINPUT53), .B1(new_n929), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n927), .A2(new_n928), .ZN(new_n944));
  INV_X1    g758(.A(new_n914), .ZN(new_n945));
  AND4_X1   g759(.A1(KEYINPUT53), .A2(new_n944), .A3(new_n942), .A4(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(KEYINPUT54), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT53), .ZN(new_n948));
  INV_X1    g762(.A(new_n927), .ZN(new_n949));
  INV_X1    g763(.A(new_n928), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n942), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n929), .A2(KEYINPUT53), .A3(new_n942), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT54), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n900), .A2(new_n904), .A3(new_n947), .A4(new_n956), .ZN(new_n957));
  AOI211_X1 g771(.A(KEYINPUT119), .B(KEYINPUT51), .C1(new_n871), .C2(new_n885), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n888), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(G952), .A2(G953), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n856), .B1(new_n959), .B2(new_n960), .ZN(G75));
  NAND2_X1  g775(.A1(new_n953), .A2(new_n954), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n962), .A2(G902), .A3(new_n459), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT56), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n451), .A2(new_n455), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(new_n453), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n966), .B(KEYINPUT121), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT55), .Z(new_n968));
  AND3_X1   g782(.A1(new_n963), .A2(new_n964), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n963), .B2(new_n964), .ZN(new_n970));
  NOR2_X1   g784(.A1(new_n350), .A2(G952), .ZN(new_n971));
  NOR3_X1   g785(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(G51));
  NAND2_X1  g786(.A1(new_n947), .A2(new_n956), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n641), .B(KEYINPUT57), .ZN(new_n974));
  AOI21_X1  g788(.A(KEYINPUT122), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT122), .ZN(new_n976));
  INV_X1    g790(.A(new_n974), .ZN(new_n977));
  AOI211_X1 g791(.A(new_n976), .B(new_n977), .C1(new_n947), .C2(new_n956), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n757), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n828), .B(KEYINPUT123), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n962), .A2(G902), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n971), .B1(new_n979), .B2(new_n981), .ZN(G54));
  AND2_X1   g796(.A1(KEYINPUT58), .A2(G475), .ZN(new_n983));
  OAI211_X1 g797(.A(G902), .B(new_n983), .C1(new_n943), .C2(new_n946), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n679), .ZN(new_n985));
  INV_X1    g799(.A(new_n971), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n962), .A2(G902), .A3(new_n519), .A4(new_n983), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(G60));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT59), .Z(new_n991));
  AOI21_X1  g805(.A(new_n991), .B1(new_n947), .B2(new_n956), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n669), .A2(new_n671), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n986), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n993), .B2(new_n992), .ZN(G63));
  AOI21_X1  g809(.A(KEYINPUT60), .B1(G217), .B2(G902), .ZN(new_n996));
  AND3_X1   g810(.A1(KEYINPUT60), .A2(G217), .A3(G902), .ZN(new_n997));
  OAI22_X1  g811(.A1(new_n943), .A2(new_n946), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n374), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n971), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AND2_X1   g814(.A1(new_n703), .A2(new_n705), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(new_n998), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT61), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1003), .B(new_n1004), .ZN(G66));
  NAND3_X1  g819(.A1(new_n945), .A2(new_n926), .A3(new_n925), .ZN(new_n1006));
  NAND2_X1  g820(.A1(G224), .A2(G953), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n1006), .A2(G953), .B1(new_n530), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n965), .B1(G898), .B2(new_n350), .ZN(new_n1009));
  XOR2_X1   g823(.A(new_n1008), .B(new_n1009), .Z(G69));
  AND2_X1   g824(.A1(new_n940), .A2(new_n785), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n950), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n779), .A2(new_n386), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n834), .B2(new_n1013), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1014), .A2(new_n836), .A3(new_n350), .A4(new_n849), .ZN(new_n1015));
  XOR2_X1   g829(.A(new_n312), .B(new_n507), .Z(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n350), .B1(G227), .B2(G900), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n747), .A2(new_n1011), .ZN(new_n1025));
  INV_X1    g839(.A(KEYINPUT62), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n747), .A2(KEYINPUT62), .A3(new_n1011), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n847), .B1(new_n684), .B2(new_n911), .ZN(new_n1030));
  NAND4_X1  g844(.A1(new_n388), .A2(new_n648), .A3(new_n726), .A4(new_n1030), .ZN(new_n1031));
  NAND4_X1  g845(.A1(new_n836), .A2(new_n1029), .A3(new_n849), .A4(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1032), .A2(new_n350), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1017), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1016), .B1(new_n1032), .B2(new_n350), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT125), .ZN(new_n1038));
  NAND4_X1  g852(.A1(new_n1024), .A2(new_n1036), .A3(new_n1019), .A4(new_n1038), .ZN(new_n1039));
  AOI21_X1  g853(.A(new_n1022), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1040));
  OAI21_X1  g854(.A(new_n1019), .B1(new_n1037), .B2(KEYINPUT125), .ZN(new_n1041));
  AOI211_X1 g855(.A(new_n1035), .B(new_n1016), .C1(new_n1032), .C2(new_n350), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  AND2_X1   g857(.A1(new_n1039), .A2(new_n1043), .ZN(G72));
  NAND2_X1  g858(.A1(G472), .A2(G902), .ZN(new_n1045));
  XOR2_X1   g859(.A(new_n1045), .B(KEYINPUT63), .Z(new_n1046));
  OAI21_X1  g860(.A(new_n1046), .B1(new_n1032), .B2(new_n1006), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n1047), .A2(new_n735), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1014), .A2(new_n836), .A3(new_n849), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1046), .B1(new_n1049), .B2(new_n1006), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1050), .A2(new_n300), .ZN(new_n1051));
  INV_X1    g865(.A(new_n300), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1052), .A2(new_n1046), .ZN(new_n1053));
  NOR2_X1   g867(.A1(new_n1053), .A2(new_n735), .ZN(new_n1054));
  AOI21_X1  g868(.A(new_n971), .B1(new_n962), .B2(new_n1054), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1048), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  INV_X1    g870(.A(KEYINPUT127), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND4_X1  g872(.A1(new_n1048), .A2(new_n1051), .A3(KEYINPUT127), .A4(new_n1055), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n1058), .A2(new_n1059), .ZN(G57));
endmodule


