//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n725, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n812, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n933, new_n934, new_n935, new_n936, new_n937;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  INV_X1    g001(.A(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n204), .B(KEYINPUT80), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT31), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT81), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT72), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT22), .ZN(new_n209));
  INV_X1    g008(.A(G197gat), .ZN(new_n210));
  INV_X1    g009(.A(G204gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(G197gat), .A2(G204gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n209), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(G211gat), .ZN(new_n215));
  INV_X1    g014(.A(G218gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G211gat), .A2(G218gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n208), .B1(new_n214), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g019(.A1(G197gat), .A2(G204gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(G197gat), .A2(G204gat), .ZN(new_n222));
  OAI21_X1  g021(.A(KEYINPUT22), .B1(new_n221), .B2(new_n222), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n223), .A2(KEYINPUT72), .A3(new_n218), .A4(new_n217), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n218), .B1(new_n217), .B2(new_n209), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n212), .A2(new_n213), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n220), .A2(new_n224), .A3(new_n227), .ZN(new_n228));
  NOR2_X1   g027(.A1(G155gat), .A2(G162gat), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT2), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G155gat), .A2(G162gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n235));
  INV_X1    g034(.A(G141gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n234), .A2(G141gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n233), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n229), .ZN(new_n243));
  XNOR2_X1  g042(.A(G141gat), .B(G148gat), .ZN(new_n244));
  OAI211_X1 g043(.A(new_n232), .B(new_n243), .C1(new_n244), .C2(KEYINPUT2), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n242), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT77), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT77), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n242), .A2(new_n248), .A3(new_n245), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT29), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n228), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  AOI21_X1  g052(.A(KEYINPUT3), .B1(new_n228), .B2(new_n252), .ZN(new_n254));
  INV_X1    g053(.A(KEYINPUT75), .ZN(new_n255));
  AND2_X1   g054(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(KEYINPUT74), .A2(G141gat), .ZN(new_n257));
  OAI21_X1  g056(.A(G148gat), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI22_X1  g057(.A1(new_n258), .A2(new_n240), .B1(new_n232), .B2(new_n231), .ZN(new_n259));
  XNOR2_X1  g058(.A(G155gat), .B(G162gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n236), .A2(G148gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n240), .A2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n260), .B1(new_n230), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n255), .B1(new_n259), .B2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n242), .A2(KEYINPUT75), .A3(new_n245), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n254), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(G228gat), .A2(G233gat), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n253), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT82), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n269), .B1(new_n214), .B2(new_n219), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n223), .A2(KEYINPUT82), .A3(new_n218), .A4(new_n217), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(new_n227), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(KEYINPUT83), .A3(new_n252), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(new_n249), .ZN(new_n274));
  AOI21_X1  g073(.A(KEYINPUT83), .B1(new_n272), .B2(new_n252), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n246), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT84), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n253), .ZN(new_n279));
  OAI211_X1 g078(.A(KEYINPUT84), .B(new_n246), .C1(new_n274), .C2(new_n275), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n268), .B1(new_n281), .B2(new_n267), .ZN(new_n282));
  INV_X1    g081(.A(G22gat), .ZN(new_n283));
  AND2_X1   g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n282), .A2(new_n283), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n207), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n267), .ZN(new_n287));
  INV_X1    g086(.A(new_n268), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(G22gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n282), .A2(new_n283), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT85), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n206), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n286), .B1(new_n292), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n264), .A2(new_n265), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT3), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  INV_X1    g097(.A(G127gat), .ZN(new_n299));
  NOR2_X1   g098(.A1(new_n299), .A2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G127gat), .ZN(new_n302));
  OAI22_X1  g101(.A1(new_n298), .A2(KEYINPUT1), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G120gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G113gat), .ZN(new_n305));
  INV_X1    g104(.A(G113gat), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(G120gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G127gat), .B(G134gat), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT1), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT76), .B1(new_n303), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n303), .A2(new_n311), .A3(KEYINPUT76), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n251), .A2(new_n297), .A3(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n303), .A2(new_n311), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n246), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n316), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  OR2_X1    g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n318), .B1(new_n315), .B2(new_n296), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n322), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(KEYINPUT39), .A3(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n327), .B(KEYINPUT0), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(G57gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n329), .B(G85gat), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n326), .B(new_n331), .C1(KEYINPUT39), .C2(new_n323), .ZN(new_n332));
  XNOR2_X1  g131(.A(new_n332), .B(KEYINPUT40), .ZN(new_n333));
  NOR2_X1   g132(.A1(G183gat), .A2(G190gat), .ZN(new_n334));
  AND2_X1   g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(KEYINPUT24), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(KEYINPUT24), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g136(.A1(G169gat), .A2(G176gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT23), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(G169gat), .B2(G176gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(G169gat), .A2(G176gat), .ZN(new_n342));
  AND3_X1   g141(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n337), .A2(KEYINPUT25), .A3(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT66), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n345), .B1(new_n335), .B2(KEYINPUT24), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT66), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n336), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n343), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT67), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT67), .ZN(new_n353));
  AOI211_X1 g152(.A(new_n353), .B(KEYINPUT25), .C1(new_n349), .C2(new_n343), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n344), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g154(.A(KEYINPUT27), .B(G183gat), .ZN(new_n356));
  INV_X1    g155(.A(G190gat), .ZN(new_n357));
  AOI21_X1  g156(.A(KEYINPUT28), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  AND2_X1   g158(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT28), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n359), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT69), .ZN(new_n364));
  INV_X1    g163(.A(new_n335), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT68), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT26), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n366), .B1(new_n338), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n338), .A2(new_n367), .ZN(new_n369));
  OAI211_X1 g168(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n368), .A2(new_n342), .A3(new_n369), .A4(new_n370), .ZN(new_n371));
  NAND4_X1  g170(.A1(new_n363), .A2(new_n364), .A3(new_n365), .A4(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n362), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n358), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n365), .ZN(new_n375));
  OAI21_X1  g174(.A(KEYINPUT69), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  AND2_X1   g176(.A1(G226gat), .A2(G233gat), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n355), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(KEYINPUT29), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n363), .A2(new_n365), .A3(new_n371), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n381), .B1(new_n355), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n228), .B1(new_n379), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n355), .A2(new_n382), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n355), .A2(new_n377), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n387), .A2(new_n378), .B1(new_n388), .B2(new_n380), .ZN(new_n389));
  INV_X1    g188(.A(new_n228), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  OAI211_X1 g190(.A(KEYINPUT73), .B(new_n228), .C1(new_n379), .C2(new_n383), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n386), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  XNOR2_X1  g192(.A(G8gat), .B(G36gat), .ZN(new_n394));
  INV_X1    g193(.A(G64gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(G92gat), .ZN(new_n397));
  XNOR2_X1  g196(.A(new_n396), .B(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n398), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n386), .A2(new_n391), .A3(new_n392), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n399), .A2(KEYINPUT30), .A3(new_n401), .ZN(new_n402));
  OR3_X1    g201(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n398), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT79), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n259), .A2(new_n263), .A3(new_n255), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT75), .B1(new_n242), .B2(new_n245), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n303), .A2(new_n311), .A3(KEYINPUT76), .ZN(new_n408));
  OAI22_X1  g207(.A1(new_n406), .A2(new_n407), .B1(new_n408), .B2(new_n312), .ZN(new_n409));
  INV_X1    g208(.A(new_n318), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n322), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT5), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n405), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT78), .ZN(new_n414));
  OAI211_X1 g213(.A(KEYINPUT79), .B(KEYINPUT5), .C1(new_n324), .C2(new_n322), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n321), .A2(new_n322), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n413), .A2(KEYINPUT78), .A3(new_n415), .ZN(new_n419));
  AND4_X1   g218(.A1(KEYINPUT5), .A2(new_n316), .A3(new_n320), .A4(new_n322), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AND3_X1   g220(.A1(new_n418), .A2(new_n421), .A3(KEYINPUT86), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT86), .B1(new_n418), .B2(new_n421), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n330), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n333), .A2(new_n404), .A3(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n393), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT37), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n400), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n427), .B2(new_n426), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT38), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(new_n401), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n418), .A2(new_n421), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n432), .A2(new_n433), .A3(new_n331), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n417), .A2(new_n416), .B1(new_n419), .B2(new_n420), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n433), .B1(new_n435), .B2(new_n330), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n434), .B1(new_n424), .B2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT38), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n389), .A2(new_n228), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n390), .B1(new_n379), .B2(new_n383), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n440), .A2(KEYINPUT37), .A3(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n295), .B(new_n425), .C1(new_n431), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G227gat), .A2(G233gat), .ZN(new_n446));
  XOR2_X1   g245(.A(new_n446), .B(KEYINPUT64), .Z(new_n447));
  XNOR2_X1  g246(.A(new_n447), .B(KEYINPUT65), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n317), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n355), .A2(new_n377), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n355), .B2(new_n377), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n449), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT33), .ZN(new_n454));
  XNOR2_X1  g253(.A(G15gat), .B(G43gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n455), .B(G71gat), .ZN(new_n456));
  INV_X1    g255(.A(G99gat), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n456), .B(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n453), .B(KEYINPUT32), .C1(new_n454), .C2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n459), .B1(new_n453), .B2(new_n454), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n453), .A2(KEYINPUT32), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n461), .A2(KEYINPUT70), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT70), .B1(new_n461), .B2(new_n462), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n388), .A2(new_n317), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n355), .A2(new_n377), .A3(new_n450), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT34), .B1(new_n468), .B2(new_n447), .ZN(new_n469));
  NOR2_X1   g268(.A1(new_n449), .A2(KEYINPUT34), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n466), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n472), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n474), .B(new_n460), .C1(new_n463), .C2(new_n464), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n477));
  OR2_X1    g276(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n476), .B1(KEYINPUT71), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n402), .A2(new_n403), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n432), .A2(new_n331), .ZN(new_n483));
  NOR2_X1   g282(.A1(new_n436), .A2(new_n483), .ZN(new_n484));
  NOR3_X1   g283(.A1(new_n432), .A2(new_n433), .A3(new_n331), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n482), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n293), .B1(new_n284), .B2(new_n285), .ZN(new_n487));
  INV_X1    g286(.A(new_n206), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n488), .B1(new_n290), .B2(KEYINPUT85), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n290), .A2(new_n291), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n487), .A2(new_n489), .B1(new_n490), .B2(new_n207), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n445), .A2(new_n481), .A3(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT88), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n476), .A2(new_n491), .ZN(new_n495));
  OAI21_X1  g294(.A(KEYINPUT87), .B1(new_n438), .B2(new_n404), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n432), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n418), .A2(new_n421), .A3(KEYINPUT86), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n436), .B1(new_n502), .B2(new_n330), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n498), .B(new_n482), .C1(new_n503), .C2(new_n434), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT35), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n494), .B1(new_n497), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n295), .A2(new_n473), .A3(new_n475), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n482), .B1(new_n503), .B2(new_n434), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(KEYINPUT87), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n424), .A2(new_n437), .ZN(new_n511));
  INV_X1    g310(.A(new_n434), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n511), .A2(new_n512), .B1(new_n403), .B2(new_n402), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT35), .B1(new_n513), .B2(new_n498), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n510), .A2(new_n514), .A3(KEYINPUT88), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n507), .A2(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(KEYINPUT35), .B1(new_n508), .B2(new_n486), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(KEYINPUT89), .B(KEYINPUT35), .C1(new_n508), .C2(new_n486), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n493), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT14), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(G29gat), .A2(G36gat), .ZN(new_n526));
  MUX2_X1   g325(.A(new_n525), .B(KEYINPUT14), .S(new_n526), .Z(new_n527));
  INV_X1    g326(.A(KEYINPUT91), .ZN(new_n528));
  XOR2_X1   g327(.A(G43gat), .B(G50gat), .Z(new_n529));
  AOI21_X1  g328(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n527), .A2(new_n529), .ZN(new_n531));
  OAI21_X1  g330(.A(KEYINPUT15), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(KEYINPUT15), .B2(new_n530), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT17), .ZN(new_n534));
  XNOR2_X1  g333(.A(new_n533), .B(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G15gat), .B(G22gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT16), .ZN(new_n537));
  AOI21_X1  g336(.A(G1gat), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G8gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n538), .B(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n536), .A2(KEYINPUT92), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  OR2_X1    g342(.A1(new_n533), .A2(new_n542), .ZN(new_n544));
  NAND2_X1  g343(.A1(G229gat), .A2(G233gat), .ZN(new_n545));
  AND3_X1   g344(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n546), .A2(KEYINPUT18), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n533), .B(new_n542), .ZN(new_n548));
  XOR2_X1   g347(.A(new_n545), .B(KEYINPUT13), .Z(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n546), .A2(KEYINPUT18), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n547), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n553));
  XNOR2_X1  g352(.A(G113gat), .B(G141gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(G169gat), .B(G197gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n557), .B(KEYINPUT12), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n547), .A2(new_n560), .A3(new_n550), .A4(new_n551), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AND2_X1   g362(.A1(new_n395), .A2(G57gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n395), .A2(G57gat), .ZN(new_n565));
  INV_X1    g364(.A(G71gat), .ZN(new_n566));
  INV_X1    g365(.A(G78gat), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  OAI22_X1  g367(.A1(new_n564), .A2(new_n565), .B1(new_n568), .B2(KEYINPUT9), .ZN(new_n569));
  XNOR2_X1  g368(.A(G71gat), .B(G78gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT93), .ZN(new_n572));
  NAND2_X1  g371(.A1(G85gat), .A2(G92gat), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(KEYINPUT7), .ZN(new_n574));
  NAND2_X1  g373(.A1(G99gat), .A2(G106gat), .ZN(new_n575));
  INV_X1    g374(.A(G85gat), .ZN(new_n576));
  AOI22_X1  g375(.A1(KEYINPUT8), .A2(new_n575), .B1(new_n576), .B2(new_n397), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G99gat), .B(G106gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n572), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT98), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT98), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n572), .A2(new_n583), .A3(new_n580), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT99), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n579), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(new_n578), .B(new_n586), .Z(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  AOI22_X1  g387(.A1(new_n582), .A2(new_n584), .B1(new_n571), .B2(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(KEYINPUT100), .B(KEYINPUT10), .Z(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(new_n580), .B(KEYINPUT96), .Z(new_n593));
  INV_X1    g392(.A(KEYINPUT10), .ZN(new_n594));
  OR3_X1    g393(.A1(new_n593), .A2(new_n594), .A3(new_n572), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G230gat), .ZN(new_n597));
  INV_X1    g396(.A(G233gat), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G120gat), .B(G148gat), .ZN(new_n602));
  INV_X1    g401(.A(G176gat), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(new_n211), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n601), .B(new_n606), .C1(new_n600), .C2(new_n589), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n599), .B1(new_n592), .B2(new_n595), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n589), .A2(new_n600), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n605), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n563), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n572), .A2(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(G127gat), .B(G155gat), .Z(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(G183gat), .B(G211gat), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(G231gat), .A2(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  OAI21_X1  g419(.A(new_n542), .B1(new_n572), .B2(new_n613), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT95), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g422(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n624));
  XOR2_X1   g423(.A(new_n623), .B(new_n624), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n620), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n535), .A2(new_n593), .ZN(new_n628));
  NAND3_X1  g427(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n629));
  OAI211_X1 g428(.A(new_n628), .B(new_n629), .C1(new_n593), .C2(new_n533), .ZN(new_n630));
  XNOR2_X1  g429(.A(G190gat), .B(G218gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT97), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G134gat), .ZN(new_n635));
  INV_X1    g434(.A(G162gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n630), .B(new_n631), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n639), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n522), .A2(new_n612), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n484), .A2(new_n485), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g447(.A1(new_n645), .A2(new_n404), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT101), .ZN(new_n650));
  OR3_X1    g449(.A1(new_n650), .A2(new_n537), .A3(KEYINPUT42), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n537), .B1(new_n650), .B2(KEYINPUT42), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n649), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n539), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n654), .B1(KEYINPUT42), .B2(new_n649), .ZN(G1325gat));
  INV_X1    g454(.A(new_n476), .ZN(new_n656));
  AOI21_X1  g455(.A(G15gat), .B1(new_n645), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n481), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n658), .A2(G15gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n657), .B1(new_n645), .B2(new_n659), .ZN(G1326gat));
  NAND2_X1  g459(.A1(new_n645), .A2(new_n491), .ZN(new_n661));
  XNOR2_X1  g460(.A(KEYINPUT43), .B(G22gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n661), .B(new_n662), .ZN(G1327gat));
  NAND2_X1  g462(.A1(new_n522), .A2(new_n643), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n612), .A2(new_n627), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n666), .A2(new_n523), .A3(new_n646), .ZN(new_n667));
  XOR2_X1   g466(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n507), .A2(new_n515), .A3(new_n519), .A4(new_n520), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n642), .B1(new_n670), .B2(new_n493), .ZN(new_n671));
  NOR2_X1   g470(.A1(KEYINPUT103), .A2(KEYINPUT44), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n671), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(KEYINPUT103), .B(KEYINPUT44), .Z(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  AOI211_X1 g475(.A(new_n642), .B(new_n676), .C1(new_n670), .C2(new_n493), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n678), .A2(new_n612), .A3(new_n627), .ZN(new_n679));
  INV_X1    g478(.A(new_n646), .ZN(new_n680));
  OAI21_X1  g479(.A(G29gat), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n669), .A2(new_n681), .ZN(G1328gat));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n524), .A3(new_n404), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(KEYINPUT46), .ZN(new_n684));
  XOR2_X1   g483(.A(new_n684), .B(KEYINPUT104), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n683), .A2(KEYINPUT46), .ZN(new_n686));
  OAI21_X1  g485(.A(G36gat), .B1(new_n679), .B2(new_n482), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(G1329gat));
  INV_X1    g487(.A(KEYINPUT105), .ZN(new_n689));
  OAI21_X1  g488(.A(G43gat), .B1(new_n679), .B2(new_n481), .ZN(new_n690));
  NOR4_X1   g489(.A1(new_n664), .A2(G43gat), .A3(new_n476), .A4(new_n665), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT106), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n690), .B2(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT47), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1330gat));
  OR3_X1    g494(.A1(new_n679), .A2(KEYINPUT109), .A3(new_n295), .ZN(new_n696));
  OAI21_X1  g495(.A(KEYINPUT109), .B1(new_n679), .B2(new_n295), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(G50gat), .A3(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(new_n295), .B2(G50gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n491), .A2(KEYINPUT108), .A3(new_n203), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n666), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n698), .A2(KEYINPUT48), .A3(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n679), .A2(new_n295), .ZN(new_n705));
  OAI21_X1  g504(.A(new_n703), .B1(new_n705), .B2(new_n203), .ZN(new_n706));
  XOR2_X1   g505(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n704), .A2(new_n708), .ZN(G1331gat));
  NOR3_X1   g508(.A1(new_n627), .A2(new_n643), .A3(new_n562), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n522), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n611), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(new_n646), .ZN(new_n714));
  XNOR2_X1  g513(.A(new_n714), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n482), .ZN(new_n716));
  NOR2_X1   g515(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n717));
  AND2_X1   g516(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n716), .B2(new_n717), .ZN(G1333gat));
  OAI21_X1  g519(.A(G71gat), .B1(new_n712), .B2(new_n481), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n656), .A2(new_n566), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n712), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g522(.A(new_n723), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g523(.A1(new_n712), .A2(new_n295), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n567), .ZN(G1335gat));
  INV_X1    g525(.A(new_n611), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n626), .A2(new_n562), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR4_X1   g528(.A1(new_n674), .A2(new_n677), .A3(new_n727), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(G85gat), .B1(new_n731), .B2(new_n680), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n522), .A2(KEYINPUT51), .A3(new_n643), .A4(new_n728), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT110), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n671), .A2(KEYINPUT110), .A3(KEYINPUT51), .A4(new_n728), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT111), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n664), .A2(new_n729), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n739), .A2(KEYINPUT51), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT111), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n735), .A2(new_n742), .A3(new_n736), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n744), .A2(new_n576), .A3(new_n646), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n732), .B1(new_n745), .B2(new_n727), .ZN(G1336gat));
  NOR3_X1   g545(.A1(new_n727), .A2(G92gat), .A3(new_n482), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  OR2_X1    g547(.A1(new_n739), .A2(KEYINPUT112), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT51), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n739), .A2(KEYINPUT112), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n748), .B1(new_n752), .B2(new_n737), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n397), .B1(new_n730), .B2(new_n404), .ZN(new_n754));
  OAI21_X1  g553(.A(KEYINPUT52), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n678), .A2(new_n611), .A3(new_n404), .A4(new_n728), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT52), .B1(new_n756), .B2(G92gat), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n735), .A2(new_n742), .A3(new_n736), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n742), .B1(new_n735), .B2(new_n736), .ZN(new_n759));
  NOR3_X1   g558(.A1(new_n758), .A2(new_n759), .A3(new_n740), .ZN(new_n760));
  OAI211_X1 g559(.A(KEYINPUT113), .B(new_n757), .C1(new_n760), .C2(new_n748), .ZN(new_n761));
  INV_X1    g560(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n744), .A2(new_n747), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT113), .B1(new_n763), .B2(new_n757), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n755), .B1(new_n762), .B2(new_n764), .ZN(G1337gat));
  OAI21_X1  g564(.A(G99gat), .B1(new_n731), .B2(new_n481), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n744), .A2(new_n457), .A3(new_n656), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n727), .ZN(G1338gat));
  INV_X1    g567(.A(G106gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n611), .A2(new_n491), .A3(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n752), .B2(new_n737), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n769), .B1(new_n730), .B2(new_n491), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT53), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(KEYINPUT53), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n774), .B1(new_n760), .B2(new_n770), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1339gat));
  NAND3_X1  g575(.A1(new_n592), .A2(new_n599), .A3(new_n595), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n601), .A2(KEYINPUT54), .A3(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT54), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n606), .B1(new_n608), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g579(.A1(new_n778), .A2(KEYINPUT55), .A3(new_n780), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n781), .A2(new_n607), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n778), .A2(new_n780), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT55), .ZN(new_n784));
  AOI21_X1  g583(.A(KEYINPUT115), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n786));
  AOI211_X1 g585(.A(new_n786), .B(KEYINPUT55), .C1(new_n778), .C2(new_n780), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n782), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT116), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n782), .B(KEYINPUT116), .C1(new_n785), .C2(new_n787), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n563), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n545), .B1(new_n543), .B2(new_n544), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n548), .A2(new_n549), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n557), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  AND2_X1   g594(.A1(new_n561), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n611), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT117), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n642), .B1(new_n792), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n790), .A2(new_n791), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n643), .A3(new_n796), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n626), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n710), .A2(new_n727), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT114), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n710), .A2(new_n805), .A3(new_n727), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g606(.A1(new_n802), .A2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n808), .A2(new_n646), .A3(new_n482), .A4(new_n495), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n563), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(new_n306), .ZN(G1340gat));
  NOR2_X1   g610(.A1(new_n809), .A2(new_n727), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(new_n304), .ZN(G1341gat));
  NOR2_X1   g612(.A1(new_n809), .A2(new_n627), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(new_n299), .ZN(G1342gat));
  NOR2_X1   g614(.A1(new_n809), .A2(new_n642), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n301), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(KEYINPUT56), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT56), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n819), .A3(new_n301), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n818), .B(new_n820), .C1(new_n301), .C2(new_n816), .ZN(G1343gat));
  NOR3_X1   g620(.A1(new_n658), .A2(new_n680), .A3(new_n404), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n783), .A2(new_n784), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(KEYINPUT118), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT118), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n783), .A2(new_n826), .A3(new_n784), .ZN(new_n827));
  NAND4_X1  g626(.A1(new_n825), .A2(new_n782), .A3(new_n562), .A4(new_n827), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n643), .B1(new_n828), .B2(new_n797), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n626), .B1(new_n801), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n491), .B1(new_n807), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n823), .B1(new_n832), .B2(KEYINPUT57), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT57), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n834), .B(new_n491), .C1(new_n802), .C2(new_n807), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n833), .A2(new_n562), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n237), .A2(new_n238), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT119), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n808), .A2(new_n840), .A3(new_n646), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n646), .B1(new_n802), .B2(new_n807), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n404), .B1(new_n842), .B2(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n481), .A2(new_n491), .ZN(new_n844));
  XNOR2_X1  g643(.A(new_n844), .B(KEYINPUT120), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n563), .A2(G141gat), .ZN(new_n846));
  NAND4_X1  g645(.A1(new_n841), .A2(new_n843), .A3(new_n845), .A4(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT121), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n839), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n849), .A2(KEYINPUT58), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT58), .ZN(new_n851));
  NAND4_X1  g650(.A1(new_n839), .A2(new_n847), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n850), .A2(new_n852), .ZN(G1344gat));
  NOR2_X1   g652(.A1(new_n727), .A2(G148gat), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n841), .A2(new_n843), .A3(new_n845), .A4(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n833), .A2(new_n835), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n856), .B1(new_n857), .B2(new_n727), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n234), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n643), .A2(new_n796), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n788), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n627), .B1(new_n861), .B2(new_n829), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n295), .B1(new_n862), .B2(new_n803), .ZN(new_n863));
  OR3_X1    g662(.A1(new_n863), .A2(KEYINPUT122), .A3(KEYINPUT57), .ZN(new_n864));
  OAI211_X1 g663(.A(KEYINPUT57), .B(new_n491), .C1(new_n802), .C2(new_n807), .ZN(new_n865));
  OAI21_X1  g664(.A(KEYINPUT122), .B1(new_n863), .B2(KEYINPUT57), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n611), .A3(new_n822), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n856), .B1(new_n868), .B2(G148gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n855), .B1(new_n859), .B2(new_n869), .ZN(G1345gat));
  INV_X1    g669(.A(G155gat), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n857), .A2(new_n871), .A3(new_n627), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n841), .A2(new_n843), .A3(new_n626), .A4(new_n845), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n872), .B1(new_n871), .B2(new_n873), .ZN(G1346gat));
  NOR3_X1   g673(.A1(new_n857), .A2(new_n636), .A3(new_n642), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n841), .A2(new_n843), .A3(new_n643), .A4(new_n845), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n636), .B2(new_n876), .ZN(G1347gat));
  INV_X1    g676(.A(KEYINPUT123), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n508), .A2(new_n482), .ZN(new_n879));
  OAI221_X1 g678(.A(new_n680), .B1(new_n878), .B2(new_n879), .C1(new_n802), .C2(new_n807), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n878), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(G169gat), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n884), .A3(new_n562), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n808), .A2(new_n680), .A3(new_n879), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n887), .A2(new_n562), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT124), .B1(new_n888), .B2(G169gat), .ZN(new_n889));
  OAI211_X1 g688(.A(KEYINPUT124), .B(G169gat), .C1(new_n886), .C2(new_n563), .ZN(new_n890));
  INV_X1    g689(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n885), .B1(new_n889), .B2(new_n891), .ZN(G1348gat));
  AOI21_X1  g691(.A(G176gat), .B1(new_n883), .B2(new_n611), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n886), .A2(new_n603), .A3(new_n727), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n893), .A2(new_n894), .ZN(G1349gat));
  NAND3_X1  g694(.A1(new_n883), .A2(new_n626), .A3(new_n356), .ZN(new_n896));
  OAI21_X1  g695(.A(G183gat), .B1(new_n886), .B2(new_n627), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT60), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT60), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n896), .A2(new_n900), .A3(new_n897), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n899), .A2(new_n901), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n883), .A2(new_n357), .A3(new_n643), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n887), .A2(new_n643), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G190gat), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n904), .B(G190gat), .C1(new_n886), .C2(new_n642), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n903), .B1(new_n906), .B2(new_n908), .ZN(G1351gat));
  NOR2_X1   g708(.A1(new_n658), .A2(new_n482), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  OAI21_X1  g710(.A(KEYINPUT125), .B1(new_n911), .B2(new_n295), .ZN(new_n912));
  OR3_X1    g711(.A1(new_n911), .A2(KEYINPUT125), .A3(new_n295), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n808), .A2(new_n680), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n915), .A2(new_n210), .A3(new_n562), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n911), .A2(new_n646), .ZN(new_n917));
  AND2_X1   g716(.A1(new_n867), .A2(new_n917), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(new_n562), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n916), .B1(new_n919), .B2(new_n210), .ZN(G1352gat));
  NAND2_X1  g719(.A1(new_n915), .A2(new_n611), .ZN(new_n921));
  XOR2_X1   g720(.A(KEYINPUT126), .B(G204gat), .Z(new_n922));
  OAI21_X1  g721(.A(KEYINPUT62), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  OR4_X1    g722(.A1(KEYINPUT62), .A2(new_n914), .A3(new_n727), .A4(new_n922), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n867), .A2(new_n611), .A3(new_n917), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n922), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(G1353gat));
  NAND3_X1  g726(.A1(new_n915), .A2(new_n215), .A3(new_n626), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n867), .A2(new_n626), .A3(new_n917), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n929), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT63), .B1(new_n929), .B2(G211gat), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(G1354gat));
  NAND3_X1  g731(.A1(new_n918), .A2(G218gat), .A3(new_n643), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n216), .B1(new_n914), .B2(new_n642), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  OAI211_X1 g735(.A(KEYINPUT127), .B(new_n216), .C1(new_n914), .C2(new_n642), .ZN(new_n937));
  AND3_X1   g736(.A1(new_n933), .A2(new_n936), .A3(new_n937), .ZN(G1355gat));
endmodule


