//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n491, new_n492, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n575, new_n576, new_n577, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n617, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1182;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT67), .Z(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n459), .A2(G2105), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G101), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G137), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n462), .A2(G125), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(new_n463), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(new_n469), .ZN(G160));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n459), .ZN(new_n472));
  NAND2_X1  g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n463), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n463), .A2(G112), .ZN(new_n476));
  OAI21_X1  g051(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n477));
  OAI21_X1  g052(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g053(.A(G2105), .B1(new_n472), .B2(new_n473), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n478), .B1(G136), .B2(new_n479), .ZN(new_n480));
  XOR2_X1   g055(.A(new_n480), .B(KEYINPUT68), .Z(G162));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n482));
  INV_X1    g057(.A(G138), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n482), .B1(new_n464), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(KEYINPUT4), .A3(G138), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n474), .A2(G126), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  OAI211_X1 g062(.A(new_n487), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n484), .A2(new_n485), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(G164));
  INV_X1    g065(.A(KEYINPUT6), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G651), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT69), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n494), .B1(new_n491), .B2(G651), .ZN(new_n495));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n496), .A2(KEYINPUT69), .A3(KEYINPUT6), .ZN(new_n497));
  OAI211_X1 g072(.A(G543), .B(new_n493), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G50), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT69), .B1(new_n496), .B2(KEYINPUT6), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n494), .A2(new_n491), .A3(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT5), .A2(G543), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AND3_X1   g083(.A1(new_n503), .A2(new_n493), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G88), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n508), .A2(G62), .ZN(new_n511));
  AND2_X1   g086(.A1(G75), .A2(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(G651), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n500), .A2(new_n510), .A3(new_n513), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND4_X1  g090(.A1(new_n503), .A2(G89), .A3(new_n493), .A4(new_n508), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  AND2_X1   g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  OAI21_X1  g096(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n506), .A2(KEYINPUT70), .A3(new_n507), .ZN(new_n523));
  AND2_X1   g098(.A1(G63), .A2(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g100(.A1(new_n516), .A2(new_n518), .A3(new_n525), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n498), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n492), .B1(new_n501), .B2(new_n502), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(KEYINPUT71), .A3(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n526), .B1(new_n531), .B2(G51), .ZN(G168));
  INV_X1    g107(.A(G52), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n528), .B2(new_n530), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n522), .A2(new_n523), .A3(G64), .ZN(new_n535));
  NAND2_X1  g110(.A1(G77), .A2(G543), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n496), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n529), .A2(G90), .A3(new_n508), .ZN(new_n538));
  NOR3_X1   g113(.A1(new_n534), .A2(new_n537), .A3(new_n538), .ZN(G171));
  INV_X1    g114(.A(KEYINPUT72), .ZN(new_n540));
  INV_X1    g115(.A(G43), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(new_n528), .B2(new_n530), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n509), .A2(G81), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND4_X1   g119(.A1(KEYINPUT71), .A2(new_n503), .A3(G543), .A4(new_n493), .ZN(new_n545));
  AOI21_X1  g120(.A(KEYINPUT71), .B1(new_n529), .B2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(G43), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n509), .A2(G81), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(KEYINPUT72), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n522), .A2(new_n523), .ZN(new_n551));
  INV_X1    g126(.A(G56), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI22_X1  g128(.A1(new_n544), .A2(new_n549), .B1(G651), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT73), .Z(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  NAND3_X1  g135(.A1(new_n529), .A2(G53), .A3(G543), .ZN(new_n561));
  OR2_X1    g136(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n520), .A2(new_n521), .ZN(new_n566));
  INV_X1    g141(.A(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n565), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n568), .A2(G651), .ZN(new_n569));
  INV_X1    g144(.A(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n529), .A2(new_n508), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n564), .A2(new_n573), .ZN(G299));
  NAND2_X1  g149(.A1(new_n535), .A2(new_n536), .ZN(new_n575));
  AOI22_X1  g150(.A1(new_n575), .A2(G651), .B1(new_n509), .B2(G90), .ZN(new_n576));
  OAI21_X1  g151(.A(G52), .B1(new_n545), .B2(new_n546), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G301));
  OAI21_X1  g153(.A(G51), .B1(new_n545), .B2(new_n546), .ZN(new_n579));
  INV_X1    g154(.A(new_n526), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G286));
  INV_X1    g156(.A(new_n551), .ZN(new_n582));
  OAI21_X1  g157(.A(G651), .B1(new_n582), .B2(G74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n499), .A2(G49), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI211_X1 g160(.A(new_n583), .B(new_n584), .C1(new_n585), .C2(new_n571), .ZN(G288));
  NAND2_X1  g161(.A1(new_n499), .A2(G48), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n509), .A2(G86), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n508), .A2(G61), .ZN(new_n589));
  AND2_X1   g164(.A1(G73), .A2(G543), .ZN(new_n590));
  OAI21_X1  g165(.A(G651), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g166(.A1(new_n587), .A2(new_n588), .A3(new_n591), .ZN(G305));
  NAND2_X1  g167(.A1(new_n531), .A2(G47), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G60), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n551), .B2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(KEYINPUT74), .B(G85), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n596), .A2(G651), .B1(new_n509), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n593), .A2(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND3_X1  g175(.A1(new_n509), .A2(KEYINPUT10), .A3(G92), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n571), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n566), .B2(new_n606), .ZN(new_n607));
  AOI22_X1  g182(.A1(new_n601), .A2(new_n604), .B1(G651), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n531), .A2(G54), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(new_n610), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n600), .B1(new_n611), .B2(G868), .ZN(G321));
  XNOR2_X1  g188(.A(G299), .B(KEYINPUT75), .ZN(new_n614));
  MUX2_X1   g189(.A(new_n614), .B(G286), .S(G868), .Z(G297));
  MUX2_X1   g190(.A(new_n614), .B(G286), .S(G868), .Z(G280));
  INV_X1    g191(.A(G559), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n611), .B1(new_n617), .B2(G860), .ZN(G148));
  OAI21_X1  g193(.A(KEYINPUT77), .B1(new_n554), .B2(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n611), .A2(new_n617), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT76), .ZN(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  MUX2_X1   g198(.A(KEYINPUT77), .B(new_n619), .S(new_n623), .Z(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n462), .A2(new_n460), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  INV_X1    g203(.A(G2100), .ZN(new_n629));
  OR2_X1    g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n628), .A2(new_n629), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n474), .A2(G123), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n479), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n463), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(new_n636), .B(G2096), .Z(new_n637));
  NAND3_X1  g212(.A1(new_n630), .A2(new_n631), .A3(new_n637), .ZN(G156));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n640), .A2(new_n641), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(KEYINPUT14), .A3(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT80), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G1341), .B(G1348), .Z(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(KEYINPUT78), .B(KEYINPUT16), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT79), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n647), .A2(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n654), .A2(new_n655), .A3(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XNOR2_X1  g232(.A(G2084), .B(G2090), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT81), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  OR2_X1    g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT82), .B(KEYINPUT17), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n660), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n661), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n658), .B(new_n662), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n665), .A2(new_n658), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n668), .B(KEYINPUT18), .Z(new_n669));
  NOR2_X1   g244(.A1(new_n661), .A2(new_n658), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n666), .A2(new_n669), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(new_n629), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT83), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XNOR2_X1  g251(.A(G1971), .B(G1976), .ZN(new_n677));
  INV_X1    g252(.A(KEYINPUT19), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XOR2_X1   g254(.A(G1956), .B(G2474), .Z(new_n680));
  XOR2_X1   g255(.A(G1961), .B(G1966), .Z(new_n681));
  AND2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT20), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n680), .A2(new_n681), .ZN(new_n685));
  NOR3_X1   g260(.A1(new_n679), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(new_n679), .B2(new_n685), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1981), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(G1986), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT84), .ZN(new_n694));
  OR2_X1    g269(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n692), .A2(new_n694), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n695), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n696), .B1(new_n695), .B2(new_n697), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n698), .A2(new_n699), .ZN(G229));
  INV_X1    g275(.A(G16), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n701), .A2(G23), .ZN(new_n702));
  INV_X1    g277(.A(G288), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n702), .B1(new_n703), .B2(new_n701), .ZN(new_n704));
  XNOR2_X1  g279(.A(KEYINPUT33), .B(G1976), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(G6), .A2(G16), .ZN(new_n707));
  INV_X1    g282(.A(G305), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G16), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n701), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n701), .ZN(new_n713));
  INV_X1    g288(.A(G1971), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n706), .A2(new_n711), .A3(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(KEYINPUT34), .ZN(new_n718));
  NOR2_X1   g293(.A1(G16), .A2(G24), .ZN(new_n719));
  INV_X1    g294(.A(G290), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n719), .B1(new_n720), .B2(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G1986), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n479), .A2(G131), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT85), .ZN(new_n724));
  OAI21_X1  g299(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n725));
  INV_X1    g300(.A(G107), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(G2105), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(new_n474), .B2(G119), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  MUX2_X1   g304(.A(G25), .B(new_n729), .S(G29), .Z(new_n730));
  XOR2_X1   g305(.A(KEYINPUT35), .B(G1991), .Z(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(KEYINPUT86), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n730), .B(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n721), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n691), .B2(new_n734), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n717), .A2(new_n718), .A3(new_n722), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT36), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n701), .A2(G19), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT87), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(new_n554), .B2(new_n701), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(G1341), .Z(new_n741));
  NOR2_X1   g316(.A1(G5), .A2(G16), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT94), .Z(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(G301), .B2(new_n701), .ZN(new_n744));
  INV_X1    g319(.A(G1961), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n701), .A2(G20), .ZN(new_n747));
  XOR2_X1   g322(.A(new_n747), .B(KEYINPUT96), .Z(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT23), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(G299), .B2(G16), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(G1956), .ZN(new_n751));
  INV_X1    g326(.A(G1348), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n611), .A2(G16), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n753), .B1(G4), .B2(G16), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  AOI211_X1 g330(.A(new_n746), .B(new_n755), .C1(new_n752), .C2(new_n754), .ZN(new_n756));
  INV_X1    g331(.A(G29), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G32), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n460), .A2(G105), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT92), .Z(new_n760));
  INV_X1    g335(.A(G141), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(new_n464), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n474), .A2(G129), .ZN(new_n763));
  NAND3_X1  g338(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n764), .A2(KEYINPUT26), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n764), .A2(KEYINPUT26), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n763), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(new_n762), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n758), .B1(new_n768), .B2(new_n757), .ZN(new_n769));
  XOR2_X1   g344(.A(KEYINPUT27), .B(G1996), .Z(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G27), .A2(G29), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G164), .B2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n771), .B1(G2078), .B2(new_n773), .ZN(new_n774));
  NOR2_X1   g349(.A1(G168), .A2(new_n701), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n701), .B2(G21), .ZN(new_n776));
  INV_X1    g351(.A(G1966), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n773), .A2(G2078), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n774), .A2(new_n778), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n479), .A2(G140), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n474), .A2(G128), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n463), .A2(G116), .ZN(new_n784));
  OAI21_X1  g359(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n782), .B(new_n783), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n786), .A2(G29), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n757), .A2(G26), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT28), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT88), .Z(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G2067), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G2067), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n757), .A2(G33), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT89), .B(KEYINPUT25), .Z(new_n795));
  NAND3_X1  g370(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n479), .A2(G139), .ZN(new_n798));
  AOI22_X1  g373(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n797), .B(new_n798), .C1(new_n463), .C2(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT90), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n794), .B1(new_n801), .B2(new_n757), .ZN(new_n802));
  OAI211_X1 g377(.A(new_n792), .B(new_n793), .C1(G2072), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n757), .A2(G35), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G162), .B2(new_n757), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G2090), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  XOR2_X1   g383(.A(KEYINPUT31), .B(G11), .Z(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT93), .ZN(new_n810));
  INV_X1    g385(.A(G28), .ZN(new_n811));
  OR2_X1    g386(.A1(new_n811), .A2(KEYINPUT30), .ZN(new_n812));
  AOI21_X1  g387(.A(G29), .B1(new_n811), .B2(KEYINPUT30), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  XOR2_X1   g389(.A(KEYINPUT91), .B(KEYINPUT24), .Z(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(G34), .ZN(new_n816));
  NOR2_X1   g391(.A1(new_n816), .A2(G29), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n817), .B1(G160), .B2(G29), .ZN(new_n818));
  OAI221_X1 g393(.A(new_n814), .B1(new_n757), .B2(new_n636), .C1(new_n818), .C2(G2084), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(G2084), .B2(new_n818), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n805), .A2(new_n807), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n802), .A2(G2072), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n808), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR3_X1   g398(.A1(new_n781), .A2(new_n803), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n737), .A2(new_n741), .A3(new_n756), .A4(new_n824), .ZN(G150));
  INV_X1    g400(.A(G150), .ZN(G311));
  NAND3_X1  g401(.A1(new_n522), .A2(new_n523), .A3(G67), .ZN(new_n827));
  NAND2_X1  g402(.A1(G80), .A2(G543), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT97), .B(G93), .Z(new_n830));
  AOI22_X1  g405(.A1(new_n829), .A2(G651), .B1(new_n509), .B2(new_n830), .ZN(new_n831));
  OAI21_X1  g406(.A(G55), .B1(new_n545), .B2(new_n546), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT98), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n833), .B1(new_n831), .B2(new_n832), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G860), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT37), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n553), .A2(G651), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n829), .A2(G651), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n509), .A2(new_n830), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(G55), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n528), .B2(new_n530), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n846), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n542), .A2(new_n543), .A3(new_n540), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT72), .B1(new_n547), .B2(new_n548), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n841), .B(new_n847), .C1(new_n848), .C2(new_n849), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n837), .B2(new_n554), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT38), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n610), .A2(new_n617), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT39), .ZN(new_n858));
  AOI21_X1  g433(.A(G860), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(KEYINPUT39), .A3(new_n856), .ZN(new_n860));
  AOI21_X1  g435(.A(KEYINPUT99), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n856), .ZN(new_n862));
  NOR2_X1   g437(.A1(new_n853), .A2(new_n854), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AND4_X1   g439(.A1(KEYINPUT99), .A2(new_n864), .A3(new_n860), .A4(new_n838), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n840), .B1(new_n861), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n868), .B(new_n840), .C1(new_n861), .C2(new_n865), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n867), .A2(new_n869), .ZN(G145));
  XNOR2_X1  g445(.A(new_n729), .B(new_n627), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n479), .A2(G142), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n474), .A2(G130), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n463), .A2(G118), .ZN(new_n874));
  OAI21_X1  g449(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n872), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n871), .B(new_n876), .Z(new_n877));
  INV_X1    g452(.A(KEYINPUT101), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(new_n489), .B(new_n786), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n768), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n800), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n883), .A2(new_n801), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n871), .B(new_n876), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n885), .A2(KEYINPUT101), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n879), .A2(new_n882), .A3(new_n884), .A4(new_n886), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(KEYINPUT102), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n879), .A2(new_n886), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n884), .A2(new_n882), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n467), .A2(new_n468), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(G2105), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n479), .A2(G137), .B1(G101), .B2(new_n460), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n636), .ZN(new_n897));
  XNOR2_X1  g472(.A(G162), .B(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n899), .B1(new_n890), .B2(new_n885), .ZN(new_n901));
  AOI21_X1  g476(.A(G37), .B1(new_n888), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  XNOR2_X1  g478(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n902), .A3(new_n904), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(G395));
  NAND2_X1  g483(.A1(new_n544), .A2(new_n549), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n909), .A2(new_n841), .A3(new_n847), .ZN(new_n910));
  OAI21_X1  g485(.A(KEYINPUT98), .B1(new_n844), .B2(new_n846), .ZN(new_n911));
  AOI22_X1  g486(.A1(new_n909), .A2(new_n841), .B1(new_n911), .B2(new_n834), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n621), .B(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n572), .B1(new_n562), .B2(new_n563), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n915), .A2(new_n609), .A3(new_n608), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n609), .B2(new_n608), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT41), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n610), .A2(G299), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT41), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(new_n921), .A3(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n914), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n917), .A2(new_n918), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n914), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n925), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n914), .A2(new_n926), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  XNOR2_X1  g506(.A(G166), .B(G288), .ZN(new_n932));
  NOR2_X1   g507(.A1(G290), .A2(new_n708), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n720), .A2(G305), .ZN(new_n934));
  OR3_X1    g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  AND3_X1   g513(.A1(new_n929), .A2(new_n931), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n938), .B1(new_n929), .B2(new_n931), .ZN(new_n940));
  OAI21_X1  g515(.A(G868), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g517(.A(new_n941), .B1(G868), .B2(new_n837), .ZN(G331));
  INV_X1    g518(.A(G37), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT105), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(G171), .B2(G286), .ZN(new_n946));
  NAND3_X1  g521(.A1(G301), .A2(KEYINPUT105), .A3(G168), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT106), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n948), .B1(G301), .B2(G168), .ZN(new_n949));
  NAND4_X1  g524(.A1(G286), .A2(KEYINPUT106), .A3(new_n577), .A4(new_n576), .ZN(new_n950));
  AOI22_X1  g525(.A1(new_n946), .A2(new_n947), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n851), .A2(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n851), .A2(new_n951), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n953), .A2(new_n926), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n946), .A2(new_n947), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n949), .A2(new_n950), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n912), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT107), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n958), .A2(new_n959), .A3(new_n960), .A4(new_n850), .ZN(new_n961));
  OAI21_X1  g536(.A(KEYINPUT107), .B1(new_n851), .B2(new_n951), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n961), .A2(new_n962), .B1(new_n851), .B2(new_n951), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n937), .B(new_n955), .C1(new_n963), .C2(new_n924), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n954), .A2(new_n926), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n965), .A2(new_n952), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n960), .B1(new_n913), .B2(new_n958), .ZN(new_n967));
  NOR3_X1   g542(.A1(new_n851), .A2(new_n951), .A3(KEYINPUT107), .ZN(new_n968));
  OAI21_X1  g543(.A(new_n954), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n966), .B1(new_n969), .B2(new_n923), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n935), .A2(KEYINPUT108), .A3(new_n936), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT108), .B1(new_n935), .B2(new_n936), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n944), .B(new_n964), .C1(new_n970), .C2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT43), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n926), .A2(KEYINPUT110), .A3(new_n921), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n977), .B1(new_n923), .B2(KEYINPUT110), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n978), .B1(new_n954), .B2(new_n953), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n965), .B1(new_n962), .B2(new_n961), .ZN(new_n980));
  OAI22_X1  g555(.A1(new_n979), .A2(new_n980), .B1(new_n971), .B2(new_n972), .ZN(new_n981));
  AND4_X1   g556(.A1(KEYINPUT43), .A2(new_n981), .A3(new_n944), .A4(new_n964), .ZN(new_n982));
  OAI21_X1  g557(.A(KEYINPUT44), .B1(new_n976), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT109), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n974), .A2(new_n984), .A3(KEYINPUT43), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n984), .B1(new_n974), .B2(KEYINPUT43), .ZN(new_n986));
  AND4_X1   g561(.A1(new_n975), .A2(new_n981), .A3(new_n944), .A4(new_n964), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n983), .B1(new_n988), .B2(KEYINPUT44), .ZN(G397));
  NAND3_X1  g564(.A1(new_n894), .A2(G40), .A3(new_n895), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(G160), .A2(KEYINPUT111), .A3(G40), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n489), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g573(.A1(new_n994), .A2(new_n998), .A3(G1996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n768), .ZN(new_n1000));
  XOR2_X1   g575(.A(new_n1000), .B(KEYINPUT112), .Z(new_n1001));
  INV_X1    g576(.A(G2067), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n786), .B(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(G1996), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1003), .B1(new_n768), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n994), .A2(new_n998), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n1006), .B(KEYINPUT113), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1001), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(new_n1007), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n729), .B(new_n731), .ZN(new_n1010));
  XOR2_X1   g585(.A(new_n1010), .B(KEYINPUT114), .Z(new_n1011));
  OAI21_X1  g586(.A(new_n1008), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(G290), .B(G1986), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1012), .B1(new_n1006), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n996), .A2(KEYINPUT50), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n489), .A2(new_n1016), .A3(new_n995), .ZN(new_n1017));
  NAND4_X1  g592(.A1(new_n1015), .A2(new_n1017), .A3(new_n992), .A4(new_n993), .ZN(new_n1018));
  XOR2_X1   g593(.A(KEYINPUT121), .B(G2084), .Z(new_n1019));
  OR2_X1    g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n489), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n998), .A2(new_n992), .A3(new_n993), .A4(new_n1021), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n1022), .A2(KEYINPUT120), .A3(new_n777), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT120), .B1(new_n1022), .B2(new_n777), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1020), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  AND2_X1   g600(.A1(new_n1025), .A2(G8), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(G286), .ZN(new_n1027));
  OAI211_X1 g602(.A(G168), .B(new_n1020), .C1(new_n1023), .C2(new_n1024), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(G8), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1029), .A2(KEYINPUT124), .A3(KEYINPUT51), .ZN(new_n1030));
  XOR2_X1   g605(.A(KEYINPUT124), .B(KEYINPUT51), .Z(new_n1031));
  NAND3_X1  g606(.A1(new_n1028), .A2(G8), .A3(new_n1031), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1027), .A2(new_n1030), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n1034));
  XNOR2_X1  g609(.A(KEYINPUT125), .B(KEYINPUT53), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1035), .B1(new_n1022), .B2(G2078), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1018), .A2(new_n745), .ZN(new_n1037));
  AND2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT53), .ZN(new_n1039));
  NOR3_X1   g614(.A1(new_n990), .A2(new_n1039), .A3(G2078), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n998), .A2(new_n1040), .A3(new_n1021), .ZN(new_n1041));
  XNOR2_X1  g616(.A(new_n1041), .B(KEYINPUT126), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1038), .A2(G301), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1043), .A2(KEYINPUT127), .ZN(new_n1044));
  AND2_X1   g619(.A1(new_n998), .A2(new_n1021), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n992), .A2(new_n993), .ZN(new_n1046));
  NOR2_X1   g621(.A1(new_n1039), .A2(G2078), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1038), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G171), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1044), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1043), .A2(KEYINPUT127), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1034), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(G303), .A2(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT55), .ZN(new_n1055));
  OR3_X1    g630(.A1(new_n1054), .A2(KEYINPUT116), .A3(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(KEYINPUT116), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1022), .A2(new_n714), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G2090), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1046), .A2(new_n1063), .A3(new_n1017), .A4(new_n1015), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1062), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1066));
  OAI211_X1 g641(.A(G8), .B(new_n1059), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  INV_X1    g643(.A(new_n996), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1068), .B1(new_n1046), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n703), .A2(G1976), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT52), .ZN(new_n1073));
  INV_X1    g648(.A(G1976), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT52), .B1(G288), .B2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1070), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT117), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n689), .B1(new_n591), .B2(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(G305), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(G305), .A2(new_n1078), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT49), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(KEYINPUT49), .A3(new_n1080), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1070), .A3(new_n1084), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n1073), .A2(new_n1076), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1068), .B1(new_n1060), .B2(new_n1064), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1059), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT119), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT119), .ZN(new_n1091));
  NOR3_X1   g666(.A1(new_n1087), .A2(new_n1091), .A3(new_n1059), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1067), .B(new_n1086), .C1(new_n1090), .C2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G301), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1094));
  AND4_X1   g669(.A1(G301), .A2(new_n1036), .A3(new_n1037), .A4(new_n1048), .ZN(new_n1095));
  NOR3_X1   g670(.A1(new_n1094), .A2(new_n1034), .A3(new_n1095), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1022), .A2(G1996), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT58), .B(G1341), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1099), .B1(new_n1046), .B2(new_n1069), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n554), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(KEYINPUT59), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT59), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n1103), .B(new_n554), .C1(new_n1098), .C2(new_n1100), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1018), .A2(new_n752), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1046), .A2(new_n1002), .A3(new_n1069), .ZN(new_n1107));
  AND3_X1   g682(.A1(new_n1106), .A2(new_n610), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n610), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1109));
  OAI21_X1  g684(.A(KEYINPUT60), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1106), .A2(new_n1107), .A3(new_n1111), .ZN(new_n1112));
  NAND3_X1  g687(.A1(new_n1105), .A2(new_n1110), .A3(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n1114));
  NAND2_X1  g689(.A1(G299), .A2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(KEYINPUT122), .A2(KEYINPUT57), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1115), .B(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT56), .B(G2072), .Z(new_n1120));
  INV_X1    g695(.A(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1045), .A2(new_n1119), .A3(new_n1046), .A4(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(G1956), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1018), .A2(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT123), .B1(new_n1022), .B2(new_n1120), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1118), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  AND4_X1   g702(.A1(new_n1118), .A2(new_n1126), .A3(new_n1124), .A4(new_n1122), .ZN(new_n1128));
  OAI21_X1  g703(.A(KEYINPUT61), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1118), .A3(new_n1126), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1118), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1132));
  INV_X1    g707(.A(new_n1126), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1131), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1130), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1113), .B1(new_n1129), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1130), .A2(new_n1109), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1134), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1053), .B(new_n1097), .C1(new_n1137), .C2(new_n1139), .ZN(new_n1140));
  NOR2_X1   g715(.A1(new_n1093), .A2(new_n1050), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1141), .B1(new_n1033), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1033), .B1(new_n1140), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1026), .A2(G168), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  AND2_X1   g721(.A1(new_n1067), .A2(new_n1086), .ZN(new_n1147));
  OAI21_X1  g722(.A(G8), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(new_n1089), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1146), .A2(KEYINPUT63), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1093), .A2(new_n1145), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1150), .B1(KEYINPUT63), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1033), .A2(new_n1141), .A3(KEYINPUT62), .ZN(new_n1153));
  XOR2_X1   g728(.A(new_n1070), .B(KEYINPUT118), .Z(new_n1154));
  NAND2_X1  g729(.A1(new_n708), .A2(new_n689), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1085), .A2(new_n1074), .A3(new_n703), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1154), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(new_n1067), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1157), .B1(new_n1158), .B2(new_n1086), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1152), .A2(new_n1153), .A3(new_n1159), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1014), .B1(new_n1144), .B2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n1008), .A2(new_n724), .A3(new_n728), .A4(new_n731), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n786), .A2(G2067), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1009), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n999), .B(KEYINPUT46), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n768), .A2(new_n1003), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1165), .B1(new_n1007), .B2(new_n1166), .ZN(new_n1167));
  XOR2_X1   g742(.A(new_n1167), .B(KEYINPUT47), .Z(new_n1168));
  NAND3_X1  g743(.A1(new_n1006), .A2(new_n691), .A3(new_n720), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT48), .Z(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1012), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1164), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1161), .A2(new_n1172), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g748(.A1(new_n656), .A2(G319), .A3(new_n675), .ZN(new_n1175));
  NOR3_X1   g749(.A1(new_n698), .A2(new_n699), .A3(new_n1175), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n888), .A2(new_n901), .ZN(new_n1177));
  NAND2_X1  g751(.A1(new_n1177), .A2(new_n944), .ZN(new_n1178));
  AOI21_X1  g752(.A(new_n898), .B1(new_n888), .B2(new_n891), .ZN(new_n1179));
  OAI21_X1  g753(.A(new_n1176), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g754(.A1(new_n988), .A2(new_n1180), .ZN(G308));
  OR2_X1    g755(.A1(new_n986), .A2(new_n987), .ZN(new_n1182));
  OAI211_X1 g756(.A(new_n903), .B(new_n1176), .C1(new_n1182), .C2(new_n985), .ZN(G225));
endmodule


