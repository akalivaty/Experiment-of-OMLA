//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:25 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n554, new_n555, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1195, new_n1196,
    new_n1197;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G137), .A3(new_n461), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n461), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  AND2_X1   g045(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n461), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G124), .ZN(new_n476));
  XOR2_X1   g051(.A(new_n476), .B(KEYINPUT67), .Z(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n472), .B2(new_n474), .ZN(new_n481));
  OR2_X1    g056(.A1(new_n481), .A2(KEYINPUT66), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n481), .A2(KEYINPUT66), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n480), .B1(G136), .B2(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n471), .C2(new_n473), .ZN(new_n487));
  OR2_X1    g062(.A1(G102), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n490), .A3(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n471), .B2(new_n473), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n497), .C1(new_n473), .C2(new_n471), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(G164));
  INV_X1    g074(.A(KEYINPUT6), .ZN(new_n500));
  INV_X1    g075(.A(G651), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(KEYINPUT68), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT68), .ZN(new_n503));
  NAND3_X1  g078(.A1(new_n503), .A2(KEYINPUT6), .A3(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(G50), .A3(G543), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  INV_X1    g082(.A(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g086(.A1(new_n505), .A2(G88), .A3(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n511), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  OAI211_X1 g088(.A(new_n506), .B(new_n512), .C1(new_n513), .C2(new_n501), .ZN(G303));
  INV_X1    g089(.A(G303), .ZN(G166));
  NAND3_X1  g090(.A1(new_n511), .A2(G63), .A3(G651), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT69), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n503), .A2(KEYINPUT6), .A3(G651), .ZN(new_n519));
  AOI21_X1  g094(.A(KEYINPUT6), .B1(new_n503), .B2(G651), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n502), .A2(KEYINPUT69), .A3(new_n504), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n517), .B1(new_n523), .B2(G51), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(KEYINPUT70), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n502), .A2(new_n504), .B1(new_n509), .B2(new_n510), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n527), .A2(KEYINPUT7), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n526), .A2(G89), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n524), .A2(KEYINPUT70), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n531), .A2(new_n532), .ZN(G168));
  NAND2_X1  g108(.A1(new_n523), .A2(G52), .ZN(new_n534));
  NAND2_X1  g109(.A1(G77), .A2(G543), .ZN(new_n535));
  AND2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(G64), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n535), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G651), .B1(new_n526), .B2(G90), .ZN(new_n541));
  AND2_X1   g116(.A1(new_n534), .A2(new_n541), .ZN(G171));
  NAND2_X1  g117(.A1(new_n526), .A2(G81), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n521), .A2(G543), .A3(new_n522), .ZN(new_n544));
  INV_X1    g119(.A(G43), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n543), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT71), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n511), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  OR2_X1    g123(.A1(new_n548), .A2(new_n501), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  NAND4_X1  g127(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  NAND4_X1  g131(.A1(new_n521), .A2(G53), .A3(G543), .A4(new_n522), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(KEYINPUT9), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n508), .B1(new_n505), .B2(new_n518), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND4_X1  g135(.A1(new_n559), .A2(new_n560), .A3(G53), .A4(new_n522), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(G78), .A2(G543), .ZN(new_n563));
  XOR2_X1   g138(.A(KEYINPUT72), .B(G65), .Z(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n538), .ZN(new_n565));
  AOI22_X1  g140(.A1(new_n565), .A2(G651), .B1(G91), .B2(new_n526), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g142(.A(new_n567), .B(KEYINPUT73), .ZN(G299));
  XOR2_X1   g143(.A(G171), .B(KEYINPUT74), .Z(G301));
  OR2_X1    g144(.A1(new_n531), .A2(new_n532), .ZN(G286));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n571), .B(G651), .C1(new_n511), .C2(G74), .ZN(new_n572));
  NAND2_X1  g147(.A1(G74), .A2(G651), .ZN(new_n573));
  OAI211_X1 g148(.A(KEYINPUT75), .B(new_n573), .C1(new_n538), .C2(new_n501), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n521), .A2(G49), .A3(G543), .A4(new_n522), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n526), .A2(G87), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n578), .A2(KEYINPUT76), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT76), .ZN(new_n580));
  NAND4_X1  g155(.A1(new_n575), .A2(new_n576), .A3(new_n580), .A4(new_n577), .ZN(new_n581));
  AND2_X1   g156(.A1(new_n579), .A2(new_n581), .ZN(G288));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n583), .B1(new_n509), .B2(new_n510), .ZN(new_n584));
  INV_X1    g159(.A(G73), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n585), .A2(new_n508), .ZN(new_n586));
  OAI21_X1  g161(.A(G651), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n505), .A2(G86), .A3(new_n511), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n505), .A2(G48), .A3(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(G305));
  NAND2_X1  g165(.A1(new_n526), .A2(G85), .ZN(new_n591));
  AOI22_X1  g166(.A1(new_n511), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G47), .ZN(new_n593));
  OAI221_X1 g168(.A(new_n591), .B1(new_n501), .B2(new_n592), .C1(new_n544), .C2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(new_n526), .A2(G92), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n595), .B(KEYINPUT10), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n511), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n501), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n523), .A2(G54), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n601), .A2(G868), .ZN(new_n602));
  XNOR2_X1  g177(.A(G171), .B(KEYINPUT74), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G284));
  AOI21_X1  g179(.A(new_n602), .B1(G868), .B2(new_n603), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NOR2_X1   g181(.A1(G286), .A2(new_n606), .ZN(new_n607));
  XOR2_X1   g182(.A(G299), .B(KEYINPUT77), .Z(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(new_n606), .ZN(G297));
  XNOR2_X1  g184(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g185(.A(new_n601), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  NOR2_X1   g188(.A1(new_n601), .A2(G559), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT79), .ZN(new_n615));
  MUX2_X1   g190(.A(new_n550), .B(new_n615), .S(G868), .Z(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n462), .A2(new_n467), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT12), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT13), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n475), .A2(G123), .ZN(new_n622));
  NOR2_X1   g197(.A1(new_n461), .A2(G111), .ZN(new_n623));
  OAI21_X1  g198(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI221_X1 g200(.A(new_n622), .B1(new_n623), .B2(new_n624), .C1(new_n484), .C2(new_n625), .ZN(new_n626));
  AOI22_X1  g201(.A1(new_n621), .A2(G2100), .B1(G2096), .B2(new_n626), .ZN(new_n627));
  OR2_X1    g202(.A1(new_n626), .A2(G2096), .ZN(new_n628));
  OAI211_X1 g203(.A(new_n627), .B(new_n628), .C1(G2100), .C2(new_n621), .ZN(G156));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2438), .ZN(new_n631));
  XOR2_X1   g206(.A(G2427), .B(G2430), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT81), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n631), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n631), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n638), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT82), .ZN(new_n645));
  INV_X1    g220(.A(G14), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n646), .B1(new_n642), .B2(new_n643), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(G401));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT84), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2084), .B(G2090), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT83), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT85), .B(KEYINPUT17), .ZN(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n651), .B2(new_n653), .ZN(new_n656));
  AOI21_X1  g231(.A(KEYINPUT18), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  XOR2_X1   g232(.A(KEYINPUT86), .B(G2100), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(G2072), .B(G2078), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n651), .A2(new_n653), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n660), .B1(new_n661), .B2(KEYINPUT18), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n659), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1971), .B(G1976), .Z(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT19), .ZN(new_n666));
  XOR2_X1   g241(.A(G1956), .B(G2474), .Z(new_n667));
  XOR2_X1   g242(.A(G1961), .B(G1966), .Z(new_n668));
  AND2_X1   g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n666), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n666), .A2(new_n669), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n666), .A2(new_n670), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(KEYINPUT88), .ZN(new_n676));
  OR2_X1    g251(.A1(new_n675), .A2(KEYINPUT88), .ZN(new_n677));
  AOI211_X1 g252(.A(new_n671), .B(new_n674), .C1(new_n676), .C2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT89), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1981), .B(G1986), .ZN(new_n684));
  INV_X1    g259(.A(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n683), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G229));
  XOR2_X1   g262(.A(KEYINPUT31), .B(G11), .Z(new_n688));
  INV_X1    g263(.A(G29), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT30), .B(G28), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n626), .B2(new_n689), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT96), .B(G2084), .Z(new_n693));
  OAI21_X1  g268(.A(G29), .B1(new_n465), .B2(new_n469), .ZN(new_n694));
  INV_X1    g269(.A(G34), .ZN(new_n695));
  AND2_X1   g270(.A1(new_n695), .A2(KEYINPUT24), .ZN(new_n696));
  NOR2_X1   g271(.A1(new_n695), .A2(KEYINPUT24), .ZN(new_n697));
  OAI21_X1  g272(.A(new_n689), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n693), .B1(new_n694), .B2(new_n698), .ZN(new_n699));
  AND3_X1   g274(.A1(new_n694), .A2(new_n693), .A3(new_n698), .ZN(new_n700));
  NOR3_X1   g275(.A1(new_n692), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(G2078), .ZN(new_n702));
  NOR2_X1   g277(.A1(G27), .A2(G29), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n703), .B1(G164), .B2(G29), .ZN(new_n704));
  XOR2_X1   g279(.A(new_n704), .B(KEYINPUT99), .Z(new_n705));
  OAI21_X1  g280(.A(new_n701), .B1(new_n702), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n689), .A2(G33), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n708));
  XOR2_X1   g283(.A(new_n708), .B(KEYINPUT25), .Z(new_n709));
  AOI22_X1  g284(.A1(new_n462), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n709), .B1(new_n710), .B2(new_n461), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(new_n485), .B2(G139), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n707), .B1(new_n712), .B2(new_n689), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(G2072), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n705), .A2(new_n702), .ZN(new_n715));
  INV_X1    g290(.A(G16), .ZN(new_n716));
  NOR2_X1   g291(.A1(G171), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(G5), .B2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(G1961), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  NAND4_X1  g296(.A1(new_n714), .A2(new_n715), .A3(new_n720), .A4(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n716), .A2(G4), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(new_n611), .B2(new_n716), .ZN(new_n724));
  AOI211_X1 g299(.A(new_n706), .B(new_n722), .C1(G1348), .C2(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n716), .A2(G19), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n726), .B1(new_n551), .B2(new_n716), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(G1341), .Z(new_n728));
  NAND2_X1  g303(.A1(new_n689), .A2(G26), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n729), .B(KEYINPUT28), .Z(new_n730));
  OAI21_X1  g305(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n731));
  INV_X1    g306(.A(G116), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G2105), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT94), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n475), .A2(G128), .ZN(new_n735));
  INV_X1    g310(.A(G140), .ZN(new_n736));
  OAI211_X1 g311(.A(new_n734), .B(new_n735), .C1(new_n484), .C2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT95), .ZN(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n730), .B1(new_n739), .B2(G29), .ZN(new_n740));
  INV_X1    g315(.A(G2067), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G2090), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n689), .A2(G35), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(G162), .B2(new_n689), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT29), .Z(new_n746));
  AOI21_X1  g321(.A(new_n742), .B1(new_n743), .B2(new_n746), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n725), .A2(new_n728), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n716), .A2(G21), .ZN(new_n749));
  OAI21_X1  g324(.A(new_n749), .B1(G168), .B2(new_n716), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n750), .A2(G1966), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n750), .A2(G1966), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n485), .A2(G141), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT97), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n756), .B(KEYINPUT98), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT26), .ZN(new_n758));
  AND2_X1   g333(.A1(new_n467), .A2(G105), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(G129), .B2(new_n475), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n755), .A2(new_n758), .A3(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G32), .B(new_n761), .S(G29), .Z(new_n762));
  XOR2_X1   g337(.A(KEYINPUT27), .B(G1996), .Z(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n762), .A2(new_n763), .ZN(new_n765));
  OAI211_X1 g340(.A(new_n764), .B(new_n765), .C1(G1348), .C2(new_n724), .ZN(new_n766));
  NOR4_X1   g341(.A1(new_n748), .A2(new_n751), .A3(new_n752), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n689), .A2(G25), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n485), .A2(G131), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n770));
  INV_X1    g345(.A(G107), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(G2105), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(new_n475), .B2(G119), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n768), .B1(new_n775), .B2(new_n689), .ZN(new_n776));
  XOR2_X1   g351(.A(KEYINPUT35), .B(G1991), .Z(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT90), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n776), .B(new_n778), .Z(new_n779));
  INV_X1    g354(.A(KEYINPUT91), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  MUX2_X1   g356(.A(G24), .B(G290), .S(G16), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1986), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  MUX2_X1   g359(.A(G6), .B(G305), .S(G16), .Z(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  INV_X1    g361(.A(G1981), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n716), .A2(G22), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G166), .B2(new_n716), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT93), .ZN(new_n791));
  INV_X1    g366(.A(G1971), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G23), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT92), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n578), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT92), .A4(new_n577), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n794), .B1(new_n798), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT33), .B(G1976), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n788), .A2(new_n793), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(KEYINPUT34), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n779), .A2(new_n780), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n784), .A2(new_n803), .A3(new_n804), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT36), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n716), .A2(G20), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT23), .Z(new_n809));
  AOI21_X1  g384(.A(new_n809), .B1(G299), .B2(G16), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G1956), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n746), .B2(new_n743), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n812), .A2(KEYINPUT100), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n812), .A2(KEYINPUT100), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n767), .A2(new_n807), .A3(new_n813), .A4(new_n814), .ZN(G150));
  INV_X1    g390(.A(G150), .ZN(G311));
  NAND2_X1  g391(.A1(new_n611), .A2(G559), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT38), .ZN(new_n818));
  AND2_X1   g393(.A1(new_n523), .A2(G55), .ZN(new_n819));
  XNOR2_X1  g394(.A(KEYINPUT101), .B(G93), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n526), .A2(new_n820), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n511), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n821), .B1(new_n501), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n819), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n551), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n550), .B1(new_n819), .B2(new_n823), .ZN(new_n826));
  AND2_X1   g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n818), .B(new_n827), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n829));
  INV_X1    g404(.A(G860), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(KEYINPUT39), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n829), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n824), .A2(new_n830), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT37), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n832), .A2(new_n834), .ZN(G145));
  XNOR2_X1  g410(.A(new_n761), .B(new_n712), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n475), .A2(G130), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n461), .A2(G118), .ZN(new_n838));
  OAI21_X1  g413(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g415(.A(new_n840), .B1(new_n485), .B2(G142), .ZN(new_n841));
  XOR2_X1   g416(.A(new_n841), .B(new_n619), .Z(new_n842));
  XNOR2_X1  g417(.A(new_n836), .B(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n496), .A2(new_n498), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n487), .A2(new_n491), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n738), .B(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n774), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n843), .B(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n626), .B(G160), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(G162), .ZN(new_n851));
  OR2_X1    g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(G37), .B1(new_n849), .B2(new_n851), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g430(.A(G299), .B(new_n601), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n856), .A2(KEYINPUT41), .ZN(new_n857));
  XNOR2_X1  g432(.A(G299), .B(new_n611), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT41), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n857), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n825), .A2(new_n826), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n615), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n864), .B1(new_n863), .B2(new_n858), .ZN(new_n865));
  XOR2_X1   g440(.A(G303), .B(KEYINPUT102), .Z(new_n866));
  XNOR2_X1  g441(.A(new_n798), .B(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(G290), .B(G305), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OR2_X1    g446(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n865), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n871), .A2(KEYINPUT104), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n865), .B2(new_n872), .ZN(new_n875));
  OAI21_X1  g450(.A(G868), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n878), .B(G868), .C1(new_n873), .C2(new_n875), .ZN(new_n879));
  OAI211_X1 g454(.A(new_n877), .B(new_n879), .C1(G868), .C2(new_n824), .ZN(G295));
  OAI211_X1 g455(.A(new_n877), .B(new_n879), .C1(G868), .C2(new_n824), .ZN(G331));
  NOR2_X1   g456(.A1(G286), .A2(new_n603), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT106), .ZN(new_n883));
  NAND2_X1  g458(.A1(G286), .A2(G171), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(G301), .A2(G168), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n886), .A2(KEYINPUT106), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n827), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n884), .A2(new_n883), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(new_n886), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n882), .A2(new_n883), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n890), .A2(new_n862), .A3(new_n891), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n888), .A2(new_n858), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n858), .A2(new_n859), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n856), .A2(KEYINPUT41), .ZN(new_n895));
  AOI22_X1  g470(.A1(new_n888), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n869), .B1(new_n893), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NOR3_X1   g473(.A1(new_n885), .A2(new_n887), .A3(new_n827), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n862), .B1(new_n890), .B2(new_n891), .ZN(new_n900));
  OAI22_X1  g475(.A1(new_n899), .A2(new_n900), .B1(new_n857), .B2(new_n860), .ZN(new_n901));
  INV_X1    g476(.A(new_n869), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n888), .A2(new_n858), .A3(new_n892), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n906), .A2(KEYINPUT108), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT44), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n907), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n901), .A2(new_n903), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n910), .B2(new_n869), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n909), .B1(new_n911), .B2(new_n904), .ZN(new_n912));
  OAI21_X1  g487(.A(KEYINPUT109), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n905), .A2(new_n907), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n904), .A3(new_n909), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT109), .ZN(new_n916));
  NAND4_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .A4(KEYINPUT44), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n913), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT107), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n919), .B1(new_n905), .B2(KEYINPUT43), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n911), .A2(KEYINPUT107), .A3(new_n906), .A4(new_n904), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n905), .A2(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT44), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n918), .A2(new_n925), .ZN(G397));
  INV_X1    g501(.A(KEYINPUT45), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n927), .B1(G164), .B2(G1384), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(G40), .ZN(new_n930));
  NOR3_X1   g505(.A1(new_n465), .A2(new_n469), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n738), .B(new_n741), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n933), .B1(new_n934), .B2(new_n761), .ZN(new_n935));
  INV_X1    g510(.A(G1996), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT46), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n940));
  XNOR2_X1  g515(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n761), .A2(G1996), .A3(new_n933), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n942), .B(KEYINPUT110), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n761), .A2(G1996), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n934), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n933), .B2(new_n945), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n775), .A2(new_n777), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n775), .A2(new_n777), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n933), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  NOR3_X1   g525(.A1(new_n932), .A2(G1986), .A3(G290), .ZN(new_n951));
  XNOR2_X1  g526(.A(new_n951), .B(KEYINPUT127), .ZN(new_n952));
  XNOR2_X1  g527(.A(new_n952), .B(KEYINPUT48), .ZN(new_n953));
  OAI21_X1  g528(.A(new_n941), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n946), .A2(new_n947), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n738), .A2(new_n741), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n932), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(G1986), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n950), .B1(new_n933), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT116), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT114), .ZN(new_n962));
  NAND2_X1  g537(.A1(G305), .A2(G1981), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT49), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n587), .A2(new_n787), .A3(new_n588), .A4(new_n589), .ZN(new_n965));
  AND3_X1   g540(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n963), .B2(new_n965), .ZN(new_n967));
  NOR2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g543(.A(KEYINPUT111), .B1(G164), .B2(G1384), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT111), .ZN(new_n970));
  INV_X1    g545(.A(G1384), .ZN(new_n971));
  INV_X1    g546(.A(new_n498), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n497), .B1(new_n462), .B2(new_n494), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n970), .B(new_n971), .C1(new_n974), .C2(new_n492), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n975), .A3(new_n931), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(G8), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n962), .B1(new_n968), .B2(new_n977), .ZN(new_n978));
  OAI22_X1  g553(.A1(new_n538), .A2(new_n583), .B1(new_n585), .B2(new_n508), .ZN(new_n979));
  AOI21_X1  g554(.A(new_n508), .B1(new_n502), .B2(new_n504), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n979), .A2(G651), .B1(G48), .B2(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n787), .B1(new_n981), .B2(new_n588), .ZN(new_n982));
  INV_X1    g557(.A(new_n965), .ZN(new_n983));
  OAI21_X1  g558(.A(KEYINPUT49), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n986), .A2(KEYINPUT114), .A3(G8), .A4(new_n976), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n978), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n969), .A2(new_n989), .A3(new_n975), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n931), .A2(new_n743), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n990), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n846), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n928), .A2(new_n994), .A3(new_n931), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n792), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n993), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g572(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n998));
  AOI21_X1  g573(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT112), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT112), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n506), .A2(new_n512), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n511), .A2(G62), .ZN(new_n1003));
  NAND2_X1  g578(.A1(G75), .A2(G543), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n501), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT55), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n1001), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1000), .A2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n997), .A2(new_n1011), .A3(G8), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n796), .A2(G1976), .A3(new_n797), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1013), .A2(G8), .A3(new_n976), .ZN(new_n1014));
  XOR2_X1   g589(.A(KEYINPUT113), .B(G1976), .Z(new_n1015));
  NAND3_X1  g590(.A1(new_n579), .A2(new_n581), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1014), .A2(KEYINPUT52), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n988), .A2(new_n1012), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1022), .B1(new_n997), .B2(G8), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT63), .ZN(new_n1024));
  INV_X1    g599(.A(G1966), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT45), .B1(new_n969), .B2(new_n975), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n994), .A2(new_n931), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1025), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2084), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n990), .A2(new_n1029), .A3(new_n931), .A4(new_n991), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1031), .A2(G8), .A3(G168), .ZN(new_n1032));
  NOR4_X1   g607(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .A4(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n846), .A2(new_n989), .A3(new_n971), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n931), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n969), .A2(new_n975), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1035), .B1(new_n1036), .B2(KEYINPUT50), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(new_n743), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n996), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1022), .B1(new_n1039), .B2(G8), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1021), .A2(new_n1040), .A3(new_n1032), .ZN(new_n1041));
  AOI21_X1  g616(.A(KEYINPUT63), .B1(new_n1041), .B2(KEYINPUT115), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT115), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1022), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1037), .A2(new_n743), .B1(new_n792), .B2(new_n995), .ZN(new_n1045));
  INV_X1    g620(.A(G8), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n976), .A2(G8), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1017), .B1(new_n1048), .B2(new_n1013), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1051), .A3(new_n1012), .A4(new_n988), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1043), .B1(new_n1052), .B2(new_n1032), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1033), .B1(new_n1042), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n988), .ZN(new_n1055));
  OR2_X1    g630(.A1(G288), .A2(G1976), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n965), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n1048), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1012), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1051), .A2(new_n1059), .A3(new_n988), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n961), .B1(new_n1054), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1021), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1032), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1063), .A2(KEYINPUT115), .A3(new_n1047), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1053), .A2(new_n1065), .A3(new_n1024), .ZN(new_n1066));
  INV_X1    g641(.A(new_n1033), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1061), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1068), .A2(KEYINPUT116), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1062), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1028), .A2(G168), .A3(new_n1030), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(G8), .ZN(new_n1073));
  AOI21_X1  g648(.A(G168), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT51), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT51), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1072), .A2(new_n1076), .A3(G8), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT62), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT62), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1075), .A2(new_n1080), .A3(new_n1077), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n990), .A2(new_n931), .A3(new_n991), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(KEYINPUT117), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n990), .A2(new_n1084), .A3(new_n931), .A4(new_n991), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT121), .B(G1961), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1085), .A3(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT53), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n995), .B2(G2078), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(G2078), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1087), .A2(new_n1089), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n603), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1052), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1079), .A2(new_n1081), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT124), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT124), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1079), .A2(new_n1081), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G1348), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1083), .A2(new_n1101), .A3(new_n1085), .ZN(new_n1102));
  OR2_X1    g677(.A1(new_n976), .A2(G2067), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1956), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n989), .B1(new_n969), .B2(new_n975), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1105), .B1(new_n1106), .B2(new_n1035), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n1108));
  AND3_X1   g683(.A1(new_n562), .A2(new_n1108), .A3(new_n566), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n562), .B2(new_n566), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AND3_X1   g686(.A1(new_n928), .A2(new_n994), .A3(new_n931), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1107), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1104), .A2(new_n611), .A3(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n567), .A2(KEYINPUT57), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT118), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n562), .A2(new_n1108), .A3(new_n566), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT118), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n970), .B1(new_n846), .B2(new_n971), .ZN(new_n1122));
  AOI211_X1 g697(.A(KEYINPUT111), .B(G1384), .C1(new_n844), .C2(new_n845), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT50), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  AND2_X1   g699(.A1(new_n1034), .A2(new_n931), .ZN(new_n1125));
  AOI21_X1  g700(.A(G1956), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1113), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n995), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1120), .B(new_n1121), .C1(new_n1126), .C2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n1103), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(new_n611), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n601), .A4(new_n1103), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT60), .ZN(new_n1134));
  AOI22_X1  g709(.A1(new_n1132), .A2(new_n1133), .B1(new_n1134), .B2(new_n1104), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1115), .A2(KEYINPUT61), .ZN(new_n1136));
  XOR2_X1   g711(.A(KEYINPUT58), .B(G1341), .Z(new_n1137));
  AOI22_X1  g712(.A1(new_n1112), .A2(new_n936), .B1(new_n976), .B2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(KEYINPUT59), .B1(new_n1138), .B2(new_n550), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n976), .A2(new_n1137), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(G1996), .B2(new_n995), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT59), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(new_n551), .A3(new_n1142), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1136), .A2(new_n1129), .B1(new_n1139), .B2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1145), .B1(new_n1126), .B2(new_n1128), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(new_n1115), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  AOI21_X1  g723(.A(KEYINPUT119), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n1150));
  AOI211_X1 g725(.A(new_n1150), .B(KEYINPUT61), .C1(new_n1146), .C2(new_n1115), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1144), .B1(new_n1149), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT120), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1135), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1144), .B(KEYINPUT120), .C1(new_n1149), .C2(new_n1151), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1130), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1093), .A2(new_n603), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n928), .A2(new_n931), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(KEYINPUT122), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1159), .A2(new_n994), .A3(new_n1091), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1160), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1161), .A2(KEYINPUT123), .A3(G171), .ZN(new_n1162));
  AOI21_X1  g737(.A(KEYINPUT123), .B1(new_n1161), .B2(G171), .ZN(new_n1163));
  OAI211_X1 g738(.A(KEYINPUT54), .B(new_n1157), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1094), .B1(new_n603), .B2(new_n1161), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT54), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1052), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1164), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n1100), .B1(new_n1156), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g745(.A(KEYINPUT125), .B(new_n960), .C1(new_n1071), .C2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1130), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1104), .A2(new_n1134), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1115), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1139), .A2(new_n1143), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1177), .A2(new_n1178), .ZN(new_n1179));
  NOR3_X1   g754(.A1(new_n1126), .A2(new_n1145), .A3(new_n1128), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1111), .B1(new_n1107), .B2(new_n1114), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1148), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1182), .A2(new_n1150), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1147), .A2(KEYINPUT119), .A3(new_n1148), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1179), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1176), .B1(new_n1185), .B2(KEYINPUT120), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1155), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1173), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1169), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND4_X1  g765(.A1(new_n1190), .A2(new_n1100), .A3(new_n1062), .A4(new_n1070), .ZN(new_n1191));
  AOI21_X1  g766(.A(KEYINPUT125), .B1(new_n1191), .B2(new_n960), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n958), .B1(new_n1172), .B2(new_n1192), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g768(.A1(G227), .A2(new_n459), .ZN(new_n1195));
  NAND3_X1  g769(.A1(new_n686), .A2(new_n648), .A3(new_n1195), .ZN(new_n1196));
  AOI21_X1  g770(.A(new_n1196), .B1(new_n852), .B2(new_n853), .ZN(new_n1197));
  NAND2_X1  g771(.A1(new_n1197), .A2(new_n923), .ZN(G225));
  INV_X1    g772(.A(G225), .ZN(G308));
endmodule


