//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 0 0 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:44 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n684, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n920, new_n921, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n973, new_n974,
    new_n975;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  INV_X1    g001(.A(G228gat), .ZN(new_n203));
  INV_X1    g002(.A(G233gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(KEYINPUT74), .B(G155gat), .Z(new_n206));
  INV_X1    g005(.A(G162gat), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT2), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G141gat), .B(G148gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(G141gat), .ZN(new_n212));
  OR3_X1    g011(.A1(new_n212), .A2(KEYINPUT73), .A3(G148gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n208), .A2(new_n210), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g014(.A(new_n211), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT72), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n209), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(new_n209), .B2(new_n217), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n216), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n214), .A2(new_n215), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT29), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT70), .ZN(new_n225));
  XNOR2_X1  g024(.A(G211gat), .B(G218gat), .ZN(new_n226));
  XNOR2_X1  g025(.A(G197gat), .B(G204gat), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT22), .ZN(new_n228));
  INV_X1    g027(.A(G211gat), .ZN(new_n229));
  INV_X1    g028(.A(G218gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n228), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(new_n227), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  AOI21_X1  g032(.A(new_n226), .B1(new_n231), .B2(new_n227), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n225), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n227), .A2(new_n231), .ZN(new_n236));
  INV_X1    g035(.A(new_n226), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n238), .A2(KEYINPUT70), .A3(new_n232), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n224), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n214), .A2(new_n221), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT29), .B1(new_n238), .B2(new_n232), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n215), .B1(new_n244), .B2(KEYINPUT81), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n223), .B1(new_n233), .B2(new_n234), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT81), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n243), .B1(new_n245), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g048(.A(new_n205), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n205), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n243), .B2(KEYINPUT3), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n244), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n240), .B1(new_n223), .B2(new_n222), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR3_X1   g055(.A1(new_n250), .A2(new_n256), .A3(G22gat), .ZN(new_n257));
  INV_X1    g056(.A(G22gat), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n214), .A2(new_n221), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT3), .B1(new_n246), .B2(new_n247), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n244), .A2(KEYINPUT81), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n251), .B1(new_n262), .B2(new_n255), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n242), .A2(new_n253), .A3(new_n252), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n258), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT80), .B(KEYINPUT31), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n257), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(G22gat), .B1(new_n250), .B2(new_n256), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n263), .A2(new_n258), .A3(new_n264), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G78gat), .B(G106gat), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n272), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n267), .B1(new_n257), .B2(new_n265), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n269), .A2(new_n270), .A3(new_n266), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(KEYINPUT82), .B(G50gat), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NOR3_X1   g078(.A1(new_n273), .A2(new_n277), .A3(new_n279), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n272), .B1(new_n268), .B2(new_n271), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n274), .A3(new_n276), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n202), .B1(new_n280), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(G227gat), .A2(G233gat), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  XNOR2_X1  g088(.A(G127gat), .B(G134gat), .ZN(new_n290));
  XNOR2_X1  g089(.A(new_n289), .B(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(G169gat), .A2(G176gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(G169gat), .A2(G176gat), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n293), .B1(KEYINPUT23), .B2(new_n294), .ZN(new_n295));
  AND2_X1   g094(.A1(new_n293), .A2(KEYINPUT23), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  NOR2_X1   g096(.A1(new_n297), .A2(KEYINPUT25), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  INV_X1    g098(.A(G190gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n301), .B(KEYINPUT65), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(G183gat), .A2(G190gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT24), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n304), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n302), .A2(new_n305), .A3(new_n308), .A4(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n298), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n307), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n301), .A2(new_n303), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n313), .B1(new_n314), .B2(new_n308), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n297), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n311), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n294), .ZN(new_n319));
  NOR3_X1   g118(.A1(new_n319), .A2(new_n293), .A3(KEYINPUT26), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n293), .A2(KEYINPUT26), .ZN(new_n321));
  INV_X1    g120(.A(new_n306), .ZN(new_n322));
  NOR3_X1   g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT27), .B(G183gat), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(KEYINPUT68), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n326), .A2(KEYINPUT28), .A3(new_n300), .A4(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n325), .A2(new_n300), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT67), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT28), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(new_n332), .A3(new_n300), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n324), .B1(new_n328), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n292), .B1(new_n318), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n297), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n315), .A2(new_n312), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n339), .A2(KEYINPUT25), .B1(new_n298), .B2(new_n310), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n334), .A2(new_n328), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n323), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n340), .A2(new_n342), .A3(new_n291), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n285), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT32), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n336), .A2(new_n285), .A3(new_n343), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(KEYINPUT34), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT34), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n336), .A2(new_n343), .A3(new_n349), .A4(new_n285), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g150(.A(G15gat), .B(G43gat), .Z(new_n352));
  XNOR2_X1  g151(.A(G71gat), .B(G99gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n352), .B(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n285), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n318), .A2(new_n335), .A3(new_n292), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n291), .B1(new_n340), .B2(new_n342), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n356), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n360), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n354), .B1(new_n344), .B2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n364), .A2(new_n348), .A3(new_n350), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n346), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(new_n365), .A3(new_n346), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n367), .A2(KEYINPUT86), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT86), .ZN(new_n370));
  INV_X1    g169(.A(new_n368), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n366), .ZN(new_n372));
  INV_X1    g171(.A(G226gat), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n340), .B(new_n342), .C1(new_n373), .C2(new_n204), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n318), .A2(new_n335), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n373), .A2(new_n204), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n376), .A2(KEYINPUT29), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n374), .B(new_n240), .C1(new_n375), .C2(new_n377), .ZN(new_n378));
  NOR3_X1   g177(.A1(new_n318), .A2(new_n335), .A3(new_n376), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n340), .B2(new_n342), .ZN(new_n380));
  OAI21_X1  g179(.A(new_n241), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n378), .A2(new_n381), .A3(KEYINPUT30), .A4(new_n385), .ZN(new_n388));
  AND2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n378), .A2(new_n381), .A3(new_n385), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT71), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT30), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT71), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n378), .A2(new_n381), .A3(new_n393), .A4(new_n385), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n391), .A2(new_n392), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n369), .A2(new_n372), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n399));
  AND3_X1   g198(.A1(new_n399), .A2(new_n292), .A3(new_n222), .ZN(new_n400));
  NAND2_X1  g199(.A1(G225gat), .A2(G233gat), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(KEYINPUT75), .B(KEYINPUT5), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n259), .A2(KEYINPUT4), .A3(new_n291), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n291), .A2(new_n214), .A3(new_n221), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n405), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n406), .B1(new_n405), .B2(new_n409), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n403), .B(new_n404), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n399), .A2(new_n292), .A3(new_n222), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n414), .A2(new_n409), .A3(new_n405), .A4(new_n401), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n243), .A2(new_n292), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n407), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n404), .B1(new_n417), .B2(new_n402), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n415), .A2(KEYINPUT76), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(KEYINPUT76), .B1(new_n415), .B2(new_n418), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT77), .B(KEYINPUT0), .Z(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT78), .ZN(new_n423));
  XNOR2_X1  g222(.A(G1gat), .B(G29gat), .ZN(new_n424));
  XNOR2_X1  g223(.A(new_n423), .B(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G57gat), .B(G85gat), .ZN(new_n426));
  XOR2_X1   g225(.A(new_n425), .B(new_n426), .Z(new_n427));
  INV_X1    g226(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n421), .A2(KEYINPUT6), .A3(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n429), .A2(KEYINPUT85), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n421), .A2(new_n428), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT6), .ZN(new_n432));
  OAI211_X1 g231(.A(new_n413), .B(new_n427), .C1(new_n419), .C2(new_n420), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT85), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n430), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OR3_X1    g236(.A1(new_n284), .A2(new_n398), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n367), .A2(new_n368), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n279), .B1(new_n273), .B2(new_n277), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n281), .A2(new_n278), .A3(new_n282), .ZN(new_n441));
  AOI21_X1  g240(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n435), .A2(new_n397), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n202), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(KEYINPUT85), .B1(new_n434), .B2(new_n429), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n386), .B1(new_n382), .B2(KEYINPUT37), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n378), .A2(new_n381), .A3(KEYINPUT83), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n450), .B(KEYINPUT37), .C1(KEYINPUT83), .C2(new_n378), .ZN(new_n451));
  XOR2_X1   g250(.A(KEYINPUT84), .B(KEYINPUT38), .Z(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n452), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n382), .A2(KEYINPUT37), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n454), .B1(new_n455), .B2(new_n448), .ZN(new_n456));
  AND2_X1   g255(.A1(new_n391), .A2(new_n394), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n453), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n447), .A2(new_n430), .A3(new_n458), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n416), .A2(new_n407), .A3(new_n401), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n405), .A2(new_n409), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT79), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n400), .B1(new_n462), .B2(new_n410), .ZN(new_n463));
  OAI211_X1 g262(.A(KEYINPUT39), .B(new_n460), .C1(new_n463), .C2(new_n401), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n414), .B1(new_n411), .B2(new_n412), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT39), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n465), .A2(new_n466), .A3(new_n402), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n427), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT40), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g269(.A1(new_n464), .A2(KEYINPUT40), .A3(new_n427), .A4(new_n467), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n470), .A2(new_n396), .A3(new_n431), .A4(new_n471), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n472), .B1(new_n280), .B2(new_n283), .ZN(new_n473));
  OR2_X1    g272(.A1(new_n459), .A2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n443), .A2(new_n441), .A3(new_n440), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT36), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n439), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n371), .A2(new_n366), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(KEYINPUT36), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AND2_X1   g279(.A1(new_n475), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g280(.A1(new_n438), .A2(new_n446), .B1(new_n474), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G113gat), .B(G141gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(G169gat), .B(G197gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  XNOR2_X1  g284(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XNOR2_X1  g286(.A(new_n487), .B(KEYINPUT12), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT17), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g292(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g294(.A1(G43gat), .A2(G50gat), .ZN(new_n496));
  NOR2_X1   g295(.A1(G43gat), .A2(G50gat), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT15), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n491), .A2(new_n492), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n495), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT15), .ZN(new_n502));
  INV_X1    g301(.A(G43gat), .ZN(new_n503));
  INV_X1    g302(.A(G50gat), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  XNOR2_X1  g304(.A(KEYINPUT89), .B(G43gat), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n504), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n501), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g309(.A(KEYINPUT88), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n510), .A2(new_n511), .A3(new_n493), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n498), .B1(new_n512), .B2(new_n500), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n489), .B1(new_n508), .B2(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(G43gat), .B(G50gat), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n499), .B1(new_n515), .B2(KEYINPUT15), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n503), .A2(KEYINPUT89), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT89), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G43gat), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n517), .A2(new_n519), .A3(new_n504), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n522), .A3(new_n495), .ZN(new_n523));
  NOR2_X1   g322(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n494), .A2(new_n509), .B1(new_n524), .B2(new_n492), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n499), .B1(new_n525), .B2(new_n511), .ZN(new_n526));
  OAI211_X1 g325(.A(new_n523), .B(KEYINPUT17), .C1(new_n498), .C2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G1gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT16), .ZN(new_n529));
  INV_X1    g328(.A(G15gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(G22gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n258), .A2(G15gat), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g332(.A(G1gat), .B1(new_n531), .B2(new_n532), .ZN(new_n534));
  OAI21_X1  g333(.A(G8gat), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n529), .A2(new_n531), .A3(new_n532), .ZN(new_n536));
  INV_X1    g335(.A(G8gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(G15gat), .B(G22gat), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n536), .B(new_n537), .C1(G1gat), .C2(new_n538), .ZN(new_n539));
  AND2_X1   g338(.A1(new_n535), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n514), .A2(new_n527), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(G229gat), .A2(G233gat), .ZN(new_n542));
  OAI22_X1  g341(.A1(new_n526), .A2(new_n498), .B1(new_n501), .B2(new_n507), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n535), .A2(new_n539), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n543), .A2(KEYINPUT90), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT90), .B1(new_n543), .B2(new_n544), .ZN(new_n546));
  OAI211_X1 g345(.A(new_n541), .B(new_n542), .C1(new_n545), .C2(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT91), .B(KEYINPUT18), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n508), .A2(new_n513), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(new_n540), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n551), .B1(new_n545), .B2(new_n546), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n542), .B(KEYINPUT13), .Z(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT90), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n550), .B2(new_n540), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n543), .A2(KEYINPUT90), .A3(new_n544), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n558), .A2(KEYINPUT18), .A3(new_n542), .A4(new_n541), .ZN(new_n559));
  AND4_X1   g358(.A1(new_n488), .A2(new_n549), .A3(new_n554), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n554), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT93), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n559), .A2(new_n554), .A3(KEYINPUT93), .ZN(new_n564));
  AOI21_X1  g363(.A(KEYINPUT92), .B1(new_n547), .B2(new_n548), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n547), .A2(KEYINPUT92), .A3(new_n548), .ZN(new_n567));
  NAND4_X1  g366(.A1(new_n563), .A2(new_n564), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n488), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n560), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G57gat), .B(G64gat), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(G71gat), .A2(G78gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(G71gat), .A2(G78gat), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT9), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n572), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n574), .B(new_n573), .C1(new_n571), .C2(new_n576), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT21), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G231gat), .A2(G233gat), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G127gat), .B(G155gat), .ZN(new_n585));
  XOR2_X1   g384(.A(new_n585), .B(KEYINPUT20), .Z(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n584), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G183gat), .B(G211gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n584), .B(new_n586), .ZN(new_n591));
  INV_X1    g390(.A(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n540), .B1(new_n581), .B2(new_n580), .ZN(new_n595));
  XOR2_X1   g394(.A(KEYINPUT94), .B(KEYINPUT19), .Z(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n594), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(G120gat), .B(G148gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(G176gat), .B(G204gat), .ZN(new_n600));
  XOR2_X1   g399(.A(new_n599), .B(new_n600), .Z(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(KEYINPUT102), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G99gat), .A2(G106gat), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT97), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT97), .A2(G99gat), .A3(G106gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n607), .A2(KEYINPUT8), .A3(new_n608), .ZN(new_n609));
  OAI21_X1  g408(.A(G92gat), .B1(KEYINPUT7), .B2(G85gat), .ZN(new_n610));
  AND2_X1   g409(.A1(KEYINPUT7), .A2(G85gat), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(G92gat), .ZN(new_n613));
  AND3_X1   g412(.A1(new_n613), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n614));
  OAI21_X1  g413(.A(new_n609), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G99gat), .B(G106gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n609), .B(new_n616), .C1(new_n612), .C2(new_n614), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n618), .A2(KEYINPUT98), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n615), .A2(new_n621), .A3(new_n617), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n620), .A2(new_n580), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  INV_X1    g423(.A(new_n580), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n625), .A2(new_n618), .A3(new_n619), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n623), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n620), .A2(new_n622), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(KEYINPUT10), .A3(new_n625), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n604), .B1(new_n627), .B2(new_n629), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n603), .B1(new_n623), .B2(new_n626), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n602), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n627), .A2(KEYINPUT100), .A3(new_n629), .ZN(new_n633));
  AOI21_X1  g432(.A(KEYINPUT100), .B1(new_n627), .B2(new_n629), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n633), .A2(new_n634), .A3(new_n604), .ZN(new_n635));
  INV_X1    g434(.A(new_n601), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n636), .B1(new_n631), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n637), .B2(new_n631), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n632), .B1(new_n635), .B2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n628), .A2(new_n543), .ZN(new_n642));
  NAND2_X1  g441(.A1(G232gat), .A2(G233gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT95), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n514), .A2(new_n527), .ZN(new_n647));
  OAI211_X1 g446(.A(new_n642), .B(new_n646), .C1(new_n647), .C2(new_n628), .ZN(new_n648));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT99), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OR2_X1    g450(.A1(new_n647), .A2(new_n628), .ZN(new_n652));
  INV_X1    g451(.A(new_n650), .ZN(new_n653));
  NAND4_X1  g452(.A1(new_n652), .A2(new_n653), .A3(new_n646), .A4(new_n642), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n645), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(KEYINPUT96), .ZN(new_n656));
  XOR2_X1   g455(.A(G134gat), .B(G162gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  AND3_X1   g457(.A1(new_n651), .A2(new_n654), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n658), .B1(new_n651), .B2(new_n654), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n598), .A2(new_n641), .A3(new_n661), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n482), .A2(new_n570), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n664), .A2(new_n435), .ZN(new_n665));
  XNOR2_X1  g464(.A(KEYINPUT103), .B(G1gat), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n665), .B(new_n666), .ZN(G1324gat));
  XNOR2_X1  g466(.A(KEYINPUT104), .B(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n663), .A2(new_n396), .ZN(new_n669));
  XOR2_X1   g468(.A(KEYINPUT16), .B(G8gat), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n668), .B1(new_n669), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(KEYINPUT105), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n537), .B1(new_n663), .B2(new_n396), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n674), .A2(KEYINPUT106), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(KEYINPUT106), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n669), .A2(new_n671), .ZN(new_n677));
  AOI22_X1  g476(.A1(new_n675), .A2(new_n676), .B1(KEYINPUT42), .B2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n673), .A2(new_n678), .ZN(G1325gat));
  OAI21_X1  g478(.A(G15gat), .B1(new_n664), .B2(new_n480), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n369), .A2(new_n372), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n663), .A2(new_n530), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(G1326gat));
  NAND2_X1  g482(.A1(new_n440), .A2(new_n441), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n663), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT43), .B(G22gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1327gat));
  OAI211_X1 g487(.A(new_n475), .B(new_n480), .C1(new_n459), .C2(new_n473), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n284), .A2(new_n398), .A3(new_n437), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n689), .B1(new_n690), .B2(new_n445), .ZN(new_n691));
  INV_X1    g490(.A(new_n598), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n641), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(new_n661), .ZN(new_n694));
  AOI21_X1  g493(.A(KEYINPUT93), .B1(new_n559), .B2(new_n554), .ZN(new_n695));
  AND3_X1   g494(.A1(new_n547), .A2(KEYINPUT92), .A3(new_n548), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n695), .A2(new_n696), .A3(new_n565), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n488), .B1(new_n697), .B2(new_n564), .ZN(new_n698));
  OAI211_X1 g497(.A(new_n691), .B(new_n694), .C1(new_n698), .C2(new_n560), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n699), .A2(G29gat), .A3(new_n435), .ZN(new_n700));
  XOR2_X1   g499(.A(new_n700), .B(KEYINPUT45), .Z(new_n701));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n482), .B2(new_n661), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n659), .A2(new_n660), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n691), .A2(KEYINPUT44), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT107), .B1(new_n698), .B2(new_n560), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n570), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n693), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n435), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n701), .A2(new_n713), .ZN(G1328gat));
  NOR3_X1   g513(.A1(new_n699), .A2(G36gat), .A3(new_n397), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT46), .ZN(new_n716));
  OAI21_X1  g515(.A(KEYINPUT108), .B1(new_n712), .B2(new_n397), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(G36gat), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n712), .A2(KEYINPUT108), .A3(new_n397), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n716), .B1(new_n718), .B2(new_n719), .ZN(G1329gat));
  INV_X1    g519(.A(new_n480), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n703), .A2(new_n721), .A3(new_n705), .A4(new_n711), .ZN(new_n722));
  INV_X1    g521(.A(new_n506), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n681), .ZN(new_n725));
  NOR3_X1   g524(.A1(new_n699), .A2(new_n723), .A3(new_n725), .ZN(new_n726));
  NOR2_X1   g525(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(KEYINPUT109), .A2(KEYINPUT47), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n729), .B(new_n730), .ZN(G1330gat));
  OAI21_X1  g530(.A(new_n504), .B1(new_n699), .B2(new_n684), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n685), .A2(G50gat), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n712), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT110), .B(KEYINPUT48), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1331gat));
  NAND4_X1  g535(.A1(new_n710), .A2(new_n598), .A3(new_n661), .A4(new_n640), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n482), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n740), .A2(new_n435), .ZN(new_n741));
  XOR2_X1   g540(.A(new_n741), .B(G57gat), .Z(G1332gat));
  OAI22_X1  g541(.A1(new_n740), .A2(new_n397), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n743));
  XNOR2_X1  g542(.A(new_n738), .B(KEYINPUT111), .ZN(new_n744));
  XNOR2_X1  g543(.A(KEYINPUT49), .B(G64gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n744), .A2(new_n396), .A3(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1333gat));
  OAI21_X1  g546(.A(G71gat), .B1(new_n740), .B2(new_n480), .ZN(new_n748));
  INV_X1    g547(.A(G71gat), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n744), .A2(new_n749), .A3(new_n681), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(new_n750), .A3(KEYINPUT50), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(G1334gat));
  NAND2_X1  g554(.A1(new_n744), .A2(new_n685), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g556(.A1(new_n710), .A2(new_n692), .ZN(new_n758));
  INV_X1    g557(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n640), .ZN(new_n760));
  XOR2_X1   g559(.A(new_n760), .B(KEYINPUT112), .Z(new_n761));
  NAND2_X1  g560(.A1(new_n706), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g561(.A(G85gat), .B1(new_n762), .B2(new_n435), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n435), .A2(G85gat), .A3(new_n641), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n691), .A2(new_n704), .A3(new_n759), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT51), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n691), .A2(KEYINPUT51), .A3(new_n704), .A4(new_n759), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n764), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n763), .A2(new_n771), .ZN(G1336gat));
  NAND3_X1  g571(.A1(new_n767), .A2(KEYINPUT113), .A3(new_n769), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT113), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n765), .A2(new_n774), .A3(new_n766), .ZN(new_n775));
  NOR3_X1   g574(.A1(new_n397), .A2(G92gat), .A3(new_n641), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(KEYINPUT114), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n773), .A2(new_n779), .A3(new_n775), .A4(new_n776), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n703), .A2(new_n396), .A3(new_n705), .A4(new_n761), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(G92gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n778), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(KEYINPUT52), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n776), .B1(new_n768), .B2(new_n770), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT52), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n785), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n784), .A2(new_n787), .ZN(G1337gat));
  NAND4_X1  g587(.A1(new_n703), .A2(new_n721), .A3(new_n705), .A4(new_n761), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(G99gat), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n725), .A2(G99gat), .A3(new_n641), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n791), .B1(new_n768), .B2(new_n770), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT115), .ZN(G1338gat));
  NAND4_X1  g593(.A1(new_n703), .A2(new_n685), .A3(new_n705), .A4(new_n761), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G106gat), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n684), .A2(G106gat), .A3(new_n641), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n797), .B1(new_n768), .B2(new_n770), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT53), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n773), .A2(new_n775), .A3(new_n797), .ZN(new_n801));
  AND2_X1   g600(.A1(new_n801), .A2(new_n796), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n800), .B1(new_n802), .B2(new_n799), .ZN(G1339gat));
  INV_X1    g602(.A(KEYINPUT55), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n627), .A2(new_n629), .A3(new_n604), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT54), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n627), .A2(new_n629), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT100), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n604), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n627), .A2(KEYINPUT100), .A3(new_n629), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n601), .B1(new_n630), .B2(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n804), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  OR2_X1    g614(.A1(new_n635), .A2(new_n639), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT55), .B(new_n813), .C1(new_n635), .C2(new_n806), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n707), .A2(new_n709), .A3(new_n818), .ZN(new_n819));
  INV_X1    g618(.A(new_n561), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n549), .A2(new_n488), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n558), .A2(new_n541), .ZN(new_n822));
  OAI22_X1  g621(.A1(new_n822), .A2(new_n542), .B1(new_n552), .B2(new_n553), .ZN(new_n823));
  AOI22_X1  g622(.A1(new_n820), .A2(new_n821), .B1(new_n823), .B2(new_n487), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n824), .A2(new_n640), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n704), .B1(new_n819), .B2(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n823), .A2(new_n487), .ZN(new_n828));
  NOR3_X1   g627(.A1(new_n661), .A2(new_n828), .A3(new_n560), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n818), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n704), .A2(new_n824), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT116), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n692), .B1(new_n826), .B2(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n662), .B1(new_n707), .B2(new_n709), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI211_X1 g636(.A(new_n435), .B(new_n685), .C1(new_n835), .C2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n397), .A3(new_n681), .ZN(new_n839));
  NOR3_X1   g638(.A1(new_n839), .A2(new_n286), .A3(new_n570), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n838), .A2(new_n478), .ZN(new_n841));
  INV_X1    g640(.A(new_n710), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n397), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n840), .B1(new_n286), .B2(new_n843), .ZN(G1340gat));
  NOR3_X1   g643(.A1(new_n839), .A2(new_n287), .A3(new_n641), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n841), .A2(new_n397), .A3(new_n640), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n845), .B1(new_n287), .B2(new_n846), .ZN(G1341gat));
  NOR2_X1   g646(.A1(new_n692), .A2(G127gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n841), .A2(new_n397), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(G127gat), .B1(new_n839), .B2(new_n692), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1342gat));
  NAND2_X1  g650(.A1(new_n397), .A2(new_n704), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(G134gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n841), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g653(.A(new_n854), .B(KEYINPUT56), .Z(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n839), .B2(new_n661), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1343gat));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n825), .B1(new_n831), .B2(new_n570), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n661), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n860), .A2(new_n833), .A3(new_n830), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n836), .B1(new_n861), .B2(new_n692), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT57), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n684), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n858), .B1(new_n862), .B2(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n830), .A2(new_n833), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n598), .B1(new_n867), .B2(new_n860), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT117), .B(new_n864), .C1(new_n868), .C2(new_n836), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n684), .B1(new_n835), .B2(new_n837), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n866), .B(new_n869), .C1(new_n870), .C2(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n480), .A2(new_n429), .A3(new_n434), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(new_n396), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(G141gat), .B1(new_n874), .B2(new_n570), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT58), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n870), .A2(new_n873), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n570), .A2(G141gat), .ZN(new_n878));
  XNOR2_X1  g677(.A(new_n878), .B(KEYINPUT119), .ZN(new_n879));
  AND2_X1   g678(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n875), .A2(new_n876), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n874), .A2(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n871), .A2(KEYINPUT118), .A3(new_n873), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n884), .A2(new_n842), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n880), .B1(new_n886), .B2(G141gat), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(new_n876), .ZN(G1344gat));
  INV_X1    g687(.A(KEYINPUT120), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n871), .A2(KEYINPUT118), .A3(new_n873), .ZN(new_n890));
  AOI21_X1  g689(.A(KEYINPUT118), .B1(new_n871), .B2(new_n873), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n890), .A2(new_n891), .A3(new_n641), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(G148gat), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n884), .A2(new_n640), .A3(new_n885), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n896), .A2(KEYINPUT120), .A3(new_n893), .A4(G148gat), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n662), .A2(new_n698), .A3(new_n560), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT121), .ZN(new_n899));
  OR2_X1    g698(.A1(new_n898), .A2(KEYINPUT121), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n818), .A2(new_n829), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n860), .A2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT122), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n692), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n860), .A2(new_n903), .A3(new_n901), .ZN(new_n905));
  OAI211_X1 g704(.A(new_n899), .B(new_n900), .C1(new_n904), .C2(new_n905), .ZN(new_n906));
  AOI21_X1  g705(.A(KEYINPUT57), .B1(new_n906), .B2(new_n685), .ZN(new_n907));
  INV_X1    g706(.A(new_n870), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n863), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n640), .B(new_n873), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G148gat), .ZN(new_n912));
  OAI21_X1  g711(.A(KEYINPUT59), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n895), .A2(new_n897), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n877), .A2(new_n912), .A3(new_n640), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n914), .A2(new_n915), .ZN(G1345gat));
  NAND3_X1  g715(.A1(new_n877), .A2(new_n206), .A3(new_n598), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n890), .A2(new_n891), .A3(new_n692), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n917), .B1(new_n918), .B2(new_n206), .ZN(G1346gat));
  OR4_X1    g718(.A1(G162gat), .A2(new_n908), .A3(new_n852), .A4(new_n872), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n890), .A2(new_n891), .A3(new_n661), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n920), .B1(new_n921), .B2(new_n207), .ZN(G1347gat));
  NAND2_X1  g721(.A1(new_n835), .A2(new_n837), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n397), .B1(new_n429), .B2(new_n434), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  NOR3_X1   g724(.A1(new_n725), .A2(new_n685), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(G169gat), .B1(new_n927), .B2(new_n570), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n923), .A2(new_n435), .ZN(new_n929));
  AND2_X1   g728(.A1(new_n442), .A2(new_n396), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OR2_X1    g730(.A1(new_n710), .A2(G169gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n928), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  XOR2_X1   g732(.A(new_n933), .B(KEYINPUT123), .Z(G1348gat));
  OAI21_X1  g733(.A(G176gat), .B1(new_n927), .B2(new_n641), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n641), .A2(G176gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n931), .B2(new_n936), .ZN(G1349gat));
  INV_X1    g736(.A(new_n927), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n299), .B1(new_n938), .B2(new_n598), .ZN(new_n939));
  INV_X1    g738(.A(new_n931), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n598), .A2(new_n326), .A3(new_n327), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  XOR2_X1   g741(.A(new_n942), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g742(.A1(new_n940), .A2(new_n300), .A3(new_n704), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT124), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n300), .B1(new_n938), .B2(new_n704), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XOR2_X1   g747(.A(new_n948), .B(KEYINPUT126), .Z(new_n949));
  NOR2_X1   g748(.A1(new_n946), .A2(new_n947), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT125), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n945), .B1(new_n949), .B2(new_n951), .ZN(G1351gat));
  AND4_X1   g751(.A1(new_n396), .A2(new_n929), .A3(new_n685), .A4(new_n480), .ZN(new_n953));
  AOI21_X1  g752(.A(G197gat), .B1(new_n953), .B2(new_n842), .ZN(new_n954));
  OR2_X1    g753(.A1(new_n907), .A2(new_n909), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n721), .A2(new_n925), .ZN(new_n956));
  AND2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(G197gat), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n570), .A2(new_n958), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n954), .B1(new_n957), .B2(new_n959), .ZN(G1352gat));
  AOI21_X1  g759(.A(G204gat), .B1(KEYINPUT127), .B2(KEYINPUT62), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n953), .A2(new_n640), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g761(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n963));
  XNOR2_X1  g762(.A(new_n962), .B(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n955), .A2(new_n640), .A3(new_n956), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(G204gat), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1353gat));
  NAND3_X1  g766(.A1(new_n953), .A2(new_n229), .A3(new_n598), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n955), .A2(new_n598), .A3(new_n956), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n969), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n970));
  AOI21_X1  g769(.A(KEYINPUT63), .B1(new_n969), .B2(G211gat), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n968), .B1(new_n970), .B2(new_n971), .ZN(G1354gat));
  NAND3_X1  g771(.A1(new_n953), .A2(new_n230), .A3(new_n704), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n957), .A2(new_n704), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n973), .B1(new_n975), .B2(new_n230), .ZN(G1355gat));
endmodule


