//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:52 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252, new_n1253;
  INV_X1    g0000(.A(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n203), .A2(G50), .A3(G58), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  INV_X1    g0006(.A(G87), .ZN(new_n207));
  INV_X1    g0007(.A(G250), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G68), .B2(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G107), .ZN(new_n213));
  INV_X1    g0013(.A(G264), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  INV_X1    g0018(.A(G244), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n202), .C2(new_n219), .ZN(new_n220));
  INV_X1    g0020(.A(G58), .ZN(new_n221));
  INV_X1    g0021(.A(G232), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n206), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n224), .B(KEYINPUT1), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n206), .A2(G13), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  AOI211_X1 g0027(.A(new_n208), .B(new_n227), .C1(new_n210), .C2(new_n214), .ZN(new_n228));
  OR2_X1    g0028(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n228), .A2(KEYINPUT0), .ZN(new_n230));
  NAND2_X1  g0030(.A1(G1), .A2(G13), .ZN(new_n231));
  INV_X1    g0031(.A(G20), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g0034(.A(G50), .B1(G58), .B2(G68), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n229), .B(new_n230), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT64), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n225), .A2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n222), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G238), .B(G244), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G250), .B(G257), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n214), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(G270), .ZN(new_n245));
  XOR2_X1   g0045(.A(new_n242), .B(new_n245), .Z(G358));
  NOR2_X1   g0046(.A1(new_n201), .A2(new_n202), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n203), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(KEYINPUT65), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(G107), .B(G116), .Z(new_n253));
  XNOR2_X1  g0053(.A(G87), .B(G97), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n252), .B(new_n255), .ZN(G351));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(KEYINPUT3), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT3), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1698), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G222), .ZN(new_n263));
  NAND2_X1  g0063(.A1(G223), .A2(G1698), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT67), .ZN(new_n266));
  XNOR2_X1  g0066(.A(KEYINPUT3), .B(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(new_n202), .ZN(new_n268));
  OR3_X1    g0068(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n231), .B1(G33), .B2(G41), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n265), .B2(new_n268), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n269), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G1), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(G274), .ZN(new_n274));
  OR2_X1    g0074(.A1(KEYINPUT66), .A2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(KEYINPUT66), .A2(G41), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n274), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(G33), .A2(G41), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n281), .A2(G1), .A3(G13), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n273), .B1(G41), .B2(G45), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G226), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n272), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n290), .A2(G58), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT8), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n291), .B(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n232), .A2(G33), .ZN(new_n294));
  INV_X1    g0094(.A(G150), .ZN(new_n295));
  NOR2_X1   g0095(.A1(G20), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI22_X1  g0097(.A1(new_n293), .A2(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(G58), .A2(G68), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n232), .B1(new_n301), .B2(new_n217), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT70), .ZN(new_n303));
  OAI221_X1 g0103(.A(KEYINPUT69), .B1(new_n295), .B2(new_n297), .C1(new_n293), .C2(new_n294), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(new_n231), .ZN(new_n307));
  INV_X1    g0107(.A(G13), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n308), .A2(G1), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G20), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n305), .A2(new_n307), .B1(new_n217), .B2(new_n311), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n307), .B1(new_n273), .B2(G20), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G50), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n312), .A2(KEYINPUT9), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n289), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT10), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT9), .B1(new_n312), .B2(new_n314), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n287), .A2(G200), .ZN(new_n320));
  NAND4_X1  g0120(.A1(new_n316), .A2(new_n317), .A3(new_n319), .A4(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n289), .A2(new_n315), .A3(new_n320), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT10), .B1(new_n322), .B2(new_n318), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n312), .A2(new_n314), .ZN(new_n325));
  INV_X1    g0125(.A(G169), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n287), .A2(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n325), .B(new_n327), .C1(G179), .C2(new_n287), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT14), .ZN(new_n329));
  NOR2_X1   g0129(.A1(G226), .A2(G1698), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(new_n222), .B2(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n267), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n279), .B1(new_n334), .B2(new_n270), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT13), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n285), .A2(G238), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n331), .A2(new_n267), .B1(G33), .B2(G97), .ZN(new_n339));
  OAI211_X1 g0139(.A(new_n280), .B(new_n337), .C1(new_n282), .C2(new_n339), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(KEYINPUT13), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n338), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n329), .B1(new_n342), .B2(G169), .ZN(new_n343));
  AOI211_X1 g0143(.A(KEYINPUT14), .B(new_n326), .C1(new_n338), .C2(new_n341), .ZN(new_n344));
  INV_X1    g0144(.A(G179), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n343), .A2(new_n344), .A3(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n309), .A2(G20), .A3(new_n201), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n348), .B(KEYINPUT12), .ZN(new_n349));
  INV_X1    g0149(.A(new_n313), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n201), .B2(new_n350), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n297), .A2(new_n217), .B1(new_n232), .B2(G68), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n294), .A2(new_n202), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n307), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(KEYINPUT11), .ZN(new_n356));
  AOI21_X1  g0156(.A(new_n351), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n347), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(G238), .A2(G1698), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n267), .B(new_n359), .C1(new_n222), .C2(G1698), .ZN(new_n360));
  OAI211_X1 g0160(.A(new_n360), .B(new_n270), .C1(G107), .C2(new_n267), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n280), .C1(new_n219), .C2(new_n284), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G200), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT8), .B(G58), .Z(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n296), .B1(G20), .B2(G77), .ZN(new_n365));
  XNOR2_X1  g0165(.A(KEYINPUT15), .B(G87), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n365), .B1(new_n366), .B2(new_n294), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n367), .A2(new_n307), .B1(new_n202), .B2(new_n311), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n368), .B1(new_n202), .B2(new_n350), .ZN(new_n369));
  OAI221_X1 g0169(.A(new_n363), .B1(new_n288), .B2(new_n362), .C1(new_n369), .C2(KEYINPUT71), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n369), .A2(KEYINPUT71), .ZN(new_n371));
  OR2_X1    g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  OR2_X1    g0172(.A1(new_n362), .A2(G179), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n362), .A2(new_n326), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n369), .A3(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n372), .A2(KEYINPUT72), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n324), .A2(new_n328), .A3(new_n358), .A4(new_n376), .ZN(new_n377));
  OR2_X1    g0177(.A1(new_n293), .A2(new_n313), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n293), .A2(new_n310), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n307), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n221), .A2(new_n201), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n301), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n296), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT7), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n267), .B2(G20), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n261), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n386), .B1(new_n390), .B2(G68), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n382), .B1(new_n391), .B2(KEYINPUT16), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT16), .ZN(new_n393));
  OAI21_X1  g0193(.A(KEYINPUT75), .B1(new_n259), .B2(G33), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT75), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(new_n257), .A3(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n394), .A2(new_n396), .A3(new_n260), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n232), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n201), .B1(new_n398), .B2(new_n388), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n393), .B1(new_n399), .B2(new_n386), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n381), .B1(new_n392), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT77), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n402), .B1(new_n279), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n282), .A2(G232), .A3(new_n283), .ZN(new_n405));
  AOI21_X1  g0205(.A(G45), .B1(new_n275), .B2(new_n276), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n405), .B(KEYINPUT77), .C1(new_n406), .C2(new_n274), .ZN(new_n407));
  OR2_X1    g0207(.A1(G223), .A2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n218), .A2(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n258), .A2(new_n408), .A3(new_n260), .A4(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(new_n270), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n404), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G200), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT76), .B1(new_n412), .B2(new_n270), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT76), .ZN(new_n418));
  AOI211_X1 g0218(.A(new_n418), .B(new_n282), .C1(new_n410), .C2(new_n411), .ZN(new_n419));
  OAI211_X1 g0219(.A(new_n404), .B(new_n407), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n416), .B1(new_n420), .B2(G190), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n401), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n401), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n425));
  AND2_X1   g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n342), .A2(G200), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT73), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n338), .A2(new_n341), .A3(G190), .ZN(new_n430));
  AND2_X1   g0230(.A1(new_n430), .A2(new_n357), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n342), .A2(KEYINPUT73), .A3(G200), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n429), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(KEYINPUT74), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT74), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n429), .A2(new_n431), .A3(new_n435), .A4(new_n432), .ZN(new_n436));
  NOR2_X1   g0236(.A1(new_n417), .A2(new_n419), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n404), .A2(new_n407), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n345), .B1(new_n326), .B2(new_n414), .ZN(new_n440));
  INV_X1    g0240(.A(new_n400), .ZN(new_n441));
  AOI21_X1  g0241(.A(KEYINPUT7), .B1(new_n261), .B2(new_n232), .ZN(new_n442));
  AOI211_X1 g0242(.A(new_n387), .B(G20), .C1(new_n258), .C2(new_n260), .ZN(new_n443));
  OAI21_X1  g0243(.A(G68), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n386), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n444), .A2(KEYINPUT16), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n446), .A2(new_n307), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n380), .B1(new_n441), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n440), .A2(new_n448), .A3(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT18), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n414), .A2(new_n326), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n420), .B2(G179), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n450), .B1(new_n401), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n426), .A2(new_n434), .A3(new_n436), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(KEYINPUT72), .B1(new_n372), .B2(new_n375), .ZN(new_n456));
  OR3_X1    g0256(.A1(new_n377), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n219), .A2(G1698), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n267), .B(new_n458), .C1(G238), .C2(G1698), .ZN(new_n459));
  NAND2_X1  g0259(.A1(G33), .A2(G116), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n282), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n273), .A2(G45), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n462), .A2(G274), .ZN(new_n463));
  AOI211_X1 g0263(.A(new_n270), .B(new_n463), .C1(new_n208), .C2(new_n462), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(new_n415), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n267), .A2(new_n232), .A3(G68), .ZN(new_n467));
  NOR2_X1   g0267(.A1(G97), .A2(G107), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(new_n207), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n333), .A2(new_n232), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n469), .A2(KEYINPUT19), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n333), .A2(G20), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n467), .B(new_n471), .C1(KEYINPUT19), .C2(new_n472), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n473), .A2(new_n307), .B1(new_n366), .B2(new_n311), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n273), .A2(G33), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n382), .A2(new_n310), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G87), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n474), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n466), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n465), .A2(G190), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n474), .B1(new_n366), .B2(new_n476), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n465), .A2(new_n345), .ZN(new_n484));
  OAI211_X1 g0284(.A(new_n483), .B(new_n484), .C1(G169), .C2(new_n465), .ZN(new_n485));
  AND2_X1   g0285(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n258), .A2(new_n260), .A3(G244), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(G1698), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n267), .A2(G244), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(G33), .A2(G283), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n489), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n267), .A2(G250), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n262), .B1(new_n494), .B2(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n270), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT5), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n273), .B(G45), .C1(new_n497), .C2(G41), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n275), .A2(new_n497), .A3(new_n276), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n270), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(G257), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n499), .A2(new_n500), .A3(G274), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n504), .A2(new_n288), .ZN(new_n505));
  AOI21_X1  g0305(.A(new_n505), .B1(G200), .B2(new_n504), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n310), .A2(G97), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(new_n477), .B2(G97), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT78), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT6), .ZN(new_n511));
  AND2_X1   g0311(.A1(G97), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n511), .B1(new_n512), .B2(new_n468), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n232), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n297), .A2(new_n202), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n510), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n516), .ZN(new_n518));
  AND3_X1   g0318(.A1(new_n213), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  XNOR2_X1  g0319(.A(G97), .B(G107), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(new_n511), .ZN(new_n521));
  OAI211_X1 g0321(.A(KEYINPUT78), .B(new_n518), .C1(new_n521), .C2(new_n232), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n517), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n213), .B1(new_n398), .B2(new_n388), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n307), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(KEYINPUT79), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT79), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n527), .B(new_n307), .C1(new_n523), .C2(new_n524), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n509), .B1(new_n526), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n506), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n504), .A2(new_n326), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n531), .B1(G179), .B2(new_n504), .ZN(new_n532));
  NOR3_X1   g0332(.A1(new_n529), .A2(KEYINPUT80), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT80), .ZN(new_n534));
  INV_X1    g0334(.A(new_n528), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n398), .A2(new_n388), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(G107), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n537), .A2(new_n517), .A3(new_n522), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n527), .B1(new_n538), .B2(new_n307), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n508), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  AND2_X1   g0340(.A1(new_n504), .A2(new_n326), .ZN(new_n541));
  NOR2_X1   g0341(.A1(new_n504), .A2(G179), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n534), .B1(new_n540), .B2(new_n543), .ZN(new_n544));
  OAI211_X1 g0344(.A(new_n486), .B(new_n530), .C1(new_n533), .C2(new_n544), .ZN(new_n545));
  XOR2_X1   g0345(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n546));
  NAND4_X1  g0346(.A1(new_n546), .A2(new_n232), .A3(G87), .A4(new_n267), .ZN(new_n547));
  INV_X1    g0347(.A(G116), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n294), .A2(new_n548), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT23), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(G20), .B2(new_n213), .ZN(new_n551));
  NOR3_X1   g0351(.A1(new_n232), .A2(KEYINPUT23), .A3(G107), .ZN(new_n552));
  NOR3_X1   g0352(.A1(new_n549), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n258), .A2(new_n260), .A3(new_n232), .A4(G87), .ZN(new_n554));
  XNOR2_X1  g0354(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n547), .A2(new_n553), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT24), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n547), .A2(new_n553), .A3(new_n559), .A4(new_n556), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n382), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n476), .A2(new_n213), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT25), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n310), .B2(G107), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n564), .A2(KEYINPUT84), .ZN(new_n565));
  NOR3_X1   g0365(.A1(new_n561), .A2(new_n562), .A3(new_n565), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n311), .A2(KEYINPUT25), .A3(new_n213), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n567), .A2(KEYINPUT84), .A3(new_n564), .ZN(new_n568));
  AND2_X1   g0368(.A1(KEYINPUT66), .A2(G41), .ZN(new_n569));
  NOR2_X1   g0369(.A1(KEYINPUT66), .A2(G41), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(KEYINPUT5), .ZN(new_n571));
  OAI211_X1 g0371(.A(G264), .B(new_n282), .C1(new_n571), .C2(new_n498), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(new_n503), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n208), .A2(new_n262), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n210), .A2(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n267), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n282), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n573), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(G200), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(G190), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n566), .A2(new_n568), .A3(new_n581), .A4(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n558), .A2(new_n560), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n307), .ZN(new_n585));
  INV_X1    g0385(.A(new_n562), .ZN(new_n586));
  INV_X1    g0386(.A(new_n565), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n585), .A2(new_n568), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  OAI21_X1  g0388(.A(KEYINPUT85), .B1(new_n579), .B2(new_n326), .ZN(new_n589));
  INV_X1    g0389(.A(new_n578), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n590), .A2(G179), .A3(new_n503), .A4(new_n572), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT86), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n579), .A2(KEYINPUT86), .A3(G179), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT85), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n595), .B(G169), .C1(new_n573), .C2(new_n578), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n589), .A2(new_n593), .A3(new_n594), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n588), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n583), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n311), .A2(new_n548), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n382), .A2(new_n310), .A3(G116), .A4(new_n475), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n306), .A2(new_n231), .B1(G20), .B2(new_n548), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n492), .B(new_n232), .C1(G33), .C2(new_n209), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n602), .A2(KEYINPUT20), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(KEYINPUT20), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n600), .B(new_n601), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  OAI211_X1 g0406(.A(G270), .B(new_n282), .C1(new_n571), .C2(new_n498), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT81), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n501), .A2(KEYINPUT81), .A3(G270), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n270), .B1(new_n267), .B2(G303), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n262), .A2(G257), .ZN(new_n613));
  NAND2_X1  g0413(.A1(G264), .A2(G1698), .ZN(new_n614));
  AND4_X1   g0414(.A1(new_n258), .A2(new_n260), .A3(new_n613), .A4(new_n614), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n503), .B1(new_n612), .B2(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n611), .A2(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n618), .A2(new_n345), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n616), .B1(new_n609), .B2(new_n610), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT21), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n620), .A2(new_n621), .A3(new_n326), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n606), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT82), .ZN(new_n624));
  INV_X1    g0424(.A(new_n606), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n620), .A2(new_n625), .A3(new_n326), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n624), .B1(new_n626), .B2(KEYINPUT21), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n618), .A2(G169), .A3(new_n606), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(KEYINPUT82), .A3(new_n621), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n620), .A2(G190), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n625), .C1(new_n415), .C2(new_n620), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n623), .A2(new_n627), .A3(new_n629), .A4(new_n631), .ZN(new_n632));
  NOR4_X1   g0432(.A1(new_n457), .A2(new_n545), .A3(new_n599), .A4(new_n632), .ZN(G372));
  NOR3_X1   g0433(.A1(new_n377), .A2(new_n455), .A3(new_n456), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT80), .B1(new_n529), .B2(new_n532), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n540), .A2(new_n534), .A3(new_n543), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n636), .A3(new_n486), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(KEYINPUT26), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n540), .A2(new_n543), .A3(new_n639), .A4(new_n482), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n485), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n598), .A2(new_n623), .A3(new_n627), .A4(new_n629), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n583), .ZN(new_n644));
  OAI211_X1 g0444(.A(new_n638), .B(new_n642), .C1(new_n545), .C2(new_n644), .ZN(new_n645));
  AND2_X1   g0445(.A1(new_n634), .A2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(KEYINPUT18), .B1(new_n440), .B2(new_n448), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n401), .A2(new_n452), .A3(new_n450), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n375), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n433), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n358), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n649), .B1(new_n652), .B2(new_n426), .ZN(new_n653));
  INV_X1    g0453(.A(new_n324), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n328), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n646), .A2(new_n655), .ZN(G369));
  NAND3_X1  g0456(.A1(new_n623), .A2(new_n627), .A3(new_n629), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT87), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n309), .A2(new_n232), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(G213), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n660), .B2(new_n661), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n659), .A2(KEYINPUT87), .A3(KEYINPUT27), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n662), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n669), .A2(new_n625), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n657), .A2(new_n670), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n671), .A2(KEYINPUT88), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n672), .B(new_n673), .C1(new_n632), .C2(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(G330), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n669), .B1(new_n566), .B2(new_n568), .ZN(new_n677));
  OAI22_X1  g0477(.A1(new_n599), .A2(new_n677), .B1(new_n598), .B2(new_n669), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n643), .A2(new_n583), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n669), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT89), .ZN(G399));
  NOR2_X1   g0483(.A1(new_n569), .A2(new_n570), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n227), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(G1), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n468), .A2(new_n207), .A3(new_n548), .ZN(new_n688));
  OAI22_X1  g0488(.A1(new_n687), .A2(new_n688), .B1(new_n235), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n689), .B(KEYINPUT28), .ZN(new_n690));
  INV_X1    g0490(.A(new_n482), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n635), .A2(new_n636), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(new_n530), .A3(new_n583), .A4(new_n643), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n635), .A2(new_n636), .A3(new_n639), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n691), .A2(new_n529), .A3(new_n532), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n485), .B1(new_n696), .B2(new_n639), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n669), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n698), .A2(KEYINPUT29), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT29), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n645), .A2(new_n700), .A3(new_n669), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  AOI22_X1  g0502(.A1(new_n635), .A2(new_n636), .B1(new_n529), .B2(new_n506), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n599), .A2(new_n632), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n703), .A2(new_n704), .A3(new_n486), .A4(new_n669), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n579), .A2(new_n496), .A3(new_n502), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT90), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n620), .A2(new_n707), .A3(G179), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  AOI21_X1  g0509(.A(new_n707), .B1(new_n620), .B2(G179), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n465), .B(new_n706), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(KEYINPUT91), .A2(KEYINPUT30), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(KEYINPUT90), .B1(new_n618), .B2(new_n345), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n708), .ZN(new_n715));
  INV_X1    g0515(.A(new_n712), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n715), .A2(new_n465), .A3(new_n716), .A4(new_n706), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT92), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n465), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n461), .A2(new_n464), .A3(KEYINPUT92), .ZN(new_n720));
  NOR3_X1   g0520(.A1(new_n719), .A2(new_n620), .A3(new_n720), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n721), .A2(new_n345), .A3(new_n504), .A4(new_n580), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n713), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n668), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT31), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n705), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n728), .A2(G330), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n702), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n690), .B1(new_n731), .B2(G1), .ZN(G364));
  OR2_X1    g0532(.A1(new_n674), .A2(G330), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n308), .A2(G20), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G45), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n686), .A2(G1), .A3(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(new_n736), .B(KEYINPUT93), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n733), .A2(new_n675), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT94), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n742), .A2(G20), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n674), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g0545(.A(new_n231), .B1(G20), .B2(new_n326), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT98), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(new_n415), .B2(G179), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n345), .A2(KEYINPUT98), .A3(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n232), .A2(G190), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n749), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G283), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n261), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NOR3_X1   g0554(.A1(new_n288), .A2(G179), .A3(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n232), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G294), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n345), .A2(G200), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n751), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G179), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n751), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AOI22_X1  g0564(.A1(G311), .A2(new_n761), .B1(new_n764), .B2(G329), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n232), .A2(new_n345), .A3(new_n415), .ZN(new_n766));
  OR2_X1    g0566(.A1(new_n766), .A2(KEYINPUT97), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(KEYINPUT97), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n767), .A2(G190), .A3(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(G326), .ZN(new_n770));
  OAI211_X1 g0570(.A(new_n758), .B(new_n765), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n288), .A3(new_n768), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(KEYINPUT33), .B(G317), .ZN(new_n774));
  AOI211_X1 g0574(.A(new_n754), .B(new_n771), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(G303), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n232), .A2(new_n288), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n749), .A2(new_n777), .A3(new_n750), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT96), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n777), .A2(new_n780), .A3(new_n759), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n777), .B2(new_n759), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n775), .B1(new_n776), .B2(new_n778), .C1(new_n779), .C2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n756), .A2(new_n209), .ZN(new_n785));
  INV_X1    g0585(.A(new_n752), .ZN(new_n786));
  AOI22_X1  g0586(.A1(new_n786), .A2(G107), .B1(new_n761), .B2(G77), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n772), .B2(new_n201), .ZN(new_n788));
  INV_X1    g0588(.A(new_n769), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n785), .B(new_n788), .C1(G50), .C2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n778), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G87), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT32), .ZN(new_n793));
  AOI21_X1  g0593(.A(new_n793), .B1(new_n764), .B2(G159), .ZN(new_n794));
  INV_X1    g0594(.A(G159), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n763), .A2(KEYINPUT32), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n783), .ZN(new_n797));
  AOI211_X1 g0597(.A(new_n794), .B(new_n796), .C1(new_n797), .C2(G58), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n790), .A2(new_n267), .A3(new_n792), .A4(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n747), .B1(new_n784), .B2(new_n799), .ZN(new_n800));
  OR3_X1    g0600(.A1(new_n745), .A2(new_n738), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n227), .A2(new_n261), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G355), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n252), .A2(new_n278), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n227), .A2(new_n267), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(G45), .B2(new_n235), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n803), .B1(G116), .B2(new_n226), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n743), .A2(new_n746), .ZN(new_n808));
  XNOR2_X1  g0608(.A(new_n808), .B(KEYINPUT95), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n739), .B1(new_n801), .B2(new_n810), .ZN(G396));
  AOI21_X1  g0611(.A(new_n785), .B1(G116), .B2(new_n761), .ZN(new_n812));
  INV_X1    g0612(.A(G311), .ZN(new_n813));
  OAI211_X1 g0613(.A(new_n812), .B(new_n261), .C1(new_n813), .C2(new_n763), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n789), .A2(G303), .B1(G107), .B2(new_n791), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n815), .B1(new_n207), .B2(new_n752), .C1(new_n753), .C2(new_n772), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n814), .B(new_n816), .C1(G294), .C2(new_n797), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT99), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n773), .A2(G150), .B1(new_n797), .B2(G143), .ZN(new_n819));
  INV_X1    g0619(.A(G137), .ZN(new_n820));
  OAI221_X1 g0620(.A(new_n819), .B1(new_n820), .B2(new_n769), .C1(new_n795), .C2(new_n760), .ZN(new_n821));
  XOR2_X1   g0621(.A(new_n821), .B(KEYINPUT34), .Z(new_n822));
  AOI22_X1  g0622(.A1(G58), .A2(new_n757), .B1(new_n791), .B2(G50), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n786), .A2(G68), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n823), .A2(new_n267), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g0625(.A(new_n825), .B1(G132), .B2(new_n764), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT100), .Z(new_n827));
  NOR2_X1   g0627(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n746), .B1(new_n818), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n746), .A2(new_n740), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n737), .C1(G77), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n369), .A2(new_n668), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n833), .B1(new_n370), .B2(new_n371), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n834), .A2(new_n375), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n650), .A2(new_n669), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n838), .A2(new_n742), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n680), .A2(new_n703), .A3(new_n486), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n641), .B1(new_n637), .B2(KEYINPUT26), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n668), .B(new_n837), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n838), .B1(new_n645), .B2(new_n669), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n845), .A2(new_n729), .ZN(new_n846));
  XOR2_X1   g0646(.A(new_n846), .B(KEYINPUT101), .Z(new_n847));
  AOI21_X1  g0647(.A(new_n737), .B1(new_n845), .B2(new_n729), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n840), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(G384));
  AOI21_X1  g0650(.A(new_n457), .B1(new_n699), .B2(new_n701), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n851), .A2(new_n655), .ZN(new_n852));
  INV_X1    g0652(.A(new_n666), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n392), .B1(KEYINPUT16), .B2(new_n391), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n854), .A2(new_n380), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n424), .A2(new_n425), .ZN(new_n856));
  OAI211_X1 g0656(.A(new_n853), .B(new_n855), .C1(new_n649), .C2(new_n856), .ZN(new_n857));
  AOI22_X1  g0657(.A1(new_n380), .A2(new_n854), .B1(new_n452), .B2(new_n666), .ZN(new_n858));
  INV_X1    g0658(.A(new_n422), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT37), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n440), .A2(new_n448), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n448), .A2(new_n853), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n422), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n860), .B1(KEYINPUT37), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT38), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n434), .A2(new_n436), .A3(new_n347), .ZN(new_n869));
  NOR2_X1   g0669(.A1(new_n357), .A2(new_n669), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n358), .A2(new_n433), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g0674(.A(new_n836), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n868), .B(new_n874), .C1(new_n843), .C2(new_n875), .ZN(new_n876));
  XOR2_X1   g0676(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  XNOR2_X1  g0678(.A(new_n863), .B(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n862), .B1(new_n426), .B2(new_n454), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n877), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n867), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g0684(.A1(new_n358), .A2(new_n668), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n866), .A2(KEYINPUT39), .A3(new_n867), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n649), .A2(new_n666), .ZN(new_n888));
  AND3_X1   g0688(.A1(new_n876), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XOR2_X1   g0689(.A(new_n852), .B(new_n889), .Z(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n837), .B1(new_n871), .B2(new_n873), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n728), .A2(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n857), .A2(new_n864), .A3(KEYINPUT38), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n865), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n891), .B1(new_n893), .B2(new_n895), .ZN(new_n896));
  NAND4_X1  g0696(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n728), .A4(new_n892), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n634), .A2(new_n728), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n898), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n890), .B(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n273), .B2(new_n734), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT35), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n234), .B1(new_n521), .B2(new_n904), .ZN(new_n905));
  OAI211_X1 g0705(.A(new_n905), .B(G116), .C1(new_n904), .C2(new_n521), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT36), .ZN(new_n907));
  OAI21_X1  g0707(.A(G77), .B1(new_n221), .B2(new_n201), .ZN(new_n908));
  OAI22_X1  g0708(.A1(new_n908), .A2(new_n235), .B1(G50), .B2(new_n201), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n909), .A2(G1), .A3(new_n308), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n903), .A2(new_n907), .A3(new_n910), .ZN(G367));
  NAND2_X1  g0711(.A1(new_n479), .A2(new_n668), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n486), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n485), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n703), .B1(new_n529), .B2(new_n669), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n540), .A2(new_n543), .A3(new_n668), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(new_n919));
  AND2_X1   g0719(.A1(new_n657), .A2(new_n669), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n920), .A2(new_n598), .A3(new_n583), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g0722(.A(new_n922), .B(KEYINPUT42), .Z(new_n923));
  NAND3_X1  g0723(.A1(new_n918), .A2(new_n588), .A3(new_n597), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n668), .B1(new_n924), .B2(new_n692), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n915), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n679), .A2(new_n919), .ZN(new_n927));
  AND2_X1   g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n926), .A2(new_n927), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n928), .B2(new_n929), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n685), .B(KEYINPUT41), .ZN(new_n934));
  INV_X1    g0734(.A(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT103), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n918), .A2(new_n936), .A3(new_n681), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n936), .B1(new_n918), .B2(new_n681), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT45), .ZN(new_n939));
  OR3_X1    g0739(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n916), .A2(new_n680), .A3(new_n669), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT44), .Z(new_n942));
  OAI21_X1  g0742(.A(new_n939), .B1(new_n937), .B2(new_n938), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(new_n679), .ZN(new_n945));
  OR2_X1    g0745(.A1(new_n678), .A2(new_n920), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n921), .ZN(new_n947));
  OR2_X1    g0747(.A1(new_n947), .A2(KEYINPUT104), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(KEYINPUT104), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n676), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n675), .B1(KEYINPUT104), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n731), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n953), .A2(KEYINPUT105), .ZN(new_n954));
  INV_X1    g0754(.A(KEYINPUT105), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n731), .B2(new_n952), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n945), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n935), .B1(new_n957), .B2(new_n731), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n735), .A2(G1), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n932), .B(new_n933), .C1(new_n958), .C2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n757), .A2(G68), .ZN(new_n961));
  OAI221_X1 g0761(.A(new_n961), .B1(new_n217), .B2(new_n760), .C1(new_n202), .C2(new_n752), .ZN(new_n962));
  AOI211_X1 g0762(.A(new_n261), .B(new_n962), .C1(G137), .C2(new_n764), .ZN(new_n963));
  AOI22_X1  g0763(.A1(new_n789), .A2(G143), .B1(G58), .B2(new_n791), .ZN(new_n964));
  AND2_X1   g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n965), .B1(new_n295), .B2(new_n783), .C1(new_n795), .C2(new_n772), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n783), .A2(new_n776), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n791), .A2(G116), .ZN(new_n968));
  XNOR2_X1  g0768(.A(KEYINPUT106), .B(KEYINPUT46), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n968), .A2(new_n969), .B1(new_n970), .B2(new_n763), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n267), .B(new_n971), .C1(G97), .C2(new_n786), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT46), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n968), .B1(KEYINPUT106), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n761), .A2(G283), .ZN(new_n975));
  OAI22_X1  g0775(.A1(new_n769), .A2(new_n813), .B1(new_n756), .B2(new_n213), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n976), .B1(G294), .B2(new_n773), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n972), .A2(new_n974), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n966), .B1(new_n967), .B2(new_n978), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT47), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n746), .ZN(new_n981));
  INV_X1    g0781(.A(new_n805), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n809), .B1(new_n226), .B2(new_n366), .C1(new_n245), .C2(new_n982), .ZN(new_n983));
  OR2_X1    g0783(.A1(new_n914), .A2(new_n744), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n981), .A2(new_n737), .A3(new_n983), .A4(new_n984), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT107), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n960), .A2(new_n986), .ZN(G387));
  NAND2_X1  g0787(.A1(new_n952), .A2(new_n959), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n730), .B1(new_n950), .B2(new_n951), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n989), .A2(KEYINPUT111), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(KEYINPUT111), .ZN(new_n991));
  NAND4_X1  g0791(.A1(new_n990), .A2(new_n685), .A3(new_n953), .A4(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n772), .A2(new_n293), .B1(new_n778), .B2(new_n202), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n756), .A2(new_n366), .B1(new_n295), .B2(new_n763), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n752), .A2(new_n209), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n267), .B1(new_n760), .B2(new_n201), .ZN(new_n996));
  NOR4_X1   g0796(.A1(new_n993), .A2(new_n994), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n217), .B2(new_n783), .C1(new_n795), .C2(new_n769), .ZN(new_n998));
  OAI22_X1  g0798(.A1(new_n783), .A2(new_n970), .B1(new_n776), .B2(new_n760), .ZN(new_n999));
  XOR2_X1   g0799(.A(new_n999), .B(KEYINPUT108), .Z(new_n1000));
  OAI221_X1 g0800(.A(new_n1000), .B1(new_n813), .B2(new_n772), .C1(new_n779), .C2(new_n769), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT109), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT48), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G283), .A2(new_n757), .B1(new_n791), .B2(G294), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n786), .A2(G116), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n764), .A2(G326), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n261), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1005), .A2(KEYINPUT49), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n998), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n746), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n678), .A2(new_n744), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n982), .B1(new_n242), .B2(G45), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n688), .B2(new_n802), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n364), .A2(new_n217), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT50), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1017), .A2(G45), .A3(new_n247), .A4(new_n688), .ZN(new_n1018));
  OAI22_X1  g0818(.A1(new_n1015), .A2(new_n1018), .B1(G107), .B2(new_n226), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n738), .B1(new_n1019), .B2(new_n809), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1012), .A2(new_n1013), .A3(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n988), .B(new_n992), .C1(new_n1022), .C2(new_n1023), .ZN(G393));
  NAND2_X1  g0824(.A1(new_n945), .A2(new_n959), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n919), .A2(new_n743), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT112), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n809), .B1(new_n209), .B2(new_n226), .C1(new_n255), .C2(new_n982), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n778), .A2(new_n201), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n769), .A2(new_n295), .B1(new_n783), .B2(new_n795), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT51), .Z(new_n1031));
  AOI211_X1 g0831(.A(new_n1029), .B(new_n1031), .C1(G50), .C2(new_n773), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n757), .A2(G77), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n786), .A2(G87), .B1(new_n764), .B2(G143), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n261), .B1(new_n761), .B2(new_n364), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n769), .A2(new_n970), .B1(new_n783), .B2(new_n813), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT52), .Z(new_n1038));
  AOI211_X1 g0838(.A(new_n267), .B(new_n1038), .C1(G303), .C2(new_n773), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n764), .A2(G322), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n791), .A2(G283), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n786), .A2(G107), .B1(new_n761), .B2(G294), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n756), .A2(new_n548), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1036), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n738), .B1(new_n1045), .B2(new_n746), .ZN(new_n1046));
  NAND3_X1  g0846(.A1(new_n1027), .A2(new_n1028), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1025), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n945), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n953), .ZN(new_n1050));
  AND2_X1   g0850(.A1(new_n1050), .A2(new_n957), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1048), .B1(new_n1051), .B2(new_n685), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(G390));
  NAND4_X1  g0853(.A1(new_n728), .A2(G330), .A3(new_n838), .A4(new_n874), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1054), .ZN(new_n1055));
  NOR3_X1   g0855(.A1(new_n894), .A2(new_n865), .A3(new_n883), .ZN(new_n1056));
  AOI21_X1  g0856(.A(KEYINPUT39), .B1(new_n881), .B2(new_n867), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n874), .B1(new_n843), .B2(new_n875), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n885), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1058), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n882), .A2(new_n1060), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n669), .B(new_n835), .C1(new_n695), .C2(new_n697), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n836), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1062), .B1(new_n1064), .B2(new_n874), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1055), .B1(new_n1061), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n884), .A2(new_n886), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n874), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n645), .A2(new_n669), .A3(new_n838), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1068), .B1(new_n1069), .B2(new_n836), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n1067), .B1(new_n1070), .B2(new_n885), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1068), .B1(new_n1063), .B2(new_n836), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1071), .B(new_n1054), .C1(new_n1072), .C2(new_n1062), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1066), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G330), .ZN(new_n1075));
  AND3_X1   g0875(.A1(new_n723), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n1076));
  AOI21_X1  g0876(.A(KEYINPUT31), .B1(new_n723), .B2(new_n668), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1075), .B1(new_n1078), .B2(new_n705), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n874), .B1(new_n1079), .B2(new_n838), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n1080), .A2(new_n1055), .B1(new_n875), .B2(new_n843), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1068), .B1(new_n729), .B2(new_n837), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1082), .A2(new_n836), .A3(new_n1063), .A4(new_n1054), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n634), .A2(G330), .A3(new_n728), .ZN(new_n1085));
  NOR3_X1   g0885(.A1(new_n851), .A2(new_n1085), .A3(new_n655), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1074), .A2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1066), .A2(new_n1073), .A3(new_n1086), .A4(new_n1084), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1088), .A2(new_n685), .A3(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1066), .A2(new_n1073), .A3(new_n959), .ZN(new_n1091));
  INV_X1    g0891(.A(G125), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n763), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n773), .A2(G137), .B1(G50), .B2(new_n786), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n760), .B2(new_n1095), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n1093), .B(new_n1096), .C1(G128), .C2(new_n789), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n757), .A2(G159), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n791), .A2(G150), .ZN(new_n1099));
  XOR2_X1   g0899(.A(KEYINPUT113), .B(KEYINPUT53), .Z(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n267), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1102), .B1(G132), .B2(new_n797), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n1097), .A2(new_n1098), .A3(new_n1101), .A4(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1033), .B1(new_n209), .B2(new_n760), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n267), .B(new_n1105), .C1(G294), .C2(new_n764), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n773), .A2(G107), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n792), .B1(new_n769), .B2(new_n753), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G116), .B2(new_n797), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1106), .A2(new_n824), .A3(new_n1107), .A4(new_n1109), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n747), .B1(new_n1104), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n738), .B(new_n1111), .C1(new_n293), .C2(new_n830), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n1058), .B2(new_n742), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1090), .A2(new_n1091), .A3(new_n1113), .ZN(G378));
  NOR2_X1   g0914(.A1(new_n831), .A2(G50), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(G33), .A2(G41), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT114), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1117), .B(new_n217), .C1(new_n267), .C2(new_n684), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n778), .A2(new_n1095), .ZN(new_n1119));
  INV_X1    g0919(.A(G132), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n772), .A2(new_n1120), .B1(new_n820), .B2(new_n760), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1119), .B(new_n1121), .C1(G128), .C2(new_n797), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1122), .B1(new_n1092), .B2(new_n769), .C1(new_n295), .C2(new_n756), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT59), .Z(new_n1124));
  AOI21_X1  g0924(.A(new_n1117), .B1(G124), .B2(new_n764), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n1124), .B(new_n1125), .C1(new_n795), .C2(new_n752), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n961), .B1(new_n769), .B2(new_n548), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT115), .Z(new_n1128));
  NOR2_X1   g0928(.A1(new_n684), .A2(new_n267), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n366), .B2(new_n760), .C1(new_n772), .C2(new_n209), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n752), .A2(new_n221), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n783), .A2(new_n213), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n763), .A2(new_n753), .ZN(new_n1133));
  NOR4_X1   g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1128), .B(new_n1134), .C1(new_n202), .C2(new_n778), .ZN(new_n1135));
  XOR2_X1   g0935(.A(new_n1135), .B(KEYINPUT116), .Z(new_n1136));
  INV_X1    g0936(.A(KEYINPUT58), .ZN(new_n1137));
  OR2_X1    g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1139));
  AND4_X1   g0939(.A1(new_n1118), .A2(new_n1126), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n737), .B1(new_n1140), .B2(new_n747), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n324), .A2(new_n328), .ZN(new_n1142));
  XOR2_X1   g0942(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n324), .A2(new_n328), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n325), .A2(new_n853), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1144), .A2(new_n325), .A3(new_n853), .A4(new_n1146), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1115), .B(new_n1141), .C1(new_n1151), .C2(new_n741), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n896), .A2(G330), .A3(new_n897), .ZN(new_n1153));
  AND2_X1   g0953(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g0955(.A1(new_n1151), .A2(G330), .A3(new_n896), .A4(new_n897), .ZN(new_n1156));
  AND3_X1   g0956(.A1(new_n1155), .A2(new_n889), .A3(new_n1156), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n889), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1158));
  NOR2_X1   g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1152), .B1(new_n1159), .B2(new_n959), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1089), .A2(new_n1086), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1161), .A2(KEYINPUT57), .A3(new_n1159), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n685), .ZN(new_n1163));
  AOI21_X1  g0963(.A(KEYINPUT57), .B1(new_n1161), .B2(new_n1159), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1160), .B1(new_n1163), .B2(new_n1164), .ZN(G375));
  AOI22_X1  g0965(.A1(new_n789), .A2(G294), .B1(G107), .B2(new_n761), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1166), .B1(new_n548), .B2(new_n772), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT118), .Z(new_n1168));
  OAI22_X1  g0968(.A1(new_n366), .A2(new_n756), .B1(new_n778), .B2(new_n209), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n752), .A2(new_n202), .B1(new_n763), .B2(new_n776), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n261), .B1(new_n783), .B2(new_n753), .ZN(new_n1171));
  NOR4_X1   g0971(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n267), .B1(new_n769), .B2(new_n1120), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1131), .B(new_n1173), .C1(G50), .C2(new_n757), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n764), .A2(G128), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n772), .A2(new_n1095), .B1(new_n778), .B2(new_n795), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(G137), .B2(new_n797), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1174), .A2(new_n1175), .A3(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G150), .B2(new_n761), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n746), .B1(new_n1172), .B2(new_n1179), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1180), .B(new_n737), .C1(G68), .C2(new_n831), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n1068), .B2(new_n740), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1182), .B1(new_n1084), .B2(new_n959), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n934), .B(KEYINPUT117), .Z(new_n1184));
  NAND2_X1  g0984(.A1(new_n1087), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1183), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT119), .Z(G381));
  XNOR2_X1  g0988(.A(G375), .B(KEYINPUT120), .ZN(new_n1189));
  INV_X1    g0989(.A(G378), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1191), .A2(G384), .A3(G381), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n960), .A2(new_n1052), .A3(new_n986), .ZN(new_n1193));
  NOR3_X1   g0993(.A1(new_n1193), .A2(G396), .A3(G393), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1192), .A2(new_n1194), .ZN(G407));
  OAI211_X1 g0995(.A(G407), .B(G213), .C1(G343), .C2(new_n1191), .ZN(G409));
  OAI211_X1 g0996(.A(G378), .B(new_n1160), .C1(new_n1163), .C2(new_n1164), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1161), .A2(new_n1159), .A3(new_n1184), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1160), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1190), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n667), .A2(G213), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1186), .A2(KEYINPUT60), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT60), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1205));
  NAND4_X1  g1005(.A1(new_n1203), .A2(new_n685), .A3(new_n1087), .A4(new_n1205), .ZN(new_n1206));
  AND3_X1   g1006(.A1(G384), .A2(new_n1183), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(G384), .B1(new_n1183), .B2(new_n1206), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1201), .A2(new_n1202), .A3(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT121), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1210), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT62), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1201), .A2(KEYINPUT121), .A3(new_n1202), .A4(new_n1209), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT122), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1212), .A2(KEYINPUT122), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1218));
  NAND4_X1  g1018(.A1(new_n1201), .A2(KEYINPUT62), .A3(new_n1209), .A4(new_n1202), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT123), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1217), .A2(new_n1218), .A3(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n667), .A2(G213), .A3(G2897), .ZN(new_n1222));
  XOR2_X1   g1022(.A(new_n1209), .B(new_n1222), .Z(new_n1223));
  NAND2_X1  g1023(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1224));
  AOI21_X1  g1024(.A(KEYINPUT61), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1221), .A2(new_n1225), .ZN(new_n1226));
  XNOR2_X1  g1026(.A(G393), .B(G396), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(new_n1193), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1052), .B1(new_n960), .B2(new_n986), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1228), .B1(new_n1229), .B2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1230), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1232), .A2(new_n1193), .A3(new_n1227), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1226), .A2(new_n1234), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT63), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1210), .A2(new_n1237), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1234), .A2(new_n1238), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1212), .A2(new_n1237), .A3(new_n1214), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1225), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1235), .A2(new_n1236), .A3(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1234), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(new_n1221), .B2(new_n1225), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1239), .A2(new_n1225), .A3(new_n1240), .ZN(new_n1245));
  OAI21_X1  g1045(.A(KEYINPUT124), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1246), .ZN(G405));
  INV_X1    g1047(.A(new_n1209), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n1197), .B1(new_n1248), .B2(KEYINPUT125), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1249), .B1(G375), .B2(new_n1190), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1234), .B(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(KEYINPUT125), .ZN(new_n1252));
  XOR2_X1   g1052(.A(new_n1252), .B(KEYINPUT126), .Z(new_n1253));
  XNOR2_X1  g1053(.A(new_n1251), .B(new_n1253), .ZN(G402));
endmodule


