

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593;

  XNOR2_X1 U325 ( .A(n464), .B(n463), .ZN(n469) );
  XNOR2_X1 U326 ( .A(n472), .B(n471), .ZN(n531) );
  XNOR2_X1 U327 ( .A(n470), .B(KEYINPUT48), .ZN(n471) );
  XNOR2_X1 U328 ( .A(n314), .B(n313), .ZN(n315) );
  XNOR2_X1 U329 ( .A(n367), .B(KEYINPUT25), .ZN(n368) );
  XNOR2_X1 U330 ( .A(n462), .B(KEYINPUT47), .ZN(n463) );
  XNOR2_X1 U331 ( .A(n369), .B(n368), .ZN(n374) );
  INV_X1 U332 ( .A(G204GAT), .ZN(n414) );
  INV_X1 U333 ( .A(KEYINPUT106), .ZN(n470) );
  INV_X1 U334 ( .A(KEYINPUT21), .ZN(n313) );
  XNOR2_X1 U335 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U336 ( .A(n381), .B(n336), .ZN(n337) );
  XNOR2_X1 U337 ( .A(n417), .B(n416), .ZN(n421) );
  XNOR2_X1 U338 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U339 ( .A(n316), .B(n315), .ZN(n333) );
  XNOR2_X1 U340 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U341 ( .A(n429), .B(n428), .ZN(n449) );
  INV_X1 U342 ( .A(G106GAT), .ZN(n446) );
  XNOR2_X1 U343 ( .A(n482), .B(G190GAT), .ZN(n483) );
  XNOR2_X1 U344 ( .A(n446), .B(KEYINPUT44), .ZN(n447) );
  XNOR2_X1 U345 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U346 ( .A(n484), .B(n483), .ZN(G1351GAT) );
  XNOR2_X1 U347 ( .A(n455), .B(n454), .ZN(G1330GAT) );
  INV_X1 U348 ( .A(KEYINPUT86), .ZN(n344) );
  XOR2_X1 U349 ( .A(G120GAT), .B(G57GAT), .Z(n424) );
  XNOR2_X1 U350 ( .A(G134GAT), .B(G127GAT), .ZN(n293) );
  XNOR2_X1 U351 ( .A(n293), .B(KEYINPUT0), .ZN(n353) );
  XOR2_X1 U352 ( .A(n424), .B(n353), .Z(n295) );
  NAND2_X1 U353 ( .A1(G225GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U354 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U355 ( .A(n296), .B(KEYINPUT5), .Z(n299) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G1GAT), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n297), .B(G141GAT), .ZN(n430) );
  XNOR2_X1 U358 ( .A(n430), .B(KEYINPUT83), .ZN(n298) );
  XNOR2_X1 U359 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U360 ( .A(KEYINPUT81), .B(G85GAT), .Z(n301) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(G148GAT), .ZN(n300) );
  XNOR2_X1 U362 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U363 ( .A(n303), .B(n302), .Z(n311) );
  XOR2_X1 U364 ( .A(G155GAT), .B(G162GAT), .Z(n305) );
  XNOR2_X1 U365 ( .A(KEYINPUT3), .B(KEYINPUT2), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U367 ( .A(KEYINPUT80), .B(n306), .Z(n319) );
  XOR2_X1 U368 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n308) );
  XNOR2_X1 U369 ( .A(KEYINPUT6), .B(KEYINPUT82), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U371 ( .A(n319), .B(n309), .ZN(n310) );
  XNOR2_X1 U372 ( .A(n311), .B(n310), .ZN(n375) );
  XOR2_X2 U373 ( .A(KEYINPUT84), .B(n375), .Z(n522) );
  INV_X1 U374 ( .A(n522), .ZN(n530) );
  XNOR2_X1 U375 ( .A(KEYINPUT79), .B(G211GAT), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n312), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U377 ( .A(G197GAT), .B(KEYINPUT78), .ZN(n314) );
  XOR2_X1 U378 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n321) );
  XOR2_X1 U379 ( .A(G148GAT), .B(KEYINPUT71), .Z(n318) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(G78GAT), .ZN(n317) );
  XNOR2_X1 U381 ( .A(n318), .B(n317), .ZN(n423) );
  XNOR2_X1 U382 ( .A(n319), .B(n423), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U384 ( .A(n333), .B(n322), .ZN(n330) );
  NAND2_X1 U385 ( .A1(G228GAT), .A2(G233GAT), .ZN(n328) );
  XOR2_X1 U386 ( .A(KEYINPUT77), .B(KEYINPUT23), .Z(n324) );
  XNOR2_X1 U387 ( .A(G22GAT), .B(G141GAT), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n326) );
  XOR2_X1 U389 ( .A(G50GAT), .B(G218GAT), .Z(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U392 ( .A(n330), .B(n329), .ZN(n477) );
  XOR2_X1 U393 ( .A(KEYINPUT28), .B(n477), .Z(n528) );
  AND2_X1 U394 ( .A1(n530), .A2(n528), .ZN(n342) );
  XOR2_X1 U395 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n332) );
  XNOR2_X1 U396 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n331) );
  XNOR2_X1 U397 ( .A(n332), .B(n331), .ZN(n354) );
  XNOR2_X1 U398 ( .A(KEYINPUT85), .B(n333), .ZN(n335) );
  XOR2_X1 U399 ( .A(G8GAT), .B(G169GAT), .Z(n437) );
  XOR2_X1 U400 ( .A(G36GAT), .B(n437), .Z(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n338) );
  XOR2_X1 U402 ( .A(G218GAT), .B(G190GAT), .Z(n381) );
  AND2_X1 U403 ( .A1(G226GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n354), .B(n339), .ZN(n341) );
  XOR2_X1 U405 ( .A(G176GAT), .B(G92GAT), .Z(n340) );
  XOR2_X1 U406 ( .A(G64GAT), .B(n340), .Z(n422) );
  XOR2_X1 U407 ( .A(n341), .B(n422), .Z(n496) );
  INV_X1 U408 ( .A(n496), .ZN(n473) );
  XNOR2_X1 U409 ( .A(KEYINPUT27), .B(n473), .ZN(n529) );
  NAND2_X1 U410 ( .A1(n342), .A2(n529), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n363) );
  XOR2_X1 U412 ( .A(KEYINPUT74), .B(G120GAT), .Z(n346) );
  XNOR2_X1 U413 ( .A(G113GAT), .B(G169GAT), .ZN(n345) );
  XNOR2_X1 U414 ( .A(n346), .B(n345), .ZN(n362) );
  XOR2_X1 U415 ( .A(G176GAT), .B(G71GAT), .Z(n348) );
  XNOR2_X1 U416 ( .A(G15GAT), .B(G99GAT), .ZN(n347) );
  XNOR2_X1 U417 ( .A(n348), .B(n347), .ZN(n350) );
  XOR2_X1 U418 ( .A(G43GAT), .B(G190GAT), .Z(n349) );
  XNOR2_X1 U419 ( .A(n350), .B(n349), .ZN(n358) );
  XNOR2_X1 U420 ( .A(KEYINPUT64), .B(KEYINPUT76), .ZN(n351) );
  XNOR2_X1 U421 ( .A(n351), .B(KEYINPUT75), .ZN(n352) );
  XOR2_X1 U422 ( .A(n352), .B(KEYINPUT20), .Z(n356) );
  XNOR2_X1 U423 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U424 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n358), .B(n357), .ZN(n360) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U427 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n362), .B(n361), .ZN(n533) );
  NAND2_X1 U429 ( .A1(n363), .A2(n533), .ZN(n364) );
  XNOR2_X1 U430 ( .A(n364), .B(KEYINPUT87), .ZN(n378) );
  OR2_X1 U431 ( .A1(n533), .A2(n496), .ZN(n365) );
  XNOR2_X1 U432 ( .A(KEYINPUT89), .B(n365), .ZN(n366) );
  NOR2_X1 U433 ( .A1(n477), .A2(n366), .ZN(n369) );
  INV_X1 U434 ( .A(KEYINPUT90), .ZN(n367) );
  XOR2_X1 U435 ( .A(KEYINPUT27), .B(n473), .Z(n372) );
  NAND2_X1 U436 ( .A1(n533), .A2(n477), .ZN(n370) );
  XNOR2_X1 U437 ( .A(n370), .B(KEYINPUT26), .ZN(n371) );
  XNOR2_X1 U438 ( .A(KEYINPUT88), .B(n371), .ZN(n576) );
  NOR2_X1 U439 ( .A1(n372), .A2(n576), .ZN(n373) );
  NOR2_X1 U440 ( .A1(n374), .A2(n373), .ZN(n376) );
  NOR2_X1 U441 ( .A1(n376), .A2(n375), .ZN(n377) );
  NOR2_X1 U442 ( .A1(n378), .A2(n377), .ZN(n491) );
  XOR2_X1 U443 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n380) );
  XNOR2_X1 U444 ( .A(KEYINPUT9), .B(KEYINPUT72), .ZN(n379) );
  XNOR2_X1 U445 ( .A(n380), .B(n379), .ZN(n395) );
  XOR2_X1 U446 ( .A(n381), .B(G92GAT), .Z(n383) );
  NAND2_X1 U447 ( .A1(G232GAT), .A2(G233GAT), .ZN(n382) );
  XNOR2_X1 U448 ( .A(n383), .B(n382), .ZN(n387) );
  XOR2_X1 U449 ( .A(KEYINPUT65), .B(G134GAT), .Z(n385) );
  XNOR2_X1 U450 ( .A(G162GAT), .B(G106GAT), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U452 ( .A(n387), .B(n386), .Z(n393) );
  XNOR2_X1 U453 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n388) );
  XNOR2_X1 U454 ( .A(n388), .B(G29GAT), .ZN(n389) );
  XOR2_X1 U455 ( .A(n389), .B(KEYINPUT8), .Z(n391) );
  XNOR2_X1 U456 ( .A(G43GAT), .B(G50GAT), .ZN(n390) );
  XNOR2_X1 U457 ( .A(n391), .B(n390), .ZN(n442) );
  XOR2_X1 U458 ( .A(G99GAT), .B(G85GAT), .Z(n425) );
  XNOR2_X1 U459 ( .A(n442), .B(n425), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U461 ( .A(n395), .B(n394), .ZN(n561) );
  XOR2_X1 U462 ( .A(KEYINPUT36), .B(n561), .Z(n590) );
  NOR2_X1 U463 ( .A1(n491), .A2(n590), .ZN(n412) );
  XOR2_X1 U464 ( .A(G64GAT), .B(G57GAT), .Z(n397) );
  XNOR2_X1 U465 ( .A(G211GAT), .B(G78GAT), .ZN(n396) );
  XNOR2_X1 U466 ( .A(n397), .B(n396), .ZN(n411) );
  XNOR2_X1 U467 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n398) );
  XNOR2_X1 U468 ( .A(n398), .B(KEYINPUT69), .ZN(n417) );
  XOR2_X1 U469 ( .A(n417), .B(G183GAT), .Z(n400) );
  XOR2_X1 U470 ( .A(G22GAT), .B(G15GAT), .Z(n438) );
  XNOR2_X1 U471 ( .A(n438), .B(G8GAT), .ZN(n399) );
  XNOR2_X1 U472 ( .A(n400), .B(n399), .ZN(n404) );
  XOR2_X1 U473 ( .A(KEYINPUT12), .B(KEYINPUT73), .Z(n402) );
  NAND2_X1 U474 ( .A1(G231GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U475 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U476 ( .A(n404), .B(n403), .Z(n409) );
  XOR2_X1 U477 ( .A(KEYINPUT14), .B(G127GAT), .Z(n406) );
  XNOR2_X1 U478 ( .A(G1GAT), .B(G155GAT), .ZN(n405) );
  XNOR2_X1 U479 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U480 ( .A(n407), .B(KEYINPUT15), .ZN(n408) );
  XNOR2_X1 U481 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U482 ( .A(n411), .B(n410), .ZN(n488) );
  NAND2_X1 U483 ( .A1(n412), .A2(n488), .ZN(n413) );
  XOR2_X1 U484 ( .A(KEYINPUT37), .B(n413), .Z(n450) );
  NAND2_X1 U485 ( .A1(G230GAT), .A2(G233GAT), .ZN(n415) );
  XOR2_X1 U486 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n419) );
  XNOR2_X1 U487 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n418) );
  XNOR2_X1 U488 ( .A(n419), .B(n418), .ZN(n420) );
  XOR2_X1 U489 ( .A(n421), .B(n420), .Z(n429) );
  XNOR2_X1 U490 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U491 ( .A(n425), .B(n424), .Z(n426) );
  XOR2_X1 U492 ( .A(n449), .B(KEYINPUT41), .Z(n539) );
  XOR2_X1 U493 ( .A(n430), .B(KEYINPUT67), .Z(n432) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n431) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n436) );
  XOR2_X1 U496 ( .A(G197GAT), .B(KEYINPUT29), .Z(n434) );
  XNOR2_X1 U497 ( .A(KEYINPUT66), .B(KEYINPUT30), .ZN(n433) );
  XNOR2_X1 U498 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U499 ( .A(n436), .B(n435), .Z(n440) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U502 ( .A(n442), .B(n441), .Z(n456) );
  INV_X1 U503 ( .A(n456), .ZN(n578) );
  NOR2_X1 U504 ( .A1(n539), .A2(n578), .ZN(n443) );
  XOR2_X1 U505 ( .A(n443), .B(KEYINPUT99), .Z(n512) );
  INV_X1 U506 ( .A(n512), .ZN(n444) );
  NOR2_X1 U507 ( .A1(n450), .A2(n444), .ZN(n445) );
  XOR2_X1 U508 ( .A(KEYINPUT102), .B(n445), .Z(n526) );
  NOR2_X1 U509 ( .A1(n526), .A2(n528), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(G1339GAT) );
  XOR2_X1 U511 ( .A(KEYINPUT68), .B(n456), .Z(n565) );
  NAND2_X1 U512 ( .A1(n565), .A2(n449), .ZN(n487) );
  NOR2_X1 U513 ( .A1(n450), .A2(n487), .ZN(n451) );
  XOR2_X1 U514 ( .A(KEYINPUT38), .B(n451), .Z(n509) );
  NOR2_X1 U515 ( .A1(n509), .A2(n533), .ZN(n455) );
  XNOR2_X1 U516 ( .A(KEYINPUT40), .B(KEYINPUT98), .ZN(n453) );
  INV_X1 U517 ( .A(G43GAT), .ZN(n452) );
  INV_X1 U518 ( .A(n488), .ZN(n585) );
  OR2_X1 U519 ( .A1(n539), .A2(n456), .ZN(n458) );
  INV_X1 U520 ( .A(KEYINPUT46), .ZN(n457) );
  XNOR2_X1 U521 ( .A(n458), .B(n457), .ZN(n459) );
  NOR2_X1 U522 ( .A1(n585), .A2(n459), .ZN(n461) );
  INV_X1 U523 ( .A(n561), .ZN(n460) );
  NAND2_X1 U524 ( .A1(n461), .A2(n460), .ZN(n464) );
  XOR2_X1 U525 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n462) );
  NOR2_X1 U526 ( .A1(n590), .A2(n488), .ZN(n465) );
  XNOR2_X1 U527 ( .A(n465), .B(KEYINPUT45), .ZN(n466) );
  NAND2_X1 U528 ( .A1(n466), .A2(n449), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n467), .A2(n565), .ZN(n468) );
  NOR2_X1 U530 ( .A1(n469), .A2(n468), .ZN(n472) );
  NAND2_X1 U531 ( .A1(n473), .A2(n531), .ZN(n475) );
  XOR2_X1 U532 ( .A(KEYINPUT54), .B(KEYINPUT118), .Z(n474) );
  XNOR2_X1 U533 ( .A(n475), .B(n474), .ZN(n476) );
  NAND2_X1 U534 ( .A1(n476), .A2(n522), .ZN(n577) );
  NOR2_X1 U535 ( .A1(n477), .A2(n577), .ZN(n478) );
  XNOR2_X1 U536 ( .A(n478), .B(KEYINPUT55), .ZN(n480) );
  INV_X1 U537 ( .A(KEYINPUT119), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(n481) );
  NOR2_X1 U539 ( .A1(n533), .A2(n481), .ZN(n571) );
  NAND2_X1 U540 ( .A1(n571), .A2(n561), .ZN(n484) );
  XOR2_X1 U541 ( .A(KEYINPUT121), .B(KEYINPUT58), .Z(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT34), .B(KEYINPUT92), .Z(n486) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT93), .ZN(n485) );
  XNOR2_X1 U544 ( .A(n486), .B(n485), .ZN(n495) );
  INV_X1 U545 ( .A(n487), .ZN(n493) );
  NOR2_X1 U546 ( .A1(n561), .A2(n488), .ZN(n489) );
  XOR2_X1 U547 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  NOR2_X1 U548 ( .A1(n491), .A2(n490), .ZN(n492) );
  XOR2_X1 U549 ( .A(KEYINPUT91), .B(n492), .Z(n511) );
  NAND2_X1 U550 ( .A1(n493), .A2(n511), .ZN(n501) );
  NOR2_X1 U551 ( .A1(n522), .A2(n501), .ZN(n494) );
  XOR2_X1 U552 ( .A(n495), .B(n494), .Z(G1324GAT) );
  NOR2_X1 U553 ( .A1(n496), .A2(n501), .ZN(n497) );
  XOR2_X1 U554 ( .A(KEYINPUT94), .B(n497), .Z(n498) );
  XNOR2_X1 U555 ( .A(G8GAT), .B(n498), .ZN(G1325GAT) );
  NOR2_X1 U556 ( .A1(n533), .A2(n501), .ZN(n500) );
  XNOR2_X1 U557 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n499) );
  XNOR2_X1 U558 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U559 ( .A1(n528), .A2(n501), .ZN(n503) );
  XNOR2_X1 U560 ( .A(G22GAT), .B(KEYINPUT95), .ZN(n502) );
  XNOR2_X1 U561 ( .A(n503), .B(n502), .ZN(G1327GAT) );
  XNOR2_X1 U562 ( .A(KEYINPUT96), .B(KEYINPUT39), .ZN(n505) );
  NOR2_X1 U563 ( .A1(n522), .A2(n509), .ZN(n504) );
  XNOR2_X1 U564 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(n506), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n509), .A2(n496), .ZN(n508) );
  XNOR2_X1 U567 ( .A(G36GAT), .B(KEYINPUT97), .ZN(n507) );
  XNOR2_X1 U568 ( .A(n508), .B(n507), .ZN(G1329GAT) );
  NOR2_X1 U569 ( .A1(n509), .A2(n528), .ZN(n510) );
  XOR2_X1 U570 ( .A(G50GAT), .B(n510), .Z(G1331GAT) );
  NAND2_X1 U571 ( .A1(n512), .A2(n511), .ZN(n518) );
  NOR2_X1 U572 ( .A1(n522), .A2(n518), .ZN(n514) );
  XNOR2_X1 U573 ( .A(KEYINPUT100), .B(KEYINPUT42), .ZN(n513) );
  XNOR2_X1 U574 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U575 ( .A(G57GAT), .B(n515), .Z(G1332GAT) );
  NOR2_X1 U576 ( .A1(n496), .A2(n518), .ZN(n516) );
  XOR2_X1 U577 ( .A(G64GAT), .B(n516), .Z(G1333GAT) );
  NOR2_X1 U578 ( .A1(n533), .A2(n518), .ZN(n517) );
  XOR2_X1 U579 ( .A(G71GAT), .B(n517), .Z(G1334GAT) );
  NOR2_X1 U580 ( .A1(n528), .A2(n518), .ZN(n520) );
  XNOR2_X1 U581 ( .A(KEYINPUT43), .B(KEYINPUT101), .ZN(n519) );
  XNOR2_X1 U582 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U583 ( .A(G78GAT), .B(n521), .Z(G1335GAT) );
  NOR2_X1 U584 ( .A1(n522), .A2(n526), .ZN(n523) );
  XOR2_X1 U585 ( .A(G85GAT), .B(n523), .Z(G1336GAT) );
  NOR2_X1 U586 ( .A1(n526), .A2(n496), .ZN(n525) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(KEYINPUT103), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n525), .B(n524), .ZN(G1337GAT) );
  NOR2_X1 U589 ( .A1(n526), .A2(n533), .ZN(n527) );
  XOR2_X1 U590 ( .A(G99GAT), .B(n527), .Z(G1338GAT) );
  INV_X1 U591 ( .A(n528), .ZN(n536) );
  AND2_X1 U592 ( .A1(n530), .A2(n529), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n532), .A2(n531), .ZN(n552) );
  NOR2_X1 U594 ( .A1(n533), .A2(n552), .ZN(n534) );
  XNOR2_X1 U595 ( .A(n534), .B(KEYINPUT107), .ZN(n535) );
  NOR2_X1 U596 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U597 ( .A(KEYINPUT108), .B(n537), .ZN(n549) );
  NAND2_X1 U598 ( .A1(n565), .A2(n549), .ZN(n538) );
  XNOR2_X1 U599 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT109), .Z(n541) );
  INV_X1 U601 ( .A(n539), .ZN(n567) );
  NAND2_X1 U602 ( .A1(n567), .A2(n549), .ZN(n540) );
  XNOR2_X1 U603 ( .A(n541), .B(n540), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT110), .B(KEYINPUT49), .Z(n542) );
  XNOR2_X1 U605 ( .A(n543), .B(n542), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT111), .Z(n545) );
  NAND2_X1 U607 ( .A1(n585), .A2(n549), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT112), .B(KEYINPUT51), .Z(n548) );
  XNOR2_X1 U611 ( .A(G134GAT), .B(KEYINPUT113), .ZN(n547) );
  XNOR2_X1 U612 ( .A(n548), .B(n547), .ZN(n551) );
  NAND2_X1 U613 ( .A1(n549), .A2(n561), .ZN(n550) );
  XOR2_X1 U614 ( .A(n551), .B(n550), .Z(G1343GAT) );
  XOR2_X1 U615 ( .A(G141GAT), .B(KEYINPUT115), .Z(n555) );
  NOR2_X1 U616 ( .A1(n576), .A2(n552), .ZN(n553) );
  XNOR2_X1 U617 ( .A(n553), .B(KEYINPUT114), .ZN(n562) );
  NAND2_X1 U618 ( .A1(n562), .A2(n578), .ZN(n554) );
  XNOR2_X1 U619 ( .A(n555), .B(n554), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n557) );
  NAND2_X1 U621 ( .A1(n567), .A2(n562), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NAND2_X1 U624 ( .A1(n562), .A2(n585), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(KEYINPUT116), .ZN(n560) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  XOR2_X1 U627 ( .A(G162GAT), .B(KEYINPUT117), .Z(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  NAND2_X1 U630 ( .A1(n571), .A2(n565), .ZN(n566) );
  XNOR2_X1 U631 ( .A(n566), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U632 ( .A1(n571), .A2(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U635 ( .A(n570), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n585), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n572), .B(KEYINPUT120), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G183GAT), .B(n573), .ZN(G1350GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT60), .Z(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n582) );
  XOR2_X1 U642 ( .A(G197GAT), .B(KEYINPUT59), .Z(n580) );
  NOR2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n586), .A2(n578), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U647 ( .A(G204GAT), .B(KEYINPUT61), .Z(n584) );
  INV_X1 U648 ( .A(n586), .ZN(n589) );
  OR2_X1 U649 ( .A1(n589), .A2(n449), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  XOR2_X1 U651 ( .A(G211GAT), .B(KEYINPUT125), .Z(n588) );
  NAND2_X1 U652 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1354GAT) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n592) );
  XNOR2_X1 U655 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n591) );
  XNOR2_X1 U656 ( .A(n592), .B(n591), .ZN(n593) );
  XOR2_X1 U657 ( .A(G218GAT), .B(n593), .Z(G1355GAT) );
endmodule

