//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  AND2_X1   g001(.A1(G211gat), .A2(G218gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(G211gat), .A2(G218gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  AND2_X1   g004(.A1(G197gat), .A2(G204gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(G197gat), .A2(G204gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g007(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n205), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(G197gat), .B(G204gat), .ZN(new_n212));
  INV_X1    g011(.A(new_n209), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NOR3_X1   g019(.A1(new_n219), .A2(G169gat), .A3(G176gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(G169gat), .A2(G176gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n221), .A2(KEYINPUT64), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225));
  INV_X1    g024(.A(G169gat), .ZN(new_n226));
  INV_X1    g025(.A(G176gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n226), .A2(new_n227), .A3(KEYINPUT23), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n225), .B1(new_n228), .B2(new_n222), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n220), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G183gat), .ZN(new_n231));
  INV_X1    g030(.A(G190gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n235));
  OAI211_X1 g034(.A(new_n233), .B(new_n234), .C1(new_n235), .C2(KEYINPUT65), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n236), .B1(KEYINPUT65), .B2(new_n235), .ZN(new_n237));
  OAI21_X1  g036(.A(KEYINPUT25), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n231), .A2(KEYINPUT27), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT27), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(G183gat), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n239), .A2(new_n241), .A3(new_n232), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT66), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(KEYINPUT28), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT28), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n245), .A2(KEYINPUT66), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n222), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n218), .A2(new_n249), .ZN(new_n250));
  NOR3_X1   g049(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI22_X1  g051(.A1(new_n242), .A2(new_n247), .B1(new_n250), .B2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n239), .A2(new_n241), .A3(new_n232), .ZN(new_n254));
  INV_X1    g053(.A(new_n244), .ZN(new_n255));
  AOI22_X1  g054(.A1(new_n254), .A2(new_n255), .B1(G183gat), .B2(G190gat), .ZN(new_n256));
  INV_X1    g055(.A(new_n235), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n257), .A2(new_n233), .A3(new_n234), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT25), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n259), .B1(new_n217), .B2(KEYINPUT23), .ZN(new_n260));
  NOR3_X1   g059(.A1(new_n260), .A2(new_n223), .A3(new_n221), .ZN(new_n261));
  AOI22_X1  g060(.A1(new_n253), .A2(new_n256), .B1(new_n258), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(KEYINPUT29), .B1(new_n238), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G226gat), .A2(G233gat), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n216), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n264), .B1(new_n238), .B2(new_n262), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n238), .A2(new_n262), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n267), .B1(new_n270), .B2(new_n264), .ZN(new_n271));
  OAI211_X1 g070(.A(new_n215), .B(new_n266), .C1(new_n271), .C2(new_n216), .ZN(new_n272));
  INV_X1    g071(.A(new_n267), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n273), .B1(new_n265), .B2(new_n263), .ZN(new_n274));
  INV_X1    g073(.A(new_n215), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G8gat), .B(G36gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(G64gat), .B(G92gat), .ZN(new_n278));
  XOR2_X1   g077(.A(new_n277), .B(new_n278), .Z(new_n279));
  NAND4_X1  g078(.A1(new_n272), .A2(new_n276), .A3(KEYINPUT30), .A4(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n280), .B(KEYINPUT75), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT30), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n272), .A2(new_n276), .ZN(new_n283));
  INV_X1    g082(.A(new_n279), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(new_n284), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT80), .ZN(new_n289));
  OR2_X1    g088(.A1(G141gat), .A2(G148gat), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT2), .ZN(new_n291));
  NAND2_X1  g090(.A1(G141gat), .A2(G148gat), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G162gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G155gat), .ZN(new_n295));
  INV_X1    g094(.A(G155gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G162gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n293), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT76), .B(G155gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n291), .B1(new_n300), .B2(G162gat), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n290), .A2(new_n295), .A3(new_n297), .A4(new_n292), .ZN(new_n302));
  OAI211_X1 g101(.A(KEYINPUT77), .B(new_n299), .C1(new_n301), .C2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n306));
  OAI21_X1  g105(.A(G162gat), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT2), .ZN(new_n308));
  AND4_X1   g107(.A1(new_n290), .A2(new_n295), .A3(new_n297), .A4(new_n292), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT77), .B1(new_n310), .B2(new_n299), .ZN(new_n311));
  OAI21_X1  g110(.A(KEYINPUT3), .B1(new_n304), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT3), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n313), .A3(new_n299), .ZN(new_n314));
  XNOR2_X1  g113(.A(G127gat), .B(G134gat), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n316));
  INV_X1    g115(.A(G113gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n317), .A2(G120gat), .ZN(new_n318));
  INV_X1    g117(.A(G120gat), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n319), .A2(G113gat), .ZN(new_n320));
  OAI211_X1 g119(.A(new_n315), .B(new_n316), .C1(new_n318), .C2(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n316), .B1(new_n318), .B2(new_n320), .ZN(new_n322));
  INV_X1    g121(.A(G127gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT67), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT67), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(G127gat), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n324), .A2(new_n326), .A3(new_n327), .A4(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n322), .A2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT68), .B1(new_n323), .B2(G134gat), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT67), .B(G127gat), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n330), .B1(new_n331), .B2(G134gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n321), .B1(new_n329), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n312), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(G225gat), .A2(G233gat), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n338), .A2(KEYINPUT5), .ZN(new_n339));
  INV_X1    g138(.A(new_n332), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(new_n328), .A3(new_n322), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n308), .A2(new_n309), .B1(new_n293), .B2(new_n298), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT4), .ZN(new_n343));
  NAND4_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .A4(new_n321), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n299), .B1(new_n301), .B2(new_n302), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT4), .B1(new_n333), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT78), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n341), .A2(new_n342), .A3(new_n321), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n348), .B1(new_n349), .B2(KEYINPUT4), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n336), .B(new_n339), .C1(new_n347), .C2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT77), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n313), .B1(new_n353), .B2(new_n303), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n337), .B1(new_n354), .B2(new_n334), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n344), .A2(new_n346), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n333), .A2(new_n345), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n353), .A2(new_n303), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n358), .B1(new_n359), .B2(new_n333), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT5), .B1(new_n360), .B2(new_n337), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n351), .B1(new_n357), .B2(new_n361), .ZN(new_n362));
  XNOR2_X1  g161(.A(G1gat), .B(G29gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT0), .ZN(new_n364));
  XNOR2_X1  g163(.A(G57gat), .B(G85gat), .ZN(new_n365));
  XOR2_X1   g164(.A(new_n364), .B(new_n365), .Z(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  AND4_X1   g166(.A1(new_n289), .A2(new_n362), .A3(KEYINPUT6), .A4(new_n367), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n353), .A2(new_n303), .B1(new_n341), .B2(new_n321), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n338), .B1(new_n369), .B2(new_n358), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n370), .B(KEYINPUT5), .C1(new_n355), .C2(new_n356), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n366), .B1(new_n371), .B2(new_n351), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n289), .B1(new_n372), .B2(KEYINPUT6), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n362), .A2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT6), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n371), .A2(new_n366), .A3(new_n351), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(KEYINPUT35), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G22gat), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT29), .B1(new_n210), .B2(new_n214), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n313), .B1(new_n381), .B2(KEYINPUT81), .ZN(new_n382));
  AND3_X1   g181(.A1(new_n215), .A2(KEYINPUT81), .A3(new_n269), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n345), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n314), .A2(new_n269), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(new_n275), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(G228gat), .A2(G233gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT82), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT82), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n387), .A2(new_n391), .A3(new_n388), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n359), .B1(KEYINPUT3), .B2(new_n381), .ZN(new_n394));
  INV_X1    g193(.A(new_n388), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n386), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n380), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n391), .B1(new_n387), .B2(new_n388), .ZN(new_n398));
  AOI211_X1 g197(.A(KEYINPUT82), .B(new_n395), .C1(new_n384), .C2(new_n386), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n380), .B(new_n396), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  OAI21_X1  g200(.A(G78gat), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(G78gat), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n404), .A2(new_n405), .A3(new_n400), .ZN(new_n406));
  XNOR2_X1  g205(.A(KEYINPUT31), .B(G50gat), .ZN(new_n407));
  XNOR2_X1  g206(.A(new_n407), .B(KEYINPUT83), .ZN(new_n408));
  XNOR2_X1  g207(.A(new_n408), .B(G106gat), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n402), .A2(new_n406), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n409), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n404), .A2(new_n405), .A3(new_n400), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n405), .B1(new_n404), .B2(new_n400), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  AND4_X1   g213(.A1(new_n288), .A2(new_n379), .A3(new_n410), .A4(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT71), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT64), .B1(new_n221), .B2(new_n223), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n228), .A2(new_n225), .A3(new_n222), .ZN(new_n418));
  AOI22_X1  g217(.A1(new_n417), .A2(new_n418), .B1(new_n219), .B2(new_n218), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n235), .A2(KEYINPUT65), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n421), .A3(new_n233), .A4(new_n234), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n259), .B1(new_n419), .B2(new_n422), .ZN(new_n423));
  NOR2_X1   g222(.A1(new_n221), .A2(new_n223), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n258), .A2(new_n424), .A3(new_n259), .A4(new_n220), .ZN(new_n425));
  OAI22_X1  g224(.A1(new_n242), .A2(new_n244), .B1(new_n231), .B2(new_n232), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n244), .A2(new_n246), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n428), .A2(new_n217), .ZN(new_n429));
  OAI22_X1  g228(.A1(new_n254), .A2(new_n427), .B1(new_n429), .B2(new_n251), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n425), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(KEYINPUT69), .B1(new_n423), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT69), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n238), .A2(new_n262), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n434), .A3(new_n333), .ZN(new_n435));
  INV_X1    g234(.A(G227gat), .ZN(new_n436));
  INV_X1    g235(.A(G233gat), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n268), .A2(KEYINPUT69), .A3(new_n341), .A4(new_n321), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(KEYINPUT70), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT70), .ZN(new_n442));
  NAND4_X1  g241(.A1(new_n435), .A2(new_n439), .A3(new_n442), .A4(new_n438), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT32), .ZN(new_n445));
  XNOR2_X1  g244(.A(G15gat), .B(G43gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(G71gat), .B(G99gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n445), .B1(new_n449), .B2(KEYINPUT33), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n416), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n450), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT71), .B(new_n452), .C1(new_n441), .C2(new_n443), .ZN(new_n453));
  AOI22_X1  g252(.A1(new_n441), .A2(new_n443), .B1(new_n445), .B2(KEYINPUT33), .ZN(new_n454));
  OAI22_X1  g253(.A1(new_n451), .A2(new_n453), .B1(new_n454), .B2(new_n448), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n435), .A2(new_n439), .ZN(new_n456));
  INV_X1    g255(.A(new_n438), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT72), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n458), .A2(new_n459), .A3(KEYINPUT34), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT34), .B1(new_n458), .B2(new_n459), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  OAI221_X1 g263(.A(new_n462), .B1(new_n454), .B2(new_n448), .C1(new_n451), .C2(new_n453), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT73), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT73), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n455), .A2(new_n467), .A3(new_n463), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n202), .B1(new_n415), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT35), .ZN(new_n471));
  AND4_X1   g270(.A1(new_n464), .A2(new_n414), .A3(new_n410), .A4(new_n465), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT75), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n280), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n280), .A2(new_n473), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n286), .B(new_n285), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT79), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n378), .B(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n374), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n471), .B1(new_n472), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n470), .A2(new_n480), .ZN(new_n481));
  AND3_X1   g280(.A1(new_n415), .A2(new_n202), .A3(new_n469), .ZN(new_n482));
  INV_X1    g281(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n478), .A2(new_n374), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(new_n288), .ZN(new_n485));
  INV_X1    g284(.A(new_n410), .ZN(new_n486));
  INV_X1    g285(.A(new_n414), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n487), .A2(new_n486), .ZN(new_n489));
  OAI21_X1  g288(.A(new_n336), .B1(new_n347), .B2(new_n350), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n338), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT39), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n492), .B1(new_n360), .B2(new_n337), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n490), .A2(new_n492), .A3(new_n338), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n494), .A2(new_n366), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT40), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n372), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n476), .B(new_n498), .C1(new_n497), .C2(new_n496), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n284), .B1(new_n283), .B2(KEYINPUT37), .ZN(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n275), .B(new_n266), .C1(new_n271), .C2(new_n216), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT37), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n503), .B1(new_n274), .B2(new_n215), .ZN(new_n504));
  AOI21_X1  g303(.A(KEYINPUT38), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n283), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n501), .A2(new_n505), .B1(new_n506), .B2(new_n279), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n506), .A2(new_n503), .ZN(new_n508));
  OAI21_X1  g307(.A(KEYINPUT38), .B1(new_n508), .B2(new_n500), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n507), .A2(new_n509), .A3(new_n374), .A4(new_n378), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n499), .A3(new_n510), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n488), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT36), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n466), .A2(new_n513), .A3(new_n468), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n464), .A2(new_n465), .A3(KEYINPUT36), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g315(.A1(new_n481), .A2(new_n483), .B1(new_n512), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(G229gat), .A2(G233gat), .ZN(new_n518));
  XOR2_X1   g317(.A(new_n518), .B(KEYINPUT13), .Z(new_n519));
  INV_X1    g318(.A(G50gat), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT15), .B1(new_n520), .B2(G43gat), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n521), .B1(G43gat), .B2(new_n520), .ZN(new_n522));
  XNOR2_X1  g321(.A(KEYINPUT14), .B(G29gat), .ZN(new_n523));
  INV_X1    g322(.A(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(G29gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n522), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT85), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n522), .B1(new_n525), .B2(new_n527), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n520), .A2(G43gat), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n520), .A2(G43gat), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n531), .B1(new_n532), .B2(KEYINPUT87), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n533), .B1(KEYINPUT87), .B2(new_n532), .ZN(new_n534));
  XNOR2_X1  g333(.A(KEYINPUT86), .B(KEYINPUT15), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G15gat), .B(G22gat), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT16), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n537), .B1(new_n538), .B2(G1gat), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n539), .B1(G1gat), .B2(new_n537), .ZN(new_n540));
  XOR2_X1   g339(.A(new_n540), .B(G8gat), .Z(new_n541));
  AND3_X1   g340(.A1(new_n529), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n541), .B1(new_n529), .B2(new_n536), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n519), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  XOR2_X1   g343(.A(new_n544), .B(KEYINPUT89), .Z(new_n545));
  INV_X1    g344(.A(KEYINPUT17), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n536), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n529), .B2(new_n536), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n541), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT88), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n550), .A2(KEYINPUT88), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n553), .A2(KEYINPUT18), .A3(new_n518), .A4(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n549), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(new_n547), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(new_n552), .A3(new_n541), .ZN(new_n558));
  INV_X1    g357(.A(new_n543), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n554), .A2(new_n558), .A3(new_n518), .A4(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT18), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n545), .A2(new_n555), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G113gat), .B(G141gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n564), .B(G197gat), .ZN(new_n565));
  XOR2_X1   g364(.A(KEYINPUT11), .B(G169gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT12), .Z(new_n568));
  NAND2_X1  g367(.A1(new_n563), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  INV_X1    g369(.A(new_n568), .ZN(new_n571));
  NAND4_X1  g370(.A1(new_n545), .A2(new_n555), .A3(new_n562), .A4(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n569), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n563), .A2(KEYINPUT90), .A3(new_n568), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g374(.A(G57gat), .B(G64gat), .Z(new_n576));
  INV_X1    g375(.A(G71gat), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n577), .A2(new_n405), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n576), .B1(KEYINPUT9), .B2(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G71gat), .B(G78gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(KEYINPUT21), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G231gat), .A2(G233gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  XOR2_X1   g384(.A(G127gat), .B(G155gat), .Z(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT20), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n585), .B(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G183gat), .B(G211gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n588), .B(new_n589), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n541), .B1(new_n582), .B2(new_n581), .ZN(new_n591));
  XOR2_X1   g390(.A(KEYINPUT91), .B(KEYINPUT19), .Z(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  OR2_X1    g393(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n590), .A2(new_n594), .ZN(new_n596));
  AND2_X1   g395(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AND2_X1   g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n604), .A2(KEYINPUT93), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n606), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT93), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n599), .A2(new_n603), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(new_n605), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n581), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT10), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n579), .B(new_n580), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n615), .A2(new_n608), .A3(new_n611), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n613), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n612), .A2(new_n607), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n615), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT95), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G230gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n617), .A2(KEYINPUT95), .A3(new_n619), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n613), .A2(new_n616), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n622), .ZN(new_n627));
  XNOR2_X1  g426(.A(G120gat), .B(G148gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(G176gat), .B(G204gat), .ZN(new_n629));
  XOR2_X1   g428(.A(new_n628), .B(new_n629), .Z(new_n630));
  NAND3_X1  g429(.A1(new_n625), .A2(new_n627), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n617), .A2(new_n619), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(new_n621), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n627), .ZN(new_n634));
  INV_X1    g433(.A(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n529), .A2(new_n536), .ZN(new_n639));
  AND2_X1   g438(.A1(G232gat), .A2(G233gat), .ZN(new_n640));
  AOI22_X1  g439(.A1(new_n639), .A2(new_n618), .B1(KEYINPUT41), .B2(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT94), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n557), .A2(new_n607), .A3(new_n612), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n640), .A2(KEYINPUT41), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT92), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n644), .A2(new_n646), .ZN(new_n647));
  OR2_X1    g446(.A1(new_n644), .A2(new_n646), .ZN(new_n648));
  XNOR2_X1  g447(.A(G190gat), .B(G218gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(G134gat), .B(G162gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  AND3_X1   g450(.A1(new_n647), .A2(new_n648), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n648), .B2(new_n647), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n597), .A2(new_n638), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n517), .A2(new_n575), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n484), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(KEYINPUT96), .B(G1gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(G1324gat));
  XOR2_X1   g460(.A(KEYINPUT16), .B(G8gat), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n657), .A2(new_n476), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n657), .ZN(new_n664));
  OAI21_X1  g463(.A(G8gat), .B1(new_n664), .B2(new_n288), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n663), .ZN(new_n666));
  MUX2_X1   g465(.A(new_n663), .B(new_n666), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g466(.A(G15gat), .B1(new_n664), .B2(new_n516), .ZN(new_n668));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n657), .A2(new_n669), .A3(new_n469), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(new_n670), .ZN(G1326gat));
  INV_X1    g470(.A(new_n489), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(KEYINPUT43), .B(G22gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(G1327gat));
  NAND3_X1  g474(.A1(new_n516), .A2(new_n488), .A3(new_n511), .ZN(new_n676));
  NAND4_X1  g475(.A1(new_n414), .A2(new_n464), .A3(new_n410), .A4(new_n465), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT35), .B1(new_n485), .B2(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n288), .A2(new_n379), .A3(new_n414), .A4(new_n410), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n468), .B2(new_n466), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n678), .B1(new_n680), .B2(new_n202), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n676), .B1(new_n681), .B2(new_n482), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n597), .A2(new_n575), .A3(new_n637), .ZN(new_n683));
  AND3_X1   g482(.A1(new_n682), .A2(new_n654), .A3(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n526), .A3(new_n658), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT44), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n687), .B1(new_n517), .B2(new_n655), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(KEYINPUT44), .A3(new_n654), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n688), .A2(new_n689), .A3(new_n683), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND4_X1  g491(.A1(new_n688), .A2(KEYINPUT97), .A3(new_n689), .A4(new_n683), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n692), .A2(new_n658), .A3(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n686), .B1(new_n694), .B2(new_n526), .ZN(G1328gat));
  AOI21_X1  g494(.A(G36gat), .B1(KEYINPUT98), .B2(KEYINPUT46), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n684), .A2(new_n476), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(KEYINPUT98), .A2(KEYINPUT46), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n692), .A2(new_n476), .A3(new_n693), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n699), .B1(new_n700), .B2(new_n524), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT99), .ZN(G1329gat));
  INV_X1    g501(.A(G43gat), .ZN(new_n703));
  AND3_X1   g502(.A1(new_n684), .A2(new_n703), .A3(new_n469), .ZN(new_n704));
  INV_X1    g503(.A(new_n516), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n692), .A2(new_n705), .A3(new_n693), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(G43gat), .ZN(new_n707));
  INV_X1    g506(.A(new_n690), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n703), .B1(new_n708), .B2(new_n705), .ZN(new_n709));
  INV_X1    g508(.A(KEYINPUT47), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n704), .A2(new_n710), .ZN(new_n711));
  OAI22_X1  g510(.A1(new_n707), .A2(KEYINPUT47), .B1(new_n709), .B2(new_n711), .ZN(G1330gat));
  OAI21_X1  g511(.A(G50gat), .B1(new_n690), .B2(new_n489), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n684), .A2(new_n520), .A3(new_n672), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n713), .A2(KEYINPUT48), .A3(new_n715), .ZN(new_n716));
  NAND3_X1  g515(.A1(new_n692), .A2(new_n672), .A3(new_n693), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n714), .B1(new_n717), .B2(G50gat), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n718), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g518(.A(new_n597), .ZN(new_n720));
  INV_X1    g519(.A(new_n575), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n720), .A2(new_n721), .A3(new_n654), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n722), .A2(new_n637), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n682), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n484), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(G57gat), .Z(G1332gat));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n288), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  OAI21_X1  g530(.A(G71gat), .B1(new_n724), .B2(new_n516), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n469), .A2(new_n577), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n732), .B1(new_n724), .B2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(new_n734), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g534(.A1(new_n724), .A2(new_n489), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n736), .B(new_n405), .ZN(G1335gat));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT100), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n482), .A2(new_n470), .A3(new_n480), .ZN(new_n740));
  INV_X1    g539(.A(new_n676), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n739), .B(new_n654), .C1(new_n740), .C2(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n720), .A2(new_n575), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n739), .B1(new_n682), .B2(new_n654), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n738), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT100), .B1(new_n517), .B2(new_n655), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n748), .A2(KEYINPUT51), .A3(new_n744), .A4(new_n742), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n638), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n601), .A3(new_n658), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n743), .A2(new_n638), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n688), .A2(new_n689), .A3(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G85gat), .B1(new_n753), .B2(new_n484), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(G1336gat));
  NAND4_X1  g554(.A1(new_n688), .A2(new_n476), .A3(new_n689), .A4(new_n752), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G92gat), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT101), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n756), .A2(KEYINPUT101), .A3(G92gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n288), .A2(G92gat), .ZN(new_n762));
  INV_X1    g561(.A(new_n762), .ZN(new_n763));
  AOI211_X1 g562(.A(new_n638), .B(new_n763), .C1(new_n747), .C2(new_n749), .ZN(new_n764));
  OAI21_X1  g563(.A(KEYINPUT52), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n762), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT103), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n764), .A2(KEYINPUT103), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT52), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .A4(new_n757), .ZN(new_n773));
  OAI211_X1 g572(.A(KEYINPUT102), .B(KEYINPUT52), .C1(new_n761), .C2(new_n764), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n767), .A2(new_n773), .A3(new_n774), .ZN(G1337gat));
  INV_X1    g574(.A(G99gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n750), .A2(new_n776), .A3(new_n469), .ZN(new_n777));
  OAI21_X1  g576(.A(G99gat), .B1(new_n753), .B2(new_n516), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(G1338gat));
  XOR2_X1   g578(.A(KEYINPUT104), .B(G106gat), .Z(new_n780));
  OAI21_X1  g579(.A(new_n780), .B1(new_n753), .B2(new_n489), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n489), .A2(G106gat), .A3(new_n638), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n783), .B1(new_n747), .B2(new_n749), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT105), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g585(.A(KEYINPUT105), .B(new_n783), .C1(new_n747), .C2(new_n749), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT106), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  OAI211_X1 g589(.A(KEYINPUT106), .B(KEYINPUT53), .C1(new_n786), .C2(new_n787), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT107), .ZN(new_n792));
  OR2_X1    g591(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT53), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n784), .A2(new_n792), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n793), .A2(new_n794), .A3(new_n781), .A4(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n790), .A2(new_n791), .A3(new_n796), .ZN(G1339gat));
  INV_X1    g596(.A(KEYINPUT109), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT54), .B1(new_n632), .B2(new_n621), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n623), .B2(new_n624), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT108), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g601(.A(new_n624), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n803), .A2(new_n620), .A3(new_n622), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT108), .B1(new_n804), .B2(new_n799), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n635), .B1(new_n633), .B2(KEYINPUT54), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n802), .A2(new_n805), .A3(KEYINPUT55), .A4(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n798), .B1(new_n808), .B2(new_n631), .ZN(new_n809));
  INV_X1    g608(.A(new_n799), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n625), .A2(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n806), .B1(new_n811), .B2(KEYINPUT108), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT55), .B1(new_n812), .B2(new_n802), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n808), .A2(new_n798), .A3(new_n631), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n814), .A2(new_n574), .A3(new_n573), .A4(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n518), .B1(new_n553), .B2(new_n554), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n542), .A2(new_n543), .A3(new_n519), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n567), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n572), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n637), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n654), .B1(new_n816), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(new_n815), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n823), .A2(new_n809), .A3(new_n813), .ZN(new_n824));
  AND3_X1   g623(.A1(new_n824), .A2(new_n654), .A3(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n720), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  NOR4_X1   g625(.A1(new_n720), .A2(new_n721), .A3(new_n637), .A4(new_n654), .ZN(new_n827));
  INV_X1    g626(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n469), .A2(new_n489), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR3_X1   g630(.A1(new_n831), .A2(new_n484), .A3(new_n476), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n317), .B1(new_n832), .B2(new_n721), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT110), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n829), .A2(new_n658), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n677), .A2(new_n476), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(new_n838), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n839), .A2(new_n317), .A3(new_n721), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n834), .A2(new_n840), .ZN(G1340gat));
  AOI21_X1  g640(.A(new_n319), .B1(new_n832), .B2(new_n637), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT111), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n839), .A2(new_n319), .A3(new_n637), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(G1341gat));
  AOI21_X1  g644(.A(new_n331), .B1(new_n832), .B2(new_n597), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n597), .A2(new_n331), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n846), .B1(new_n839), .B2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT112), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n848), .B(new_n849), .ZN(G1342gat));
  OR3_X1    g649(.A1(new_n838), .A2(G134gat), .A3(new_n655), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  INV_X1    g651(.A(new_n832), .ZN(new_n853));
  OAI21_X1  g652(.A(G134gat), .B1(new_n853), .B2(new_n655), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n854), .A3(new_n855), .ZN(G1343gat));
  INV_X1    g655(.A(KEYINPUT58), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n484), .A2(new_n476), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n516), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT113), .ZN(new_n860));
  INV_X1    g659(.A(new_n802), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n807), .B1(new_n800), .B2(new_n801), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n812), .A2(KEYINPUT113), .A3(new_n802), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT55), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AND2_X1   g665(.A1(new_n808), .A2(new_n631), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n573), .A3(new_n574), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n821), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n655), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n824), .A2(new_n654), .A3(new_n820), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n597), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n672), .B1(new_n872), .B2(new_n827), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n859), .B1(new_n873), .B2(KEYINPUT57), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n489), .B1(new_n826), .B2(new_n828), .ZN(new_n875));
  INV_X1    g674(.A(KEYINPUT57), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n878), .B2(new_n575), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n857), .B1(new_n879), .B2(KEYINPUT115), .ZN(new_n880));
  OR2_X1    g679(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n835), .A2(KEYINPUT114), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n516), .A2(new_n672), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n883), .A2(new_n476), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n575), .A2(G141gat), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n879), .B1(new_n885), .B2(new_n887), .ZN(new_n888));
  XNOR2_X1  g687(.A(new_n880), .B(new_n888), .ZN(G1344gat));
  INV_X1    g688(.A(new_n885), .ZN(new_n890));
  INV_X1    g689(.A(G148gat), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n890), .A2(new_n891), .A3(new_n637), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT59), .ZN(new_n893));
  NAND4_X1  g692(.A1(new_n814), .A2(KEYINPUT117), .A3(new_n654), .A4(new_n815), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n820), .ZN(new_n895));
  AOI21_X1  g694(.A(KEYINPUT117), .B1(new_n824), .B2(new_n654), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n870), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n827), .B1(new_n897), .B2(new_n720), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n876), .B1(new_n898), .B2(new_n489), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT118), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  AOI211_X1 g700(.A(new_n876), .B(new_n489), .C1(new_n826), .C2(new_n828), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(KEYINPUT118), .B(new_n876), .C1(new_n898), .C2(new_n489), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n638), .B1(new_n859), .B2(KEYINPUT116), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n905), .B(new_n906), .C1(KEYINPUT116), .C2(new_n859), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n893), .B1(new_n907), .B2(G148gat), .ZN(new_n908));
  INV_X1    g707(.A(new_n878), .ZN(new_n909));
  AOI211_X1 g708(.A(KEYINPUT59), .B(new_n891), .C1(new_n909), .C2(new_n637), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n892), .B1(new_n908), .B2(new_n910), .ZN(G1345gat));
  AOI21_X1  g710(.A(new_n300), .B1(new_n890), .B2(new_n597), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n597), .A2(new_n300), .ZN(new_n913));
  XOR2_X1   g712(.A(new_n913), .B(KEYINPUT119), .Z(new_n914));
  AOI21_X1  g713(.A(new_n912), .B1(new_n909), .B2(new_n914), .ZN(G1346gat));
  NOR3_X1   g714(.A1(new_n878), .A2(new_n294), .A3(new_n655), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n890), .A2(new_n654), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n916), .B1(new_n917), .B2(new_n294), .ZN(G1347gat));
  NOR2_X1   g717(.A1(new_n658), .A2(new_n288), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n829), .A2(new_n830), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g719(.A1(new_n920), .A2(new_n226), .A3(new_n575), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n658), .B1(new_n826), .B2(new_n828), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n677), .A2(new_n288), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT120), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n721), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n921), .B1(new_n926), .B2(new_n226), .ZN(G1348gat));
  NAND3_X1  g726(.A1(new_n925), .A2(new_n227), .A3(new_n637), .ZN(new_n928));
  OAI21_X1  g727(.A(G176gat), .B1(new_n920), .B2(new_n638), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n928), .A2(new_n929), .ZN(G1349gat));
  OAI21_X1  g729(.A(G183gat), .B1(new_n920), .B2(new_n720), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT121), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n597), .A2(new_n239), .A3(new_n241), .ZN(new_n933));
  AND3_X1   g732(.A1(new_n925), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n925), .B2(new_n933), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n931), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  OR2_X1    g736(.A1(new_n920), .A2(new_n655), .ZN(new_n938));
  AND2_X1   g737(.A1(new_n938), .A2(G190gat), .ZN(new_n939));
  OR2_X1    g738(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(KEYINPUT61), .A3(new_n941), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n939), .A2(KEYINPUT122), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT61), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n655), .A2(G190gat), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n943), .A2(new_n944), .B1(new_n925), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n942), .A2(new_n946), .ZN(G1351gat));
  INV_X1    g746(.A(G197gat), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n516), .A2(new_n919), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n902), .B1(new_n899), .B2(new_n900), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n949), .B1(new_n950), .B2(new_n904), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n948), .B1(new_n951), .B2(new_n721), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n883), .A2(new_n288), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n922), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n954), .A2(new_n948), .A3(new_n721), .ZN(new_n955));
  XNOR2_X1  g754(.A(new_n955), .B(KEYINPUT123), .ZN(new_n956));
  OAI21_X1  g755(.A(KEYINPUT124), .B1(new_n952), .B2(new_n956), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n955), .B(new_n958), .ZN(new_n959));
  INV_X1    g758(.A(KEYINPUT124), .ZN(new_n960));
  AOI211_X1 g759(.A(new_n575), .B(new_n949), .C1(new_n950), .C2(new_n904), .ZN(new_n961));
  OAI211_X1 g760(.A(new_n959), .B(new_n960), .C1(new_n961), .C2(new_n948), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n957), .A2(new_n962), .ZN(G1352gat));
  INV_X1    g762(.A(KEYINPUT125), .ZN(new_n964));
  INV_X1    g763(.A(new_n949), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n905), .A2(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n964), .B1(new_n966), .B2(new_n638), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n951), .A2(KEYINPUT125), .A3(new_n637), .ZN(new_n968));
  NAND3_X1  g767(.A1(new_n967), .A2(G204gat), .A3(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n954), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n970), .A2(G204gat), .A3(new_n638), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n971), .B(KEYINPUT62), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n969), .A2(new_n972), .ZN(G1353gat));
  OR3_X1    g772(.A1(new_n970), .A2(G211gat), .A3(new_n720), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n905), .A2(new_n597), .A3(new_n965), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n975), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n976));
  AOI21_X1  g775(.A(KEYINPUT63), .B1(new_n975), .B2(G211gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1354gat));
  NAND3_X1  g777(.A1(new_n922), .A2(new_n654), .A3(new_n953), .ZN(new_n979));
  INV_X1    g778(.A(G218gat), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT126), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n981), .B(new_n982), .ZN(new_n983));
  NOR2_X1   g782(.A1(new_n655), .A2(new_n980), .ZN(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n983), .B1(new_n966), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n986), .A2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g786(.A(KEYINPUT127), .ZN(new_n988));
  OAI211_X1 g787(.A(new_n983), .B(new_n988), .C1(new_n966), .C2(new_n985), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n987), .A2(new_n989), .ZN(G1355gat));
endmodule


