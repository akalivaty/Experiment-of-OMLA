//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n608,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n680, new_n681, new_n682, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT78), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G131), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  AOI21_X1  g006(.A(KEYINPUT11), .B1(new_n192), .B2(G134), .ZN(new_n193));
  INV_X1    g007(.A(G134), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G137), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT64), .A2(G137), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT64), .A2(G137), .ZN(new_n197));
  OAI211_X1 g011(.A(KEYINPUT11), .B(G134), .C1(new_n196), .C2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n191), .B1(new_n195), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n195), .A2(new_n198), .A3(new_n191), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G104), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n203), .A2(KEYINPUT3), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT80), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G107), .ZN(new_n206));
  INV_X1    g020(.A(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT80), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n203), .A2(G107), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n203), .B2(G107), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT79), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n207), .A2(G104), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT79), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT3), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n209), .A2(new_n210), .A3(new_n212), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT81), .B1(new_n216), .B2(G101), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT80), .B(G107), .ZN(new_n218));
  OR2_X1    g032(.A1(new_n203), .A2(KEYINPUT3), .ZN(new_n219));
  OAI21_X1  g033(.A(new_n210), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n212), .A2(new_n215), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT81), .ZN(new_n223));
  INV_X1    g037(.A(G101), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n217), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G143), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G146), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G143), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n232), .A2(new_n228), .A3(new_n229), .A4(G128), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT66), .ZN(new_n234));
  XNOR2_X1  g048(.A(G143), .B(G146), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n229), .A4(G128), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n230), .B1(new_n234), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n238), .B1(G128), .B2(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n218), .A2(new_n203), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(new_n213), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G101), .ZN(new_n242));
  AND3_X1   g056(.A1(new_n226), .A2(new_n239), .A3(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n239), .B1(new_n226), .B2(new_n242), .ZN(new_n244));
  OAI211_X1 g058(.A(KEYINPUT12), .B(new_n202), .C1(new_n243), .C2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT82), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n212), .A2(new_n215), .ZN(new_n247));
  NOR2_X1   g061(.A1(new_n220), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n223), .B1(new_n248), .B2(new_n224), .ZN(new_n249));
  NOR3_X1   g063(.A1(new_n216), .A2(KEYINPUT81), .A3(G101), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n242), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n235), .A2(G128), .ZN(new_n252));
  AOI211_X1 g066(.A(new_n230), .B(new_n252), .C1(new_n234), .C2(new_n237), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n226), .A2(new_n239), .A3(new_n242), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT82), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT12), .A4(new_n202), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n202), .B1(new_n243), .B2(new_n244), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT12), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n246), .A2(new_n258), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT84), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n216), .A2(G101), .ZN(new_n265));
  OAI211_X1 g079(.A(KEYINPUT4), .B(new_n265), .C1(new_n249), .C2(new_n250), .ZN(new_n266));
  NAND2_X1  g080(.A1(KEYINPUT0), .A2(G128), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n235), .A2(new_n267), .ZN(new_n268));
  XOR2_X1   g082(.A(KEYINPUT0), .B(G128), .Z(new_n269));
  OAI21_X1  g083(.A(new_n268), .B1(new_n269), .B2(new_n235), .ZN(new_n270));
  OR2_X1    g084(.A1(new_n265), .A2(KEYINPUT4), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT10), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n255), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n226), .A2(KEYINPUT10), .A3(new_n239), .A4(new_n242), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(new_n202), .ZN(new_n277));
  XNOR2_X1  g091(.A(G110), .B(G140), .ZN(new_n278));
  INV_X1    g092(.A(G227), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G953), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n278), .B(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n246), .A2(new_n258), .A3(new_n261), .A4(KEYINPUT84), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n264), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n272), .A2(new_n274), .A3(KEYINPUT83), .A4(new_n275), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n202), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n277), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(new_n281), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n292), .A2(new_n293), .A3(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT85), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(G902), .B1(new_n284), .B2(new_n291), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n298), .A2(KEYINPUT85), .A3(new_n293), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n262), .A2(new_n289), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n281), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n282), .A2(new_n288), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n294), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G469), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n190), .B1(new_n300), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(G214), .B1(G237), .B2(G902), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n270), .A2(G125), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n309), .B1(new_n253), .B2(G125), .ZN(new_n310));
  INV_X1    g124(.A(G224), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G953), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n310), .B(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT6), .ZN(new_n315));
  NAND2_X1  g129(.A1(KEYINPUT2), .A2(G113), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT67), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g132(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(KEYINPUT2), .B2(G113), .ZN(new_n321));
  XNOR2_X1  g135(.A(G116), .B(G119), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n320), .B(new_n322), .C1(KEYINPUT2), .C2(G113), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n266), .A2(new_n326), .A3(new_n271), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT5), .ZN(new_n328));
  INV_X1    g142(.A(G119), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(new_n329), .A3(G116), .ZN(new_n330));
  OAI211_X1 g144(.A(G113), .B(new_n330), .C1(new_n323), .C2(new_n328), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n331), .A2(new_n325), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n226), .A2(KEYINPUT86), .A3(new_n242), .A4(new_n332), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n226), .A2(new_n242), .A3(new_n332), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT86), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n327), .A2(new_n333), .A3(new_n336), .ZN(new_n337));
  XOR2_X1   g151(.A(G110), .B(G122), .Z(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT87), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n338), .ZN(new_n341));
  NAND4_X1  g155(.A1(new_n327), .A2(new_n336), .A3(new_n341), .A4(new_n333), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n315), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT6), .B1(new_n337), .B2(new_n339), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n314), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n314), .B1(KEYINPUT7), .B2(new_n312), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n338), .B(KEYINPUT8), .Z(new_n347));
  INV_X1    g161(.A(new_n334), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n332), .B1(new_n226), .B2(new_n242), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n310), .A2(KEYINPUT7), .A3(new_n312), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n346), .A2(new_n342), .A3(new_n350), .A4(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n345), .A2(new_n294), .A3(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G210), .B1(G237), .B2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT88), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n345), .A2(new_n294), .A3(new_n354), .A4(new_n352), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(KEYINPUT88), .A3(new_n355), .ZN(new_n360));
  AOI21_X1  g174(.A(KEYINPUT13), .B1(new_n227), .B2(G128), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n361), .B(KEYINPUT94), .Z(new_n362));
  OAI21_X1  g176(.A(KEYINPUT95), .B1(new_n227), .B2(G128), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n227), .A2(KEYINPUT13), .A3(G128), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT95), .ZN(new_n366));
  OAI211_X1 g180(.A(new_n362), .B(new_n365), .C1(new_n366), .C2(new_n364), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G134), .ZN(new_n368));
  INV_X1    g182(.A(G122), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G116), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT93), .ZN(new_n371));
  INV_X1    g185(.A(G116), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G122), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g188(.A(new_n374), .B(new_n218), .ZN(new_n375));
  XNOR2_X1  g189(.A(G128), .B(G143), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(new_n194), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(KEYINPUT96), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n368), .A2(new_n375), .A3(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n371), .B1(KEYINPUT14), .B2(new_n373), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n373), .A2(KEYINPUT14), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT97), .ZN(new_n382));
  OAI21_X1  g196(.A(G107), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n376), .B(new_n194), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n383), .B(new_n384), .C1(new_n218), .C2(new_n374), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G217), .ZN(new_n387));
  NOR3_X1   g201(.A1(new_n188), .A2(new_n387), .A3(G953), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n379), .A2(new_n385), .A3(new_n388), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n294), .ZN(new_n393));
  INV_X1    g207(.A(G478), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(KEYINPUT15), .ZN(new_n395));
  XNOR2_X1  g209(.A(new_n393), .B(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G953), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n397), .A2(G952), .ZN(new_n398));
  INV_X1    g212(.A(G234), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  AOI211_X1 g216(.A(new_n294), .B(new_n397), .C1(G234), .C2(G237), .ZN(new_n403));
  XOR2_X1   g217(.A(KEYINPUT21), .B(G898), .Z(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n402), .B1(new_n403), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT90), .ZN(new_n407));
  INV_X1    g221(.A(G140), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G125), .ZN(new_n409));
  INV_X1    g223(.A(G125), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(G140), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(KEYINPUT89), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT89), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n414), .B1(new_n409), .B2(new_n411), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT19), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n412), .A2(KEYINPUT19), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n407), .B1(new_n418), .B2(G146), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n409), .A2(KEYINPUT16), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n409), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G146), .A3(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n400), .A2(new_n397), .A3(G214), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n423), .B(new_n227), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(G131), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n423), .B(G143), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n426), .A2(new_n191), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n416), .A2(KEYINPUT90), .A3(new_n231), .A4(new_n417), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n419), .A2(new_n422), .A3(new_n428), .A4(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n412), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n231), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n413), .A2(new_n415), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n432), .B1(new_n433), .B2(new_n231), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT18), .ZN(new_n435));
  OAI21_X1  g249(.A(new_n426), .B1(new_n435), .B2(new_n191), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n434), .B(new_n436), .C1(new_n435), .C2(new_n425), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n430), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(G113), .B(G122), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n439), .B(new_n203), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT17), .ZN(new_n443));
  OAI21_X1  g257(.A(KEYINPUT91), .B1(new_n425), .B2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n425), .A2(new_n427), .A3(new_n443), .ZN(new_n445));
  INV_X1    g259(.A(new_n422), .ZN(new_n446));
  AOI21_X1  g260(.A(G146), .B1(new_n420), .B2(new_n421), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT91), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n424), .A2(new_n449), .A3(KEYINPUT17), .A4(G131), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n444), .A2(new_n445), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n440), .A3(new_n437), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(G475), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(KEYINPUT20), .A3(new_n454), .A4(new_n294), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n440), .B1(new_n451), .B2(new_n437), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT92), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n452), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n457), .B(new_n294), .C1(new_n459), .C2(new_n456), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G475), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n440), .B1(new_n430), .B2(new_n437), .ZN(new_n462));
  INV_X1    g276(.A(new_n452), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n454), .B(new_n294), .C1(new_n462), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT20), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n455), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n396), .A2(new_n406), .A3(new_n467), .ZN(new_n468));
  AND3_X1   g282(.A1(new_n359), .A2(new_n360), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g283(.A1(new_n307), .A2(new_n308), .A3(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT76), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n472), .B1(new_n329), .B2(G128), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n329), .A2(G128), .ZN(new_n474));
  INV_X1    g288(.A(G128), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT23), .A3(G119), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  XOR2_X1   g291(.A(KEYINPUT24), .B(G110), .Z(new_n478));
  XNOR2_X1  g292(.A(G119), .B(G128), .ZN(new_n479));
  OAI22_X1  g293(.A1(new_n477), .A2(G110), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n422), .A3(new_n432), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT72), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(G110), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n479), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n484), .B(new_n485), .C1(new_n446), .C2(new_n447), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n480), .A2(KEYINPUT72), .A3(new_n422), .A4(new_n432), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT73), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT73), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n483), .A2(new_n486), .A3(new_n490), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n489), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n397), .A2(G221), .A3(G234), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT22), .B(G137), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n495), .B(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n471), .B1(new_n492), .B2(new_n498), .ZN(new_n499));
  AOI211_X1 g313(.A(KEYINPUT76), .B(new_n497), .C1(new_n489), .C2(new_n491), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n488), .A2(new_n498), .ZN(new_n501));
  NOR3_X1   g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n399), .B2(G217), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g318(.A(new_n504), .B(KEYINPUT77), .Z(new_n505));
  INV_X1    g319(.A(new_n499), .ZN(new_n506));
  INV_X1    g320(.A(new_n501), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n492), .A2(new_n471), .A3(new_n498), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n506), .A2(new_n294), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT25), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n502), .A2(KEYINPUT25), .A3(new_n294), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(G217), .B1(new_n399), .B2(G902), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT71), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n513), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n505), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G472), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n194), .A2(G137), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(KEYINPUT65), .ZN(new_n522));
  NOR3_X1   g336(.A1(new_n196), .A2(new_n197), .A3(G134), .ZN(new_n523));
  OAI21_X1  g337(.A(G131), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n201), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n525), .A2(new_n253), .ZN(new_n526));
  INV_X1    g340(.A(new_n201), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n270), .B1(new_n527), .B2(new_n199), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n520), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n239), .A2(new_n201), .A3(new_n524), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n531), .A2(KEYINPUT30), .A3(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n532), .A3(new_n326), .ZN(new_n533));
  INV_X1    g347(.A(new_n326), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n528), .B(new_n534), .C1(new_n253), .C2(new_n525), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n400), .A2(new_n397), .A3(G210), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n537), .B(KEYINPUT27), .Z(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT26), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n539), .B(new_n224), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT69), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n535), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(KEYINPUT68), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT68), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n535), .A2(new_n547), .A3(new_n544), .ZN(new_n548));
  AND2_X1   g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n326), .B1(new_n526), .B2(new_n529), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n544), .B1(new_n550), .B2(new_n535), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n552), .A3(new_n540), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT29), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT69), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n536), .A2(new_n555), .A3(new_n541), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n543), .A2(new_n553), .A3(new_n554), .A4(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT70), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n550), .A2(new_n558), .A3(new_n535), .ZN(new_n559));
  OAI211_X1 g373(.A(KEYINPUT70), .B(new_n326), .C1(new_n526), .C2(new_n529), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(KEYINPUT28), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n541), .A2(new_n554), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  AND2_X1   g377(.A1(new_n563), .A2(new_n294), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n519), .B1(new_n557), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n546), .A2(new_n548), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n541), .B1(new_n566), .B2(new_n551), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n533), .A2(new_n535), .A3(new_n540), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT31), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT31), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n533), .A2(new_n570), .A3(new_n535), .A4(new_n540), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n567), .A2(new_n569), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT32), .B1(new_n572), .B2(new_n573), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n565), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n518), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n470), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(G101), .ZN(G3));
  AND4_X1   g393(.A1(KEYINPUT85), .A2(new_n292), .A3(new_n293), .A4(new_n294), .ZN(new_n580));
  AOI21_X1  g394(.A(KEYINPUT85), .B1(new_n298), .B2(new_n293), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n306), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n518), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n572), .A2(new_n294), .ZN(new_n584));
  AOI22_X1  g398(.A1(new_n584), .A2(G472), .B1(new_n572), .B2(new_n573), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n582), .A2(new_n583), .A3(new_n189), .A4(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT98), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n307), .A2(KEYINPUT98), .A3(new_n583), .A4(new_n585), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n356), .A2(new_n358), .ZN(new_n591));
  INV_X1    g405(.A(new_n308), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n406), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT33), .B1(new_n388), .B2(KEYINPUT99), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n392), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n595), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n390), .A2(new_n391), .A3(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n394), .A2(G902), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n393), .A2(new_n394), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n467), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n594), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n590), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT34), .B(G104), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G6));
  INV_X1    g421(.A(new_n467), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n396), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n594), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n590), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT100), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT35), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n613), .B(new_n207), .ZN(G9));
  AND3_X1   g428(.A1(new_n582), .A2(new_n189), .A3(new_n308), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n498), .A2(KEYINPUT36), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n492), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n503), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n517), .A2(new_n618), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n615), .A2(new_n469), .A3(new_n585), .A4(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT37), .Z(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G110), .ZN(G12));
  INV_X1    g436(.A(G900), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n403), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n609), .B1(new_n401), .B2(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(new_n565), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n574), .A2(new_n575), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n626), .A2(new_n627), .B1(new_n517), .B2(new_n618), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n592), .B1(new_n356), .B2(new_n358), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n307), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(G128), .ZN(G30));
  NAND2_X1  g446(.A1(new_n624), .A2(new_n401), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT39), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n307), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT40), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n359), .A2(new_n360), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT38), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n396), .A2(new_n467), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n619), .A2(new_n592), .A3(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n639), .B1(KEYINPUT102), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n536), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n541), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n540), .B1(new_n559), .B2(new_n560), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n645), .A2(G902), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n627), .B1(new_n519), .B2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT101), .Z(new_n649));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n641), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n637), .A2(new_n643), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n227), .ZN(G45));
  NAND3_X1  g467(.A1(new_n602), .A2(new_n467), .A3(new_n633), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(KEYINPUT103), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT103), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n602), .A2(new_n467), .A3(new_n656), .A4(new_n633), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n307), .A2(new_n630), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n307), .A2(new_n630), .A3(KEYINPUT104), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G146), .ZN(G48));
  OR2_X1    g479(.A1(new_n298), .A2(new_n293), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n189), .B(new_n666), .C1(new_n580), .C2(new_n581), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT105), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT106), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n300), .A2(KEYINPUT105), .A3(new_n189), .A4(new_n666), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n670), .B1(new_n669), .B2(new_n671), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n577), .B(new_n604), .C1(new_n672), .C2(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT41), .B(G113), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT107), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n674), .B(new_n676), .ZN(G15));
  OAI211_X1 g491(.A(new_n577), .B(new_n610), .C1(new_n672), .C2(new_n673), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G116), .ZN(G18));
  NAND2_X1  g493(.A1(new_n669), .A2(new_n671), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n681), .A2(new_n468), .A3(new_n629), .A4(new_n628), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G119), .ZN(G21));
  AND2_X1   g497(.A1(new_n549), .A2(new_n561), .ZN(new_n684));
  OAI211_X1 g498(.A(new_n569), .B(new_n571), .C1(new_n684), .C2(new_n540), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n573), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n584), .A2(G472), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n594), .A2(new_n518), .A3(new_n640), .A4(new_n688), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n672), .B2(new_n673), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G122), .ZN(G24));
  AND3_X1   g505(.A1(new_n655), .A2(KEYINPUT109), .A3(new_n657), .ZN(new_n692));
  AOI21_X1  g506(.A(KEYINPUT109), .B1(new_n655), .B2(new_n657), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g508(.A1(new_n513), .A2(new_n516), .B1(new_n503), .B2(new_n617), .ZN(new_n695));
  OAI21_X1  g509(.A(KEYINPUT108), .B1(new_n695), .B2(new_n688), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT108), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n685), .A2(new_n573), .B1(new_n584), .B2(G472), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n619), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  AND2_X1   g514(.A1(new_n694), .A2(new_n700), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n629), .A3(new_n669), .A4(new_n671), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G125), .ZN(G27));
  AOI21_X1  g517(.A(new_n592), .B1(new_n359), .B2(new_n360), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n582), .A2(new_n577), .A3(new_n704), .A4(new_n189), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n706), .A2(KEYINPUT42), .A3(new_n694), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT42), .ZN(new_n708));
  INV_X1    g522(.A(new_n694), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n708), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G131), .ZN(G33));
  INV_X1    g526(.A(new_n625), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT110), .B(G134), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G36));
  NAND2_X1  g530(.A1(new_n608), .A2(new_n602), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT43), .ZN(new_n718));
  NOR3_X1   g532(.A1(new_n718), .A2(new_n585), .A3(new_n695), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n720));
  INV_X1    g534(.A(new_n704), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(KEYINPUT44), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n304), .B(KEYINPUT45), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(G469), .A2(G902), .ZN(new_n726));
  AOI21_X1  g540(.A(KEYINPUT46), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n727), .B1(new_n297), .B2(new_n299), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n725), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n190), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(new_n634), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT111), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  OAI211_X1 g548(.A(new_n722), .B(new_n723), .C1(new_n733), .C2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G137), .ZN(G39));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n730), .A2(new_n737), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n738), .A2(new_n739), .A3(new_n721), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n740), .A2(new_n576), .A3(new_n518), .A4(new_n659), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G140), .ZN(G42));
  NOR3_X1   g556(.A1(new_n680), .A2(new_n518), .A3(new_n721), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n743), .A2(new_n402), .A3(new_n649), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n744), .A2(new_n603), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n718), .A2(new_n401), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n680), .A2(new_n721), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(KEYINPUT48), .A3(new_n577), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT48), .ZN(new_n750));
  INV_X1    g564(.A(new_n748), .ZN(new_n751));
  INV_X1    g565(.A(new_n577), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n745), .A2(new_n398), .A3(new_n749), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n300), .A2(new_n666), .ZN(new_n755));
  OAI22_X1  g569(.A1(new_n738), .A2(new_n739), .B1(new_n189), .B2(new_n755), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n747), .A2(new_n518), .A3(new_n688), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(new_n704), .A3(new_n757), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n744), .A2(new_n467), .A3(new_n602), .ZN(new_n759));
  NOR2_X1   g573(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n308), .A2(new_n760), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n639), .A2(new_n681), .A3(new_n757), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(KEYINPUT116), .A2(KEYINPUT50), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n762), .A2(new_n763), .B1(new_n748), .B2(new_n700), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n758), .A2(new_n759), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT117), .ZN(new_n767));
  OR3_X1    g581(.A1(new_n766), .A2(new_n767), .A3(KEYINPUT51), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT51), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT117), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n769), .A2(KEYINPUT117), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n754), .B1(new_n768), .B2(new_n772), .ZN(new_n773));
  AND4_X1   g587(.A1(new_n674), .A2(new_n678), .A3(new_n682), .A4(new_n690), .ZN(new_n774));
  INV_X1    g588(.A(new_n714), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n396), .A2(new_n467), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n628), .A2(new_n776), .A3(new_n633), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n307), .B(new_n704), .C1(new_n701), .C2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT42), .B1(new_n706), .B2(new_n694), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n780));
  OAI211_X1 g594(.A(new_n775), .B(new_n778), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n609), .A2(new_n603), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n638), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n588), .A2(new_n589), .A3(new_n593), .A4(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n784), .A2(new_n578), .A3(new_n620), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n648), .A2(new_n695), .ZN(new_n787));
  AOI211_X1 g601(.A(new_n592), .B(new_n640), .C1(new_n356), .C2(new_n358), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n307), .A2(new_n633), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n664), .A2(new_n631), .A3(new_n702), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(KEYINPUT52), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n702), .A2(new_n631), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n792), .A2(new_n793), .A3(new_n664), .A4(new_n789), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n774), .A2(new_n786), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(KEYINPUT114), .B1(new_n797), .B2(KEYINPUT54), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(KEYINPUT115), .B1(new_n795), .B2(new_n796), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n791), .A2(new_n794), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n714), .B1(new_n707), .B2(new_n710), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n307), .A2(new_n308), .A3(new_n469), .A4(new_n585), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n619), .A2(new_n803), .B1(new_n470), .B2(new_n577), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n802), .A2(new_n804), .A3(new_n778), .A4(new_n784), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n674), .A2(new_n678), .A3(new_n682), .A4(new_n690), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT115), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n801), .A2(new_n807), .A3(new_n808), .A4(KEYINPUT53), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n795), .A2(new_n796), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n800), .A2(new_n809), .A3(new_n810), .A4(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n797), .A2(KEYINPUT114), .A3(KEYINPUT54), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n773), .A2(new_n799), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n681), .A2(new_n629), .A3(new_n757), .ZN(new_n815));
  OAI22_X1  g629(.A1(new_n814), .A2(new_n815), .B1(G952), .B2(G953), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n639), .B1(KEYINPUT49), .B2(new_n755), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT112), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n755), .A2(KEYINPUT49), .ZN(new_n819));
  NOR3_X1   g633(.A1(new_n717), .A2(new_n190), .A3(new_n592), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n819), .A2(new_n583), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n817), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  OAI211_X1 g636(.A(new_n822), .B(new_n649), .C1(new_n818), .C2(new_n821), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(KEYINPUT113), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n816), .A2(new_n824), .ZN(G75));
  NAND3_X1  g639(.A1(new_n800), .A2(new_n811), .A3(new_n809), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(G210), .A3(G902), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT56), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  OR2_X1    g643(.A1(new_n343), .A2(new_n344), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(new_n314), .Z(new_n831));
  XNOR2_X1  g645(.A(new_n831), .B(KEYINPUT55), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n832), .B1(new_n833), .B2(new_n828), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n829), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n397), .A2(G952), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n827), .B(new_n828), .C1(new_n833), .C2(new_n832), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT119), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n835), .A2(new_n841), .A3(new_n838), .A4(new_n837), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(G51));
  NAND2_X1  g657(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(KEYINPUT120), .A3(new_n812), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n826), .A2(new_n846), .A3(KEYINPUT54), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n726), .B(KEYINPUT57), .Z(new_n848));
  NAND3_X1  g662(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n292), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n826), .A2(G469), .A3(G902), .A4(new_n724), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n836), .B1(new_n850), .B2(new_n851), .ZN(G54));
  NAND4_X1  g666(.A1(new_n826), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n853));
  INV_X1    g667(.A(new_n453), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n853), .A2(new_n854), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n856), .A3(new_n836), .ZN(G60));
  NAND2_X1  g671(.A1(G478), .A2(G902), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT59), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n813), .A2(new_n812), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n860), .B2(new_n798), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n596), .A2(new_n598), .ZN(new_n862));
  INV_X1    g676(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n836), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n845), .A2(new_n862), .A3(new_n847), .A4(new_n859), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(G63));
  NAND2_X1  g680(.A1(G217), .A2(G902), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT60), .Z(new_n868));
  NAND2_X1  g682(.A1(new_n826), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n502), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n826), .A2(new_n617), .A3(new_n868), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(KEYINPUT61), .A3(new_n837), .A4(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n873), .A2(KEYINPUT122), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n836), .B1(new_n869), .B2(new_n870), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT122), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT61), .A4(new_n872), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT61), .B1(new_n875), .B2(new_n872), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(KEYINPUT121), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT121), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n881), .B(KEYINPUT61), .C1(new_n875), .C2(new_n872), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n878), .B1(new_n880), .B2(new_n882), .ZN(G66));
  OR2_X1    g697(.A1(new_n806), .A2(new_n785), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n397), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n397), .B1(new_n404), .B2(G224), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n887));
  OR2_X1    g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n887), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n885), .A2(new_n888), .A3(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(G898), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n830), .B1(new_n891), .B2(G953), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n890), .B(new_n892), .Z(G69));
  NAND2_X1  g707(.A1(new_n530), .A2(new_n532), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n418), .ZN(new_n895));
  NAND2_X1  g709(.A1(G900), .A2(G953), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n735), .A2(new_n741), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n577), .B(new_n788), .C1(new_n733), .C2(new_n734), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n802), .B(KEYINPUT127), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n664), .A3(new_n792), .ZN(new_n901));
  OR3_X1    g715(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n895), .B(new_n896), .C1(new_n902), .C2(G953), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n895), .B(KEYINPUT124), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n792), .A2(new_n664), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT62), .ZN(new_n906));
  OR3_X1    g720(.A1(new_n652), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n652), .B2(new_n905), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OR4_X1    g723(.A1(new_n752), .A2(new_n635), .A3(new_n721), .A4(new_n782), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(new_n735), .A3(new_n741), .A4(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n904), .B1(new_n911), .B2(new_n397), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT125), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n903), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(G953), .B1(new_n279), .B2(new_n623), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT126), .Z(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n916), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n903), .B(new_n918), .C1(new_n914), .C2(new_n915), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(G72));
  NAND2_X1  g736(.A1(G472), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT63), .Z(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n902), .B2(new_n884), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n925), .A2(new_n541), .A3(new_n644), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n911), .B2(new_n884), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n836), .B1(new_n927), .B2(new_n645), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n543), .A2(new_n568), .A3(new_n556), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n797), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n926), .A2(new_n928), .A3(new_n930), .ZN(G57));
endmodule


