

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720;

  NOR2_X1 U369 ( .A1(n617), .A2(n613), .ZN(n638) );
  INV_X1 U370 ( .A(KEYINPUT23), .ZN(n409) );
  OR2_X2 U371 ( .A1(n683), .A2(G902), .ZN(n417) );
  XNOR2_X2 U372 ( .A(n698), .B(G146), .ZN(n486) );
  XNOR2_X2 U373 ( .A(n442), .B(n365), .ZN(n698) );
  XNOR2_X1 U374 ( .A(G143), .B(G128), .ZN(n418) );
  NOR2_X1 U375 ( .A1(n597), .A2(n685), .ZN(n355) );
  NAND2_X1 U376 ( .A1(n362), .A2(n359), .ZN(n364) );
  NAND2_X1 U377 ( .A1(n384), .A2(n350), .ZN(n702) );
  INV_X1 U378 ( .A(n688), .ZN(n362) );
  XNOR2_X1 U379 ( .A(n525), .B(n524), .ZN(n688) );
  NAND2_X1 U380 ( .A1(n392), .A2(n523), .ZN(n525) );
  XNOR2_X1 U381 ( .A(n506), .B(n372), .ZN(n716) );
  XNOR2_X1 U382 ( .A(n501), .B(n500), .ZN(n649) );
  XNOR2_X1 U383 ( .A(n537), .B(n463), .ZN(n559) );
  XNOR2_X1 U384 ( .A(n479), .B(n416), .ZN(n415) );
  XNOR2_X1 U385 ( .A(n406), .B(n403), .ZN(n476) );
  XNOR2_X1 U386 ( .A(n448), .B(KEYINPUT20), .ZN(n478) );
  XNOR2_X1 U387 ( .A(n453), .B(n387), .ZN(n699) );
  XNOR2_X1 U388 ( .A(n408), .B(n407), .ZN(n406) );
  XNOR2_X1 U389 ( .A(n418), .B(n370), .ZN(n455) );
  XNOR2_X1 U390 ( .A(n409), .B(KEYINPUT24), .ZN(n408) );
  XNOR2_X1 U391 ( .A(G128), .B(KEYINPUT73), .ZN(n407) );
  XOR2_X1 U392 ( .A(G104), .B(G110), .Z(n480) );
  XNOR2_X1 U393 ( .A(n477), .B(n699), .ZN(n683) );
  XNOR2_X1 U394 ( .A(n476), .B(n475), .ZN(n477) );
  NOR2_X1 U395 ( .A1(n676), .A2(n685), .ZN(n677) );
  INV_X1 U396 ( .A(n702), .ZN(n359) );
  NOR2_X1 U397 ( .A1(n665), .A2(n685), .ZN(n666) );
  XNOR2_X1 U398 ( .A(n388), .B(G125), .ZN(n453) );
  INV_X1 U399 ( .A(G146), .ZN(n388) );
  NAND2_X1 U400 ( .A1(n715), .A2(n606), .ZN(n382) );
  INV_X1 U401 ( .A(n716), .ZN(n371) );
  XNOR2_X1 U402 ( .A(n367), .B(n428), .ZN(n365) );
  XNOR2_X1 U403 ( .A(n369), .B(n368), .ZN(n367) );
  INV_X1 U404 ( .A(KEYINPUT4), .ZN(n368) );
  OR2_X1 U405 ( .A1(G237), .A2(G902), .ZN(n459) );
  INV_X1 U406 ( .A(G469), .ZN(n487) );
  NOR2_X1 U407 ( .A1(G902), .A2(n667), .ZN(n488) );
  XNOR2_X1 U408 ( .A(n379), .B(n378), .ZN(n452) );
  XNOR2_X1 U409 ( .A(G119), .B(G116), .ZN(n378) );
  XNOR2_X1 U410 ( .A(n419), .B(G113), .ZN(n379) );
  XNOR2_X1 U411 ( .A(G101), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U412 ( .A(n455), .B(G134), .ZN(n442) );
  XOR2_X1 U413 ( .A(G122), .B(G107), .Z(n449) );
  XNOR2_X1 U414 ( .A(KEYINPUT10), .B(G140), .ZN(n387) );
  NAND2_X1 U415 ( .A1(n371), .A2(n394), .ZN(n393) );
  XNOR2_X1 U416 ( .A(n382), .B(n495), .ZN(n507) );
  XNOR2_X1 U417 ( .A(n376), .B(KEYINPUT21), .ZN(n375) );
  NAND2_X1 U418 ( .A1(n478), .A2(G221), .ZN(n377) );
  INV_X1 U419 ( .A(KEYINPUT93), .ZN(n376) );
  NOR2_X1 U420 ( .A1(G953), .A2(G237), .ZN(n429) );
  XNOR2_X1 U421 ( .A(n366), .B(G131), .ZN(n428) );
  INV_X1 U422 ( .A(KEYINPUT70), .ZN(n366) );
  NAND2_X1 U423 ( .A1(n625), .A2(n357), .ZN(n516) );
  XNOR2_X1 U424 ( .A(n353), .B(KEYINPUT81), .ZN(n545) );
  OR2_X1 U425 ( .A1(n528), .A2(n529), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n391), .B(n390), .ZN(n511) );
  XNOR2_X1 U427 ( .A(n436), .B(G475), .ZN(n390) );
  OR2_X1 U428 ( .A1(n673), .A2(G902), .ZN(n391) );
  XNOR2_X1 U429 ( .A(G116), .B(KEYINPUT98), .ZN(n439) );
  XOR2_X1 U430 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n440) );
  XOR2_X1 U431 ( .A(G143), .B(KEYINPUT95), .Z(n431) );
  XNOR2_X1 U432 ( .A(G113), .B(KEYINPUT12), .ZN(n425) );
  XOR2_X1 U433 ( .A(KEYINPUT11), .B(G122), .Z(n426) );
  INV_X1 U434 ( .A(KEYINPUT79), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n400), .B(KEYINPUT78), .ZN(n399) );
  INV_X1 U436 ( .A(KEYINPUT18), .ZN(n400) );
  XNOR2_X1 U437 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U438 ( .A(n453), .B(n454), .ZN(n401) );
  NOR2_X1 U439 ( .A1(n649), .A2(n502), .ZN(n503) );
  XNOR2_X1 U440 ( .A(n460), .B(KEYINPUT80), .ZN(n461) );
  XNOR2_X1 U441 ( .A(n552), .B(n358), .ZN(n491) );
  INV_X1 U442 ( .A(KEYINPUT1), .ZN(n358) );
  XNOR2_X1 U443 ( .A(n511), .B(n389), .ZN(n514) );
  INV_X1 U444 ( .A(KEYINPUT97), .ZN(n389) );
  INV_X1 U445 ( .A(KEYINPUT94), .ZN(n413) );
  XNOR2_X1 U446 ( .A(n515), .B(KEYINPUT90), .ZN(n502) );
  INV_X1 U447 ( .A(KEYINPUT25), .ZN(n416) );
  NOR2_X1 U448 ( .A1(n534), .A2(n493), .ZN(n508) );
  INV_X1 U449 ( .A(n491), .ZN(n357) );
  XNOR2_X1 U450 ( .A(n451), .B(n452), .ZN(n687) );
  INV_X1 U451 ( .A(KEYINPUT44), .ZN(n394) );
  XNOR2_X1 U452 ( .A(KEYINPUT71), .B(G137), .ZN(n369) );
  AND2_X1 U453 ( .A1(n348), .A2(n609), .ZN(n579) );
  XNOR2_X1 U454 ( .A(n465), .B(n464), .ZN(n467) );
  NAND2_X1 U455 ( .A1(G234), .A2(G237), .ZN(n464) );
  XOR2_X1 U456 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n465) );
  INV_X1 U457 ( .A(KEYINPUT48), .ZN(n385) );
  INV_X1 U458 ( .A(KEYINPUT68), .ZN(n496) );
  XNOR2_X1 U459 ( .A(n486), .B(n423), .ZN(n593) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n403) );
  XNOR2_X1 U461 ( .A(G137), .B(G119), .ZN(n405) );
  XNOR2_X1 U462 ( .A(G110), .B(KEYINPUT91), .ZN(n404) );
  XNOR2_X1 U463 ( .A(G140), .B(G107), .ZN(n484) );
  INV_X1 U464 ( .A(KEYINPUT2), .ZN(n363) );
  XNOR2_X1 U465 ( .A(n547), .B(KEYINPUT77), .ZN(n575) );
  AND2_X1 U466 ( .A1(n661), .A2(G472), .ZN(n592) );
  XNOR2_X1 U467 ( .A(n443), .B(n354), .ZN(n679) );
  XNOR2_X1 U468 ( .A(n444), .B(n445), .ZN(n354) );
  XNOR2_X1 U469 ( .A(n435), .B(n434), .ZN(n673) );
  XNOR2_X1 U470 ( .A(n699), .B(n427), .ZN(n435) );
  XNOR2_X1 U471 ( .A(n455), .B(n456), .ZN(n457) );
  XNOR2_X1 U472 ( .A(n401), .B(n397), .ZN(n456) );
  XNOR2_X1 U473 ( .A(n399), .B(n398), .ZN(n397) );
  NOR2_X1 U474 ( .A1(G952), .A2(n703), .ZN(n685) );
  NOR2_X1 U475 ( .A1(n586), .A2(n585), .ZN(n619) );
  XNOR2_X1 U476 ( .A(n402), .B(n352), .ZN(n713) );
  XNOR2_X1 U477 ( .A(n396), .B(KEYINPUT86), .ZN(n372) );
  INV_X1 U478 ( .A(KEYINPUT35), .ZN(n396) );
  XNOR2_X1 U479 ( .A(n490), .B(n383), .ZN(n715) );
  XNOR2_X1 U480 ( .A(KEYINPUT32), .B(KEYINPUT64), .ZN(n383) );
  XNOR2_X1 U481 ( .A(n512), .B(KEYINPUT100), .ZN(n617) );
  AND2_X1 U482 ( .A1(n513), .A2(n514), .ZN(n512) );
  NOR2_X1 U483 ( .A1(n561), .A2(n560), .ZN(n611) );
  NOR2_X1 U484 ( .A1(n514), .A2(n513), .ZN(n613) );
  INV_X1 U485 ( .A(n502), .ZN(n518) );
  XNOR2_X1 U486 ( .A(n381), .B(n471), .ZN(n515) );
  INV_X1 U487 ( .A(n515), .ZN(n380) );
  NOR2_X1 U488 ( .A1(n584), .A2(n357), .ZN(n347) );
  XNOR2_X1 U489 ( .A(n377), .B(n375), .ZN(n530) );
  AND2_X1 U490 ( .A1(n574), .A2(n573), .ZN(n348) );
  AND2_X1 U491 ( .A1(n373), .A2(n579), .ZN(n349) );
  AND2_X1 U492 ( .A1(n720), .A2(n587), .ZN(n350) );
  AND2_X1 U493 ( .A1(n472), .A2(n621), .ZN(n351) );
  XOR2_X1 U494 ( .A(KEYINPUT106), .B(KEYINPUT40), .Z(n352) );
  XNOR2_X1 U495 ( .A(G902), .B(KEYINPUT15), .ZN(n458) );
  XNOR2_X2 U496 ( .A(n548), .B(KEYINPUT39), .ZN(n580) );
  NOR2_X1 U497 ( .A1(n702), .A2(n363), .ZN(n360) );
  XNOR2_X1 U498 ( .A(n386), .B(n385), .ZN(n384) );
  NOR2_X1 U499 ( .A1(KEYINPUT83), .A2(n566), .ZN(n567) );
  NOR2_X1 U500 ( .A1(n569), .A2(n568), .ZN(n574) );
  NAND2_X1 U501 ( .A1(n362), .A2(n360), .ZN(n661) );
  AND2_X1 U502 ( .A1(n661), .A2(G475), .ZN(n411) );
  INV_X1 U503 ( .A(n582), .ZN(n583) );
  XNOR2_X1 U504 ( .A(n536), .B(KEYINPUT103), .ZN(n582) );
  NAND2_X1 U505 ( .A1(n374), .A2(n349), .ZN(n386) );
  XNOR2_X1 U506 ( .A(n355), .B(n598), .ZN(G57) );
  AND2_X1 U507 ( .A1(n491), .A2(n356), .ZN(n626) );
  INV_X1 U508 ( .A(n625), .ZN(n356) );
  NOR2_X1 U509 ( .A1(n509), .A2(n357), .ZN(n510) );
  NAND2_X1 U510 ( .A1(n539), .A2(n357), .ZN(n540) );
  NAND2_X1 U511 ( .A1(n362), .A2(n361), .ZN(n591) );
  NOR2_X1 U512 ( .A1(n702), .A2(n458), .ZN(n361) );
  XNOR2_X1 U513 ( .A(n364), .B(n363), .ZN(n654) );
  INV_X1 U514 ( .A(n717), .ZN(n373) );
  XNOR2_X1 U515 ( .A(n558), .B(KEYINPUT46), .ZN(n374) );
  NAND2_X1 U516 ( .A1(n380), .A2(n351), .ZN(n473) );
  NAND2_X1 U517 ( .A1(n559), .A2(n470), .ZN(n381) );
  NAND2_X1 U518 ( .A1(n395), .A2(n393), .ZN(n392) );
  NAND2_X1 U519 ( .A1(n507), .A2(n716), .ZN(n395) );
  NOR2_X2 U520 ( .A1(n713), .A2(n712), .ZN(n558) );
  NAND2_X1 U521 ( .A1(n580), .A2(n613), .ZN(n402) );
  AND2_X1 U522 ( .A1(n662), .A2(n661), .ZN(n681) );
  NAND2_X1 U523 ( .A1(n662), .A2(n410), .ZN(n663) );
  AND2_X1 U524 ( .A1(n661), .A2(G210), .ZN(n410) );
  NAND2_X1 U525 ( .A1(n662), .A2(n411), .ZN(n674) );
  NAND2_X1 U526 ( .A1(n412), .A2(n546), .ZN(n547) );
  XNOR2_X1 U527 ( .A(n541), .B(KEYINPUT104), .ZN(n412) );
  XNOR2_X2 U528 ( .A(n414), .B(n413), .ZN(n541) );
  NAND2_X1 U529 ( .A1(n625), .A2(n552), .ZN(n414) );
  XNOR2_X2 U530 ( .A(n417), .B(n415), .ZN(n620) );
  INV_X1 U531 ( .A(n620), .ZN(n532) );
  XNOR2_X1 U532 ( .A(n499), .B(KEYINPUT33), .ZN(n500) );
  XNOR2_X1 U533 ( .A(n452), .B(n422), .ZN(n423) );
  INV_X1 U534 ( .A(n619), .ZN(n587) );
  INV_X1 U535 ( .A(KEYINPUT45), .ZN(n524) );
  NAND2_X1 U536 ( .A1(n634), .A2(n586), .ZN(n537) );
  XNOR2_X1 U537 ( .A(n687), .B(n457), .ZN(n660) );
  XNOR2_X1 U538 ( .A(n594), .B(KEYINPUT62), .ZN(n595) );
  XNOR2_X1 U539 ( .A(n596), .B(n595), .ZN(n597) );
  INV_X1 U540 ( .A(KEYINPUT63), .ZN(n598) );
  INV_X2 U541 ( .A(G953), .ZN(n703) );
  XOR2_X1 U542 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n421) );
  NAND2_X1 U543 ( .A1(n429), .A2(G210), .ZN(n420) );
  XNOR2_X1 U544 ( .A(n421), .B(n420), .ZN(n422) );
  NOR2_X1 U545 ( .A1(n593), .A2(G902), .ZN(n424) );
  XNOR2_X1 U546 ( .A(G472), .B(n424), .ZN(n549) );
  INV_X2 U547 ( .A(n549), .ZN(n542) );
  XOR2_X1 U548 ( .A(KEYINPUT6), .B(n542), .Z(n534) );
  XNOR2_X1 U549 ( .A(KEYINPUT96), .B(KEYINPUT13), .ZN(n436) );
  XNOR2_X1 U550 ( .A(n426), .B(n425), .ZN(n427) );
  XNOR2_X1 U551 ( .A(n428), .B(G104), .ZN(n433) );
  NAND2_X1 U552 ( .A1(G214), .A2(n429), .ZN(n430) );
  XNOR2_X1 U553 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U554 ( .A(n433), .B(n432), .ZN(n434) );
  NAND2_X1 U555 ( .A1(n703), .A2(G234), .ZN(n438) );
  XNOR2_X1 U556 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n437) );
  XNOR2_X1 U557 ( .A(n438), .B(n437), .ZN(n474) );
  NAND2_X1 U558 ( .A1(n474), .A2(G217), .ZN(n445) );
  XNOR2_X1 U559 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U560 ( .A(n441), .B(KEYINPUT99), .Z(n444) );
  XNOR2_X1 U561 ( .A(n442), .B(n449), .ZN(n443) );
  NOR2_X1 U562 ( .A1(G902), .A2(n679), .ZN(n446) );
  XOR2_X1 U563 ( .A(G478), .B(n446), .Z(n513) );
  INV_X1 U564 ( .A(n513), .ZN(n504) );
  NAND2_X1 U565 ( .A1(n511), .A2(n504), .ZN(n636) );
  INV_X1 U566 ( .A(n636), .ZN(n472) );
  NAND2_X1 U567 ( .A1(n458), .A2(G234), .ZN(n447) );
  XNOR2_X1 U568 ( .A(n447), .B(KEYINPUT92), .ZN(n448) );
  NAND2_X1 U569 ( .A1(G214), .A2(n459), .ZN(n634) );
  XNOR2_X1 U570 ( .A(KEYINPUT16), .B(n480), .ZN(n450) );
  XNOR2_X1 U571 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U572 ( .A1(G224), .A2(n703), .ZN(n454) );
  INV_X1 U573 ( .A(n458), .ZN(n588) );
  NOR2_X1 U574 ( .A1(n660), .A2(n588), .ZN(n462) );
  NAND2_X1 U575 ( .A1(G210), .A2(n459), .ZN(n460) );
  XNOR2_X2 U576 ( .A(n462), .B(n461), .ZN(n586) );
  XNOR2_X1 U577 ( .A(KEYINPUT19), .B(KEYINPUT66), .ZN(n463) );
  NOR2_X1 U578 ( .A1(G898), .A2(n703), .ZN(n686) );
  NAND2_X1 U579 ( .A1(n467), .A2(G902), .ZN(n466) );
  XNOR2_X1 U580 ( .A(n466), .B(KEYINPUT89), .ZN(n526) );
  NAND2_X1 U581 ( .A1(n686), .A2(n526), .ZN(n469) );
  NAND2_X1 U582 ( .A1(G952), .A2(n467), .ZN(n647) );
  NOR2_X1 U583 ( .A1(G953), .A2(n647), .ZN(n529) );
  INV_X1 U584 ( .A(n529), .ZN(n468) );
  NAND2_X1 U585 ( .A1(n469), .A2(n468), .ZN(n470) );
  XOR2_X1 U586 ( .A(KEYINPUT67), .B(KEYINPUT0), .Z(n471) );
  XNOR2_X1 U587 ( .A(n473), .B(KEYINPUT22), .ZN(n493) );
  NAND2_X1 U588 ( .A1(G221), .A2(n474), .ZN(n475) );
  NAND2_X1 U589 ( .A1(G217), .A2(n478), .ZN(n479) );
  XOR2_X1 U590 ( .A(G101), .B(n480), .Z(n482) );
  NAND2_X1 U591 ( .A1(G227), .A2(n703), .ZN(n481) );
  XNOR2_X1 U592 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U593 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U594 ( .A(n486), .B(n485), .ZN(n667) );
  XNOR2_X2 U595 ( .A(n488), .B(n487), .ZN(n552) );
  NOR2_X1 U596 ( .A1(n620), .A2(n491), .ZN(n489) );
  NAND2_X1 U597 ( .A1(n508), .A2(n489), .ZN(n490) );
  NAND2_X1 U598 ( .A1(n532), .A2(n491), .ZN(n492) );
  NOR2_X1 U599 ( .A1(n493), .A2(n492), .ZN(n494) );
  INV_X1 U600 ( .A(n542), .ZN(n624) );
  NAND2_X1 U601 ( .A1(n494), .A2(n624), .ZN(n606) );
  NOR2_X1 U602 ( .A1(KEYINPUT44), .A2(KEYINPUT87), .ZN(n495) );
  INV_X1 U603 ( .A(n530), .ZN(n621) );
  NAND2_X1 U604 ( .A1(n620), .A2(n621), .ZN(n497) );
  XNOR2_X2 U605 ( .A(n497), .B(n496), .ZN(n625) );
  INV_X1 U606 ( .A(n516), .ZN(n498) );
  NAND2_X1 U607 ( .A1(n498), .A2(n534), .ZN(n501) );
  XOR2_X1 U608 ( .A(KEYINPUT74), .B(KEYINPUT102), .Z(n499) );
  XNOR2_X1 U609 ( .A(n503), .B(KEYINPUT34), .ZN(n505) );
  NOR2_X1 U610 ( .A1(n511), .A2(n504), .ZN(n577) );
  NAND2_X1 U611 ( .A1(n505), .A2(n577), .ZN(n506) );
  NAND2_X1 U612 ( .A1(n508), .A2(n620), .ZN(n509) );
  XOR2_X1 U613 ( .A(KEYINPUT101), .B(n510), .Z(n714) );
  XNOR2_X1 U614 ( .A(n638), .B(KEYINPUT85), .ZN(n564) );
  INV_X1 U615 ( .A(n564), .ZN(n521) );
  NOR2_X1 U616 ( .A1(n624), .A2(n516), .ZN(n630) );
  NAND2_X1 U617 ( .A1(n380), .A2(n630), .ZN(n517) );
  XNOR2_X1 U618 ( .A(n517), .B(KEYINPUT31), .ZN(n616) );
  NAND2_X1 U619 ( .A1(n518), .A2(n541), .ZN(n519) );
  NOR2_X1 U620 ( .A1(n542), .A2(n519), .ZN(n601) );
  NOR2_X1 U621 ( .A1(n616), .A2(n601), .ZN(n520) );
  NOR2_X1 U622 ( .A1(n521), .A2(n520), .ZN(n522) );
  NOR2_X1 U623 ( .A1(n714), .A2(n522), .ZN(n523) );
  NAND2_X1 U624 ( .A1(G953), .A2(n526), .ZN(n527) );
  NOR2_X1 U625 ( .A1(G900), .A2(n527), .ZN(n528) );
  NOR2_X1 U626 ( .A1(n545), .A2(n530), .ZN(n531) );
  NAND2_X1 U627 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U628 ( .A(KEYINPUT72), .B(n533), .ZN(n550) );
  NAND2_X1 U629 ( .A1(n613), .A2(n534), .ZN(n535) );
  NOR2_X1 U630 ( .A1(n550), .A2(n535), .ZN(n536) );
  NOR2_X1 U631 ( .A1(n582), .A2(n537), .ZN(n538) );
  XNOR2_X1 U632 ( .A(KEYINPUT36), .B(n538), .ZN(n539) );
  XNOR2_X1 U633 ( .A(n540), .B(KEYINPUT109), .ZN(n717) );
  NAND2_X1 U634 ( .A1(n542), .A2(n634), .ZN(n543) );
  XNOR2_X1 U635 ( .A(KEYINPUT30), .B(n543), .ZN(n544) );
  NOR2_X1 U636 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U637 ( .A(KEYINPUT38), .B(n586), .Z(n633) );
  NAND2_X1 U638 ( .A1(n575), .A2(n633), .ZN(n548) );
  XOR2_X1 U639 ( .A(KEYINPUT108), .B(KEYINPUT42), .Z(n557) );
  NOR2_X1 U640 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U641 ( .A(KEYINPUT28), .B(n551), .ZN(n553) );
  NAND2_X1 U642 ( .A1(n553), .A2(n552), .ZN(n560) );
  NAND2_X1 U643 ( .A1(n634), .A2(n633), .ZN(n637) );
  NOR2_X1 U644 ( .A1(n636), .A2(n637), .ZN(n555) );
  XNOR2_X1 U645 ( .A(KEYINPUT41), .B(KEYINPUT107), .ZN(n554) );
  XOR2_X1 U646 ( .A(n555), .B(n554), .Z(n650) );
  OR2_X1 U647 ( .A1(n560), .A2(n650), .ZN(n556) );
  XNOR2_X1 U648 ( .A(n557), .B(n556), .ZN(n712) );
  INV_X1 U649 ( .A(n559), .ZN(n561) );
  NAND2_X1 U650 ( .A1(KEYINPUT83), .A2(n611), .ZN(n563) );
  OR2_X1 U651 ( .A1(n638), .A2(KEYINPUT84), .ZN(n562) );
  NAND2_X1 U652 ( .A1(n563), .A2(n562), .ZN(n569) );
  NAND2_X1 U653 ( .A1(n611), .A2(n564), .ZN(n565) );
  NAND2_X1 U654 ( .A1(KEYINPUT84), .A2(n565), .ZN(n566) );
  NOR2_X1 U655 ( .A1(KEYINPUT47), .A2(n567), .ZN(n568) );
  OR2_X1 U656 ( .A1(n611), .A2(KEYINPUT83), .ZN(n571) );
  NAND2_X1 U657 ( .A1(KEYINPUT84), .A2(n638), .ZN(n570) );
  NAND2_X1 U658 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U659 ( .A1(n572), .A2(KEYINPUT47), .ZN(n573) );
  NAND2_X1 U660 ( .A1(n575), .A2(n586), .ZN(n576) );
  XNOR2_X1 U661 ( .A(KEYINPUT105), .B(n576), .ZN(n578) );
  NAND2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n609) );
  NAND2_X1 U663 ( .A1(n617), .A2(n580), .ZN(n581) );
  XNOR2_X1 U664 ( .A(n581), .B(KEYINPUT110), .ZN(n720) );
  NAND2_X1 U665 ( .A1(n583), .A2(n634), .ZN(n584) );
  XNOR2_X1 U666 ( .A(n347), .B(KEYINPUT43), .ZN(n585) );
  NAND2_X1 U667 ( .A1(n588), .A2(KEYINPUT2), .ZN(n589) );
  XOR2_X1 U668 ( .A(KEYINPUT65), .B(n589), .Z(n590) );
  NAND2_X2 U669 ( .A1(n591), .A2(n590), .ZN(n662) );
  NAND2_X1 U670 ( .A1(n592), .A2(n662), .ZN(n596) );
  XOR2_X1 U671 ( .A(n593), .B(KEYINPUT111), .Z(n594) );
  NAND2_X1 U672 ( .A1(n601), .A2(n613), .ZN(n599) );
  XNOR2_X1 U673 ( .A(n599), .B(KEYINPUT112), .ZN(n600) );
  XNOR2_X1 U674 ( .A(G104), .B(n600), .ZN(G6) );
  XOR2_X1 U675 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n603) );
  NAND2_X1 U676 ( .A1(n601), .A2(n617), .ZN(n602) );
  XNOR2_X1 U677 ( .A(n603), .B(n602), .ZN(n605) );
  XOR2_X1 U678 ( .A(G107), .B(KEYINPUT27), .Z(n604) );
  XNOR2_X1 U679 ( .A(n605), .B(n604), .ZN(G9) );
  XNOR2_X1 U680 ( .A(G110), .B(n606), .ZN(G12) );
  XOR2_X1 U681 ( .A(G128), .B(KEYINPUT29), .Z(n608) );
  NAND2_X1 U682 ( .A1(n611), .A2(n617), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n608), .B(n607), .ZN(G30) );
  XNOR2_X1 U684 ( .A(G143), .B(KEYINPUT114), .ZN(n610) );
  XNOR2_X1 U685 ( .A(n610), .B(n609), .ZN(G45) );
  NAND2_X1 U686 ( .A1(n611), .A2(n613), .ZN(n612) );
  XNOR2_X1 U687 ( .A(n612), .B(G146), .ZN(G48) );
  XOR2_X1 U688 ( .A(G113), .B(KEYINPUT115), .Z(n615) );
  NAND2_X1 U689 ( .A1(n616), .A2(n613), .ZN(n614) );
  XNOR2_X1 U690 ( .A(n615), .B(n614), .ZN(G15) );
  NAND2_X1 U691 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U692 ( .A(n618), .B(G116), .ZN(G18) );
  XOR2_X1 U693 ( .A(G140), .B(n619), .Z(G42) );
  NOR2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  XNOR2_X1 U695 ( .A(n622), .B(KEYINPUT49), .ZN(n623) );
  NAND2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n628) );
  XNOR2_X1 U697 ( .A(n626), .B(KEYINPUT50), .ZN(n627) );
  NOR2_X1 U698 ( .A1(n628), .A2(n627), .ZN(n629) );
  NOR2_X1 U699 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U700 ( .A(KEYINPUT51), .B(n631), .Z(n632) );
  NOR2_X1 U701 ( .A1(n650), .A2(n632), .ZN(n644) );
  NOR2_X1 U702 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U703 ( .A1(n636), .A2(n635), .ZN(n641) );
  NOR2_X1 U704 ( .A1(n638), .A2(n637), .ZN(n639) );
  XOR2_X1 U705 ( .A(KEYINPUT117), .B(n639), .Z(n640) );
  NOR2_X1 U706 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U707 ( .A1(n642), .A2(n649), .ZN(n643) );
  NOR2_X1 U708 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U709 ( .A(n645), .B(KEYINPUT52), .ZN(n646) );
  NOR2_X1 U710 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U711 ( .A(n648), .B(KEYINPUT118), .ZN(n652) );
  NOR2_X1 U712 ( .A1(n650), .A2(n649), .ZN(n651) );
  NOR2_X1 U713 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U714 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U715 ( .A1(n655), .A2(G953), .ZN(n656) );
  XNOR2_X1 U716 ( .A(n656), .B(KEYINPUT53), .ZN(G75) );
  XOR2_X1 U717 ( .A(KEYINPUT88), .B(KEYINPUT82), .Z(n658) );
  XNOR2_X1 U718 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n657) );
  XNOR2_X1 U719 ( .A(n658), .B(n657), .ZN(n659) );
  XNOR2_X1 U720 ( .A(n660), .B(n659), .ZN(n664) );
  XNOR2_X1 U721 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U722 ( .A(n666), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U723 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n669) );
  XNOR2_X1 U724 ( .A(n667), .B(KEYINPUT57), .ZN(n668) );
  XNOR2_X1 U725 ( .A(n669), .B(n668), .ZN(n671) );
  NAND2_X1 U726 ( .A1(n681), .A2(G469), .ZN(n670) );
  XNOR2_X1 U727 ( .A(n671), .B(n670), .ZN(n672) );
  NOR2_X1 U728 ( .A1(n685), .A2(n672), .ZN(G54) );
  XOR2_X1 U729 ( .A(n673), .B(KEYINPUT59), .Z(n675) );
  XNOR2_X1 U730 ( .A(n675), .B(n674), .ZN(n676) );
  XNOR2_X1 U731 ( .A(n677), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U732 ( .A1(G478), .A2(n681), .ZN(n678) );
  XNOR2_X1 U733 ( .A(n679), .B(n678), .ZN(n680) );
  NOR2_X1 U734 ( .A1(n685), .A2(n680), .ZN(G63) );
  NAND2_X1 U735 ( .A1(G217), .A2(n681), .ZN(n682) );
  XNOR2_X1 U736 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U737 ( .A1(n685), .A2(n684), .ZN(G66) );
  XNOR2_X1 U738 ( .A(KEYINPUT122), .B(KEYINPUT121), .ZN(n697) );
  NOR2_X1 U739 ( .A1(n687), .A2(n686), .ZN(n695) );
  NOR2_X1 U740 ( .A1(G953), .A2(n688), .ZN(n689) );
  XOR2_X1 U741 ( .A(KEYINPUT120), .B(n689), .Z(n693) );
  NAND2_X1 U742 ( .A1(G953), .A2(G224), .ZN(n690) );
  XNOR2_X1 U743 ( .A(KEYINPUT61), .B(n690), .ZN(n691) );
  NAND2_X1 U744 ( .A1(n691), .A2(G898), .ZN(n692) );
  NAND2_X1 U745 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U746 ( .A(n695), .B(n694), .Z(n696) );
  XNOR2_X1 U747 ( .A(n697), .B(n696), .ZN(G69) );
  XNOR2_X1 U748 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n701) );
  XNOR2_X1 U749 ( .A(n698), .B(n699), .ZN(n700) );
  XNOR2_X1 U750 ( .A(n701), .B(n700), .ZN(n705) );
  XNOR2_X1 U751 ( .A(n702), .B(n705), .ZN(n704) );
  NAND2_X1 U752 ( .A1(n704), .A2(n703), .ZN(n710) );
  XNOR2_X1 U753 ( .A(G227), .B(n705), .ZN(n706) );
  NAND2_X1 U754 ( .A1(n706), .A2(G900), .ZN(n707) );
  NAND2_X1 U755 ( .A1(n707), .A2(G953), .ZN(n708) );
  XOR2_X1 U756 ( .A(KEYINPUT125), .B(n708), .Z(n709) );
  NAND2_X1 U757 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U758 ( .A(KEYINPUT126), .B(n711), .ZN(G72) );
  XOR2_X1 U759 ( .A(G137), .B(n712), .Z(G39) );
  XOR2_X1 U760 ( .A(n713), .B(G131), .Z(G33) );
  XOR2_X1 U761 ( .A(G101), .B(n714), .Z(G3) );
  XNOR2_X1 U762 ( .A(G119), .B(n715), .ZN(G21) );
  XNOR2_X1 U763 ( .A(G122), .B(n716), .ZN(G24) );
  XNOR2_X1 U764 ( .A(n717), .B(KEYINPUT116), .ZN(n718) );
  XNOR2_X1 U765 ( .A(n718), .B(KEYINPUT37), .ZN(n719) );
  XNOR2_X1 U766 ( .A(G125), .B(n719), .ZN(G27) );
  XNOR2_X1 U767 ( .A(G134), .B(n720), .ZN(G36) );
endmodule

