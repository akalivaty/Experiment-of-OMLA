//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n569, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT65), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT66), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT68), .Z(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n460), .B1(new_n461), .B2(G2106), .ZN(G319));
  INV_X1    g037(.A(G113), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  OR3_X1    g039(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT69), .ZN(new_n465));
  OAI21_X1  g040(.A(KEYINPUT69), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n465), .B(new_n466), .C1(new_n467), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n470), .A2(G2105), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n464), .A2(G2105), .ZN(new_n474));
  AOI22_X1  g049(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NOR2_X1   g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  XNOR2_X1  g053(.A(new_n478), .B(KEYINPUT70), .ZN(new_n479));
  INV_X1    g054(.A(G2105), .ZN(new_n480));
  OAI211_X1 g055(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n473), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n470), .A2(new_n480), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n481), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  OAI211_X1 g061(.A(G138), .B(new_n480), .C1(new_n468), .C2(new_n469), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT4), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n489), .A2(new_n480), .A3(G138), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT71), .B1(new_n470), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g066(.A(KEYINPUT3), .B(G2104), .ZN(new_n492));
  AND3_X1   g067(.A1(new_n489), .A2(new_n480), .A3(G138), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT71), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n488), .A2(new_n491), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(G114), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(G2105), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n499), .B1(new_n483), .B2(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT72), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT5), .ZN(new_n504));
  OAI21_X1  g079(.A(new_n503), .B1(new_n504), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n506), .A2(KEYINPUT72), .A3(KEYINPUT5), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n505), .A2(new_n507), .B1(new_n504), .B2(G543), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT6), .B(G651), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n508), .A2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(G543), .ZN(new_n515));
  INV_X1    g090(.A(G50), .ZN(new_n516));
  OAI22_X1  g091(.A1(new_n513), .A2(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n511), .A2(new_n517), .ZN(G166));
  INV_X1    g093(.A(new_n515), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n519), .A2(G51), .B1(new_n508), .B2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n508), .A2(G89), .A3(new_n512), .ZN(new_n523));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(KEYINPUT73), .ZN(new_n527));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n523), .A2(new_n528), .A3(new_n525), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n522), .B1(new_n527), .B2(new_n529), .ZN(G168));
  AND2_X1   g105(.A1(new_n508), .A2(new_n512), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n531), .A2(G90), .B1(G52), .B2(new_n519), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n508), .A2(G64), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G651), .ZN(new_n536));
  NAND3_X1  g111(.A1(new_n532), .A2(new_n536), .A3(KEYINPUT74), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n538));
  INV_X1    g113(.A(G90), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n513), .A2(new_n539), .B1(new_n515), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n510), .B1(new_n533), .B2(new_n534), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n538), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n537), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n508), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n510), .ZN(new_n546));
  INV_X1    g121(.A(G81), .ZN(new_n547));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  OAI22_X1  g123(.A1(new_n513), .A2(new_n547), .B1(new_n515), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n546), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G860), .ZN(G153));
  AND3_X1   g126(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G36), .ZN(new_n553));
  XOR2_X1   g128(.A(new_n553), .B(KEYINPUT75), .Z(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G188));
  AOI22_X1  g132(.A1(new_n508), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n558));
  INV_X1    g133(.A(G91), .ZN(new_n559));
  OAI22_X1  g134(.A1(new_n558), .A2(new_n510), .B1(new_n513), .B2(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n519), .A2(new_n562), .A3(G53), .ZN(new_n563));
  INV_X1    g138(.A(G53), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n515), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n561), .A2(new_n566), .ZN(G299));
  INV_X1    g142(.A(G171), .ZN(G301));
  NAND2_X1  g143(.A1(new_n527), .A2(new_n529), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n569), .A2(new_n521), .ZN(G286));
  INV_X1    g145(.A(G166), .ZN(G303));
  NAND2_X1  g146(.A1(new_n531), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n508), .B2(G74), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n519), .A2(G49), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n508), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n510), .ZN(new_n577));
  INV_X1    g152(.A(G86), .ZN(new_n578));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n513), .A2(new_n578), .B1(new_n515), .B2(new_n579), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n577), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n531), .A2(G85), .B1(G47), .B2(new_n519), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n508), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n510), .B2(new_n583), .ZN(G290));
  INV_X1    g159(.A(G868), .ZN(new_n585));
  NOR2_X1   g160(.A1(G301), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g161(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n587));
  NAND3_X1  g162(.A1(new_n531), .A2(G92), .A3(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n587), .ZN(new_n589));
  INV_X1    g164(.A(G92), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n589), .B1(new_n513), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n519), .A2(G54), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n508), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(new_n510), .ZN(new_n595));
  NOR2_X1   g170(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT77), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n586), .B1(new_n597), .B2(new_n585), .ZN(G321));
  XNOR2_X1  g173(.A(G321), .B(KEYINPUT78), .ZN(G284));
  OR3_X1    g174(.A1(G168), .A2(KEYINPUT79), .A3(new_n585), .ZN(new_n600));
  OAI21_X1  g175(.A(KEYINPUT79), .B1(G168), .B2(new_n585), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n560), .B1(new_n565), .B2(new_n563), .ZN(new_n602));
  OAI211_X1 g177(.A(new_n600), .B(new_n601), .C1(G868), .C2(new_n602), .ZN(G297));
  OAI211_X1 g178(.A(new_n600), .B(new_n601), .C1(G868), .C2(new_n602), .ZN(G280));
  INV_X1    g179(.A(G559), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n597), .B1(new_n605), .B2(G860), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT80), .ZN(G148));
  NAND2_X1  g182(.A1(new_n597), .A2(new_n605), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n550), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n473), .A2(G2104), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  INV_X1    g189(.A(G2100), .ZN(new_n615));
  OR2_X1    g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n473), .A2(G135), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n483), .A2(G123), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n480), .A2(G111), .ZN(new_n620));
  OAI21_X1  g195(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n621));
  OAI211_X1 g196(.A(new_n618), .B(new_n619), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(KEYINPUT81), .B(G2096), .Z(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND3_X1  g199(.A1(new_n616), .A2(new_n617), .A3(new_n624), .ZN(G156));
  XNOR2_X1  g200(.A(G2443), .B(G2446), .ZN(new_n626));
  INV_X1    g201(.A(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(G2427), .B(G2438), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(G2430), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  INV_X1    g205(.A(G2430), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n633), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n634), .A3(new_n632), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n636), .A2(KEYINPUT14), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT16), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n640), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT14), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n630), .B(G2430), .ZN(new_n644));
  AOI21_X1  g219(.A(new_n643), .B1(new_n644), .B2(new_n634), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n642), .B1(new_n645), .B2(new_n636), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n627), .B1(new_n641), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n638), .A2(new_n640), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n645), .A2(new_n642), .A3(new_n636), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n626), .A3(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n647), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g230(.A1(new_n647), .A2(KEYINPUT82), .A3(new_n652), .A4(new_n649), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n647), .A2(new_n652), .ZN(new_n659));
  AOI21_X1  g234(.A(new_n658), .B1(new_n659), .B2(new_n648), .ZN(new_n660));
  AND3_X1   g235(.A1(new_n657), .A2(KEYINPUT83), .A3(new_n660), .ZN(new_n661));
  AOI21_X1  g236(.A(KEYINPUT83), .B1(new_n657), .B2(new_n660), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(G401));
  XNOR2_X1  g238(.A(G2096), .B(G2100), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(new_n665));
  XOR2_X1   g240(.A(G2084), .B(G2090), .Z(new_n666));
  XNOR2_X1  g241(.A(G2067), .B(G2678), .ZN(new_n667));
  OR2_X1    g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n666), .A2(new_n667), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(KEYINPUT17), .A3(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n671), .B1(new_n666), .B2(new_n667), .ZN(new_n673));
  XOR2_X1   g248(.A(G2072), .B(G2078), .Z(new_n674));
  NOR2_X1   g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n672), .A2(new_n675), .ZN(new_n676));
  OAI211_X1 g251(.A(new_n670), .B(new_n671), .C1(new_n674), .C2(new_n673), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(KEYINPUT84), .A3(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(KEYINPUT84), .B1(new_n676), .B2(new_n677), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n665), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n680), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n678), .A3(new_n664), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n681), .A2(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1971), .B(G1976), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT19), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1956), .B(G2474), .Z(new_n688));
  XOR2_X1   g263(.A(G1961), .B(G1966), .Z(new_n689));
  AND2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT20), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n688), .A2(new_n689), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n690), .A2(new_n694), .ZN(new_n695));
  MUX2_X1   g270(.A(new_n695), .B(new_n694), .S(new_n687), .Z(new_n696));
  NOR2_X1   g271(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  XOR2_X1   g274(.A(G1991), .B(G1996), .Z(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(G1981), .B(G1986), .ZN(new_n702));
  INV_X1    g277(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n699), .A2(new_n700), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n699), .A2(new_n700), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n702), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(G229));
  INV_X1    g284(.A(G16), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G23), .ZN(new_n711));
  INV_X1    g286(.A(G288), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT87), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT33), .B(G1976), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OR2_X1    g291(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n714), .A2(new_n716), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n710), .A2(G22), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G166), .B2(new_n710), .ZN(new_n720));
  INV_X1    g295(.A(G1971), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(G6), .A2(G16), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n577), .A2(new_n580), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(G16), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT32), .B(G1981), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n717), .A2(new_n718), .A3(new_n722), .A4(new_n727), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT86), .B(KEYINPUT34), .Z(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n473), .A2(G131), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n483), .A2(G119), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n480), .A2(G107), .ZN(new_n734));
  OAI21_X1  g309(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n732), .B(new_n733), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT85), .Z(new_n737));
  MUX2_X1   g312(.A(G25), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  MUX2_X1   g315(.A(G24), .B(G290), .S(G16), .Z(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1986), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n730), .A2(new_n731), .A3(new_n740), .A4(new_n743), .ZN(new_n744));
  NOR2_X1   g319(.A1(KEYINPUT88), .A2(KEYINPUT36), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT89), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n744), .B(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n474), .A2(G105), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n473), .A2(G141), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n483), .A2(G129), .ZN(new_n750));
  NAND3_X1  g325(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT26), .Z(new_n752));
  AND4_X1   g327(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(G29), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n754), .B2(G32), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT27), .B(G1996), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT24), .ZN(new_n759));
  INV_X1    g334(.A(G34), .ZN(new_n760));
  AOI21_X1  g335(.A(G29), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n761), .B1(new_n759), .B2(new_n760), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G160), .B2(new_n754), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n758), .B1(G2084), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n756), .B2(new_n757), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT31), .B(G11), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT93), .B(G28), .ZN(new_n767));
  INV_X1    g342(.A(KEYINPUT30), .ZN(new_n768));
  AOI21_X1  g343(.A(G29), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n768), .B2(new_n767), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n766), .B(new_n770), .C1(new_n622), .C2(new_n754), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n754), .A2(G26), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT28), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n492), .A2(G140), .A3(new_n480), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n492), .A2(G128), .A3(G2105), .ZN(new_n775));
  OR2_X1    g350(.A1(G104), .A2(G2105), .ZN(new_n776));
  OAI211_X1 g351(.A(new_n776), .B(G2104), .C1(G116), .C2(new_n480), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n774), .A2(new_n775), .A3(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n773), .B1(new_n779), .B2(new_n754), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(G2067), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n771), .B(new_n781), .C1(G2084), .C2(new_n763), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n754), .A2(G27), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G164), .B2(new_n754), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n784), .B(new_n443), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n550), .A2(new_n710), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n710), .B2(G19), .ZN(new_n787));
  INV_X1    g362(.A(G1341), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND4_X1  g364(.A1(new_n765), .A2(new_n782), .A3(new_n785), .A4(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n473), .A2(G139), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n480), .A2(G103), .A3(G2104), .ZN(new_n792));
  INV_X1    g367(.A(KEYINPUT25), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT91), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n492), .A2(G127), .ZN(new_n797));
  AND2_X1   g372(.A1(G115), .A2(G2104), .ZN(new_n798));
  OAI21_X1  g373(.A(G2105), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g374(.A1(new_n796), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g375(.A1(new_n800), .A2(new_n754), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n754), .B2(G33), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(new_n442), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n754), .A2(G35), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G162), .B2(new_n754), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT29), .Z(new_n806));
  INV_X1    g381(.A(G2090), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n803), .B1(new_n788), .B2(new_n787), .C1(new_n806), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n710), .A2(G20), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT23), .Z(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G299), .B2(G16), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(G1956), .ZN(new_n812));
  INV_X1    g387(.A(G1966), .ZN(new_n813));
  NOR2_X1   g388(.A1(G168), .A2(new_n710), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n814), .B1(new_n710), .B2(G21), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n812), .B1(new_n813), .B2(new_n815), .ZN(new_n816));
  NOR3_X1   g391(.A1(new_n790), .A2(new_n808), .A3(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n815), .A2(new_n813), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n802), .A2(new_n442), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT92), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n806), .A2(new_n807), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT95), .Z(new_n822));
  NAND4_X1  g397(.A1(new_n817), .A2(new_n818), .A3(new_n820), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g398(.A1(G5), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G171), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT94), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(G1961), .ZN(new_n827));
  NOR2_X1   g402(.A1(G4), .A2(G16), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(new_n597), .B2(G16), .ZN(new_n829));
  XNOR2_X1  g404(.A(KEYINPUT90), .B(G1348), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n827), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g407(.A1(new_n747), .A2(new_n823), .A3(new_n832), .ZN(G311));
  INV_X1    g408(.A(G311), .ZN(G150));
  AOI22_X1  g409(.A1(new_n508), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n510), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(G93), .ZN(new_n838));
  INV_X1    g413(.A(G55), .ZN(new_n839));
  OAI22_X1  g414(.A1(new_n513), .A2(new_n838), .B1(new_n515), .B2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g418(.A(KEYINPUT96), .B1(new_n836), .B2(new_n840), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(new_n550), .A3(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n837), .A2(new_n841), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n546), .A2(new_n549), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n846), .A2(new_n847), .A3(KEYINPUT96), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n849), .B(KEYINPUT38), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n597), .A2(G559), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n850), .B(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n854));
  NOR3_X1   g429(.A1(new_n853), .A2(new_n854), .A3(G860), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n846), .A2(G860), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(KEYINPUT37), .ZN(new_n857));
  OR2_X1    g432(.A1(new_n855), .A2(new_n857), .ZN(G145));
  XNOR2_X1  g433(.A(new_n476), .B(new_n622), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n485), .ZN(new_n860));
  INV_X1    g435(.A(new_n800), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n749), .A2(new_n750), .A3(new_n748), .A4(new_n752), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n496), .A2(new_n500), .A3(new_n778), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n778), .B1(new_n496), .B2(new_n500), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n501), .A2(new_n779), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n496), .A2(new_n500), .A3(new_n778), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n866), .A2(new_n753), .A3(new_n867), .ZN(new_n868));
  AND3_X1   g443(.A1(new_n865), .A2(new_n868), .A3(KEYINPUT97), .ZN(new_n869));
  AOI21_X1  g444(.A(KEYINPUT97), .B1(new_n865), .B2(new_n868), .ZN(new_n870));
  OR3_X1    g445(.A1(new_n861), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g446(.A1(new_n863), .A2(new_n864), .A3(new_n862), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n753), .B1(new_n866), .B2(new_n867), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT98), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT98), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n865), .A2(new_n868), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(KEYINPUT99), .B1(new_n877), .B2(new_n861), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n879));
  AOI211_X1 g454(.A(new_n879), .B(new_n800), .C1(new_n874), .C2(new_n876), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n871), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n483), .A2(G130), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n480), .A2(G118), .ZN(new_n883));
  OAI21_X1  g458(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n885), .B1(G142), .B2(new_n473), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(new_n613), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(new_n736), .Z(new_n888));
  AOI21_X1  g463(.A(new_n860), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  NOR3_X1   g464(.A1(new_n861), .A2(new_n869), .A3(new_n870), .ZN(new_n890));
  AND3_X1   g465(.A1(new_n865), .A2(new_n868), .A3(new_n875), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n875), .B1(new_n865), .B2(new_n868), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n861), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(new_n879), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n877), .A2(KEYINPUT99), .A3(new_n861), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n888), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g473(.A(G37), .B1(new_n889), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(KEYINPUT100), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n896), .B2(new_n897), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n881), .A2(KEYINPUT100), .A3(new_n888), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n898), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT101), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n903), .A2(new_n904), .A3(new_n860), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n904), .B1(new_n903), .B2(new_n860), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n907), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g483(.A1(new_n846), .A2(G868), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT103), .ZN(new_n910));
  OR2_X1    g485(.A1(new_n592), .A2(new_n595), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n911), .A2(G299), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n596), .A2(new_n602), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT41), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n916), .A3(new_n913), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  INV_X1    g493(.A(new_n918), .ZN(new_n919));
  AND2_X1   g494(.A1(new_n912), .A2(new_n913), .ZN(new_n920));
  XNOR2_X1  g495(.A(new_n920), .B(KEYINPUT102), .ZN(new_n921));
  XNOR2_X1  g496(.A(new_n608), .B(new_n849), .ZN(new_n922));
  MUX2_X1   g497(.A(new_n919), .B(new_n921), .S(new_n922), .Z(new_n923));
  XNOR2_X1  g498(.A(G290), .B(new_n724), .ZN(new_n924));
  XNOR2_X1  g499(.A(G166), .B(G288), .ZN(new_n925));
  XOR2_X1   g500(.A(new_n924), .B(new_n925), .Z(new_n926));
  XOR2_X1   g501(.A(new_n926), .B(KEYINPUT42), .Z(new_n927));
  AOI21_X1  g502(.A(new_n910), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n923), .B2(new_n927), .ZN(new_n929));
  OR3_X1    g504(.A1(new_n923), .A2(KEYINPUT103), .A3(new_n927), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n909), .B1(new_n931), .B2(G868), .ZN(G295));
  AOI21_X1  g507(.A(new_n909), .B1(new_n931), .B2(G868), .ZN(G331));
  NAND3_X1  g508(.A1(G286), .A2(new_n537), .A3(new_n543), .ZN(new_n934));
  NAND2_X1  g509(.A1(G171), .A2(G168), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n849), .ZN(new_n937));
  NAND4_X1  g512(.A1(new_n934), .A2(new_n935), .A3(new_n848), .A4(new_n845), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n937), .A2(new_n938), .A3(KEYINPUT105), .ZN(new_n939));
  OR3_X1    g514(.A1(new_n936), .A2(new_n849), .A3(KEYINPUT105), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(new_n920), .ZN(new_n942));
  INV_X1    g517(.A(new_n926), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n937), .A2(new_n938), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(new_n918), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n942), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G37), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n914), .B1(new_n939), .B2(new_n940), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n944), .A2(new_n918), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n926), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n946), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n917), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n912), .A2(KEYINPUT106), .A3(new_n916), .A4(new_n913), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(new_n915), .A3(new_n954), .ZN(new_n955));
  OAI22_X1  g530(.A1(new_n941), .A2(new_n955), .B1(new_n921), .B2(new_n944), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n926), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n957), .A2(new_n947), .A3(new_n946), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n959));
  OAI221_X1 g534(.A(KEYINPUT44), .B1(KEYINPUT43), .B2(new_n951), .C1(new_n959), .C2(KEYINPUT107), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(KEYINPUT107), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT43), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n957), .A2(new_n946), .A3(new_n963), .A4(new_n947), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n966));
  OAI22_X1  g541(.A1(new_n960), .A2(new_n961), .B1(new_n965), .B2(new_n966), .ZN(G397));
  AOI21_X1  g542(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n969));
  AND3_X1   g544(.A1(new_n472), .A2(G40), .A3(new_n475), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(G2067), .ZN(new_n972));
  XNOR2_X1  g547(.A(new_n778), .B(new_n972), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT109), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n971), .A2(new_n976), .A3(new_n753), .ZN(new_n977));
  NOR2_X1   g552(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n971), .A2(G1996), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n753), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT108), .ZN(new_n981));
  INV_X1    g556(.A(new_n971), .ZN(new_n982));
  INV_X1    g557(.A(new_n739), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n736), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n978), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  XNOR2_X1  g561(.A(G290), .B(G1986), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n986), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n990));
  INV_X1    g565(.A(G8), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n990), .B1(G166), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n968), .A2(KEYINPUT45), .ZN(new_n994));
  AND2_X1   g569(.A1(new_n994), .A2(new_n970), .ZN(new_n995));
  INV_X1    g570(.A(G1384), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n501), .A2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT110), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n969), .A2(KEYINPUT110), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n995), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT50), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n970), .B1(new_n968), .B2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n997), .A2(KEYINPUT50), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  XOR2_X1   g582(.A(KEYINPUT111), .B(G2090), .Z(new_n1008));
  AOI22_X1  g583(.A1(new_n1003), .A2(new_n721), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT115), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  XNOR2_X1  g586(.A(KEYINPUT113), .B(G8), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1012), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1013), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n993), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n993), .B(KEYINPUT112), .ZN(new_n1016));
  NOR2_X1   g591(.A1(new_n1009), .A2(new_n991), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n712), .A2(G1976), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1012), .B1(new_n970), .B2(new_n968), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  INV_X1    g597(.A(G1976), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT52), .B1(G288), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1019), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1020), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1028), .B1(G305), .B2(G1981), .ZN(new_n1029));
  INV_X1    g604(.A(G1981), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n724), .A2(KEYINPUT114), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NOR2_X1   g607(.A1(new_n724), .A2(new_n1030), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1032), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT49), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1027), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1033), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(KEYINPUT49), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1026), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1015), .A2(new_n1018), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(KEYINPUT124), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT124), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1015), .A2(new_n1043), .A3(new_n1018), .A4(new_n1040), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  AOI21_X1  g620(.A(KEYINPUT57), .B1(new_n561), .B2(KEYINPUT117), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G299), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n561), .B(new_n566), .C1(KEYINPUT117), .C2(KEYINPUT57), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT56), .B(G2072), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n995), .A2(new_n1001), .A3(new_n1002), .A4(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(G1956), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1052), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1049), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(G1348), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1055), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n970), .A2(new_n972), .A3(new_n968), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n597), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1051), .A2(new_n1049), .A3(new_n1053), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1054), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n995), .A2(new_n1001), .A3(new_n976), .A4(new_n1002), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT118), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n970), .A2(new_n968), .ZN(new_n1065));
  XOR2_X1   g640(.A(KEYINPUT58), .B(G1341), .Z(new_n1066));
  AOI22_X1  g641(.A1(new_n1063), .A2(new_n1064), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AND3_X1   g642(.A1(new_n995), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1068), .A2(KEYINPUT118), .A3(new_n976), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n847), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g645(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  XNOR2_X1  g647(.A(new_n1070), .B(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1054), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1074), .A2(KEYINPUT61), .A3(new_n1061), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT60), .ZN(new_n1076));
  AOI21_X1  g651(.A(new_n1076), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1059), .B1(new_n597), .B2(new_n1077), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT61), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1061), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(new_n1054), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1059), .B(new_n1079), .C1(new_n597), .C2(new_n1077), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1075), .A2(new_n1081), .A3(new_n1084), .A4(new_n1085), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1062), .B1(new_n1073), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(G2084), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n999), .A2(new_n970), .A3(new_n994), .ZN(new_n1089));
  AOI22_X1  g664(.A1(new_n1007), .A2(new_n1088), .B1(new_n1089), .B2(new_n813), .ZN(new_n1090));
  NOR2_X1   g665(.A1(G168), .A2(new_n1012), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1090), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT121), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n1090), .B2(new_n991), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1096), .A2(new_n1098), .A3(new_n1092), .ZN(new_n1099));
  AND2_X1   g674(.A1(new_n1099), .A2(KEYINPUT51), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n1090), .A2(new_n1012), .ZN(new_n1101));
  NOR3_X1   g676(.A1(new_n1101), .A2(KEYINPUT51), .A3(new_n1091), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1094), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n1068), .B2(new_n443), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1007), .A2(G1961), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AND2_X1   g681(.A1(new_n999), .A2(new_n994), .ZN(new_n1107));
  OR2_X1    g682(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1108));
  NAND2_X1  g683(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n472), .A2(KEYINPUT53), .A3(G40), .A4(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1111), .B1(KEYINPUT122), .B2(new_n475), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1107), .B(new_n1112), .C1(KEYINPUT122), .C2(new_n475), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  XNOR2_X1  g689(.A(G171), .B(KEYINPUT54), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1107), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n970), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1106), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1118), .B2(new_n1115), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1087), .A2(new_n1103), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT62), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1121), .B(new_n1094), .C1(new_n1100), .C2(new_n1102), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1102), .B1(new_n1099), .B2(KEYINPUT51), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT62), .B1(new_n1123), .B2(new_n1093), .ZN(new_n1124));
  AOI21_X1  g699(.A(G301), .B1(new_n1106), .B2(new_n1117), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1124), .A3(new_n1125), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1045), .B1(new_n1120), .B2(new_n1126), .ZN(new_n1127));
  NOR2_X1   g702(.A1(G288), .A2(G1976), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1039), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n1020), .B1(new_n1038), .B2(KEYINPUT49), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1128), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1027), .B1(new_n1131), .B2(new_n1032), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n993), .B1(new_n1009), .B2(new_n991), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1040), .A2(G168), .A3(new_n1101), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(KEYINPUT63), .ZN(new_n1135));
  NOR4_X1   g710(.A1(new_n1090), .A2(KEYINPUT63), .A3(G286), .A4(new_n1012), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1015), .A2(new_n1136), .B1(new_n1017), .B2(new_n1016), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1040), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1135), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1139), .A2(KEYINPUT116), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT116), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1135), .B(new_n1141), .C1(new_n1137), .C2(new_n1138), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n988), .B1(new_n1127), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n971), .B1(new_n753), .B2(new_n973), .ZN(new_n1145));
  OR3_X1    g720(.A1(new_n971), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT46), .B1(new_n971), .B2(G1996), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g723(.A(new_n1148), .B(KEYINPUT47), .ZN(new_n1149));
  NOR2_X1   g724(.A1(new_n737), .A2(new_n983), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n978), .A2(new_n981), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n779), .A2(new_n972), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n971), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n986), .ZN(new_n1154));
  NOR3_X1   g729(.A1(new_n971), .A2(G1986), .A3(G290), .ZN(new_n1155));
  XOR2_X1   g730(.A(new_n1155), .B(KEYINPUT48), .Z(new_n1156));
  AOI211_X1 g731(.A(new_n1149), .B(new_n1153), .C1(new_n1154), .C2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1144), .A2(new_n1157), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n1160));
  NAND3_X1  g734(.A1(new_n681), .A2(new_n683), .A3(G319), .ZN(new_n1161));
  INV_X1    g735(.A(KEYINPUT125), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g737(.A1(new_n681), .A2(new_n683), .A3(KEYINPUT125), .A4(G319), .ZN(new_n1164));
  NAND2_X1  g738(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g739(.A(new_n1165), .B1(new_n661), .B2(new_n662), .ZN(new_n1166));
  INV_X1    g740(.A(KEYINPUT126), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g742(.A(new_n1165), .B(KEYINPUT126), .C1(new_n661), .C2(new_n662), .ZN(new_n1169));
  NAND3_X1  g743(.A1(new_n1168), .A2(new_n708), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n1170), .B1(new_n962), .B2(new_n964), .ZN(new_n1171));
  AND3_X1   g745(.A1(new_n907), .A2(new_n1160), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g746(.A(new_n1160), .B1(new_n907), .B2(new_n1171), .ZN(new_n1173));
  NOR2_X1   g747(.A1(new_n1172), .A2(new_n1173), .ZN(G308));
  NAND2_X1  g748(.A1(new_n907), .A2(new_n1171), .ZN(G225));
endmodule


