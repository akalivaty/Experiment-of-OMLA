

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577;

  XNOR2_X1 U321 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n388) );
  XNOR2_X1 U322 ( .A(n389), .B(n388), .ZN(n519) );
  XNOR2_X1 U323 ( .A(n340), .B(KEYINPUT73), .ZN(n341) );
  XNOR2_X1 U324 ( .A(n342), .B(n341), .ZN(n343) );
  NOR2_X1 U325 ( .A1(n522), .A2(n447), .ZN(n554) );
  XNOR2_X1 U326 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U327 ( .A(n451), .B(n450), .ZN(G1349GAT) );
  XOR2_X1 U328 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n290) );
  XNOR2_X1 U329 ( .A(G169GAT), .B(G15GAT), .ZN(n289) );
  XNOR2_X1 U330 ( .A(n290), .B(n289), .ZN(n302) );
  XOR2_X1 U331 ( .A(G120GAT), .B(G71GAT), .Z(n339) );
  XOR2_X1 U332 ( .A(G176GAT), .B(G190GAT), .Z(n292) );
  XNOR2_X1 U333 ( .A(G43GAT), .B(G99GAT), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U335 ( .A(n339), .B(n293), .Z(n295) );
  NAND2_X1 U336 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U337 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U338 ( .A(n296), .B(KEYINPUT85), .Z(n300) );
  XOR2_X1 U339 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n298) );
  XNOR2_X1 U340 ( .A(G183GAT), .B(KEYINPUT18), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n397) );
  XNOR2_X1 U342 ( .A(n397), .B(KEYINPUT86), .ZN(n299) );
  XNOR2_X1 U343 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n307) );
  XOR2_X1 U345 ( .A(KEYINPUT82), .B(G127GAT), .Z(n304) );
  XNOR2_X1 U346 ( .A(KEYINPUT0), .B(KEYINPUT83), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n306) );
  XOR2_X1 U348 ( .A(G113GAT), .B(G134GAT), .Z(n305) );
  XOR2_X1 U349 ( .A(n306), .B(n305), .Z(n409) );
  XOR2_X1 U350 ( .A(n307), .B(n409), .Z(n457) );
  INV_X1 U351 ( .A(n457), .ZN(n513) );
  INV_X1 U352 ( .A(n513), .ZN(n522) );
  XOR2_X1 U353 ( .A(KEYINPUT65), .B(KEYINPUT75), .Z(n309) );
  XNOR2_X1 U354 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n327) );
  XOR2_X1 U356 ( .A(KEYINPUT11), .B(KEYINPUT9), .Z(n311) );
  XNOR2_X1 U357 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n310) );
  XNOR2_X1 U358 ( .A(n311), .B(n310), .ZN(n315) );
  XOR2_X1 U359 ( .A(KEYINPUT10), .B(G92GAT), .Z(n313) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G162GAT), .ZN(n312) );
  XNOR2_X1 U361 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U362 ( .A(n315), .B(n314), .Z(n325) );
  XNOR2_X1 U363 ( .A(G43GAT), .B(KEYINPUT7), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n316), .B(G29GAT), .ZN(n317) );
  XOR2_X1 U365 ( .A(n317), .B(KEYINPUT67), .Z(n319) );
  XNOR2_X1 U366 ( .A(G50GAT), .B(KEYINPUT8), .ZN(n318) );
  XNOR2_X1 U367 ( .A(n319), .B(n318), .ZN(n356) );
  XOR2_X1 U368 ( .A(G190GAT), .B(G218GAT), .Z(n392) );
  XNOR2_X1 U369 ( .A(G99GAT), .B(G85GAT), .ZN(n320) );
  XOR2_X1 U370 ( .A(n320), .B(KEYINPUT74), .Z(n330) );
  XNOR2_X1 U371 ( .A(n392), .B(n330), .ZN(n322) );
  NAND2_X1 U372 ( .A1(G232GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U373 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U374 ( .A(n356), .B(n323), .ZN(n324) );
  XNOR2_X1 U375 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U376 ( .A(n327), .B(n326), .Z(n553) );
  XNOR2_X1 U377 ( .A(KEYINPUT110), .B(KEYINPUT46), .ZN(n358) );
  XOR2_X1 U378 ( .A(KEYINPUT13), .B(KEYINPUT71), .Z(n329) );
  XNOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT70), .ZN(n328) );
  XNOR2_X1 U380 ( .A(n329), .B(n328), .ZN(n375) );
  XNOR2_X1 U381 ( .A(n375), .B(n330), .ZN(n344) );
  XOR2_X1 U382 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n332) );
  NAND2_X1 U383 ( .A1(G230GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n332), .B(n331), .ZN(n333) );
  XOR2_X1 U385 ( .A(n333), .B(KEYINPUT72), .Z(n338) );
  XOR2_X1 U386 ( .A(G64GAT), .B(G204GAT), .Z(n335) );
  XNOR2_X1 U387 ( .A(G176GAT), .B(G92GAT), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n395) );
  XNOR2_X1 U389 ( .A(G148GAT), .B(G106GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(G78GAT), .ZN(n441) );
  XNOR2_X1 U391 ( .A(n395), .B(n441), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U393 ( .A(n339), .B(KEYINPUT32), .Z(n340) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n564) );
  XNOR2_X1 U395 ( .A(KEYINPUT41), .B(n564), .ZN(n540) );
  XOR2_X1 U396 ( .A(KEYINPUT66), .B(KEYINPUT29), .Z(n346) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U399 ( .A(n347), .B(KEYINPUT30), .Z(n351) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G36GAT), .ZN(n348) );
  XNOR2_X1 U401 ( .A(n348), .B(G8GAT), .ZN(n398) );
  XNOR2_X1 U402 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n349) );
  XNOR2_X1 U403 ( .A(n349), .B(G15GAT), .ZN(n371) );
  XNOR2_X1 U404 ( .A(n398), .B(n371), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U406 ( .A(G141GAT), .B(G22GAT), .Z(n433) );
  XOR2_X1 U407 ( .A(n352), .B(n433), .Z(n354) );
  XNOR2_X1 U408 ( .A(G197GAT), .B(G113GAT), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n496) );
  INV_X1 U411 ( .A(n496), .ZN(n559) );
  NAND2_X1 U412 ( .A1(n540), .A2(n559), .ZN(n357) );
  XOR2_X1 U413 ( .A(n358), .B(n357), .Z(n359) );
  NOR2_X1 U414 ( .A1(n553), .A2(n359), .ZN(n380) );
  XOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n361) );
  XNOR2_X1 U416 ( .A(KEYINPUT81), .B(KEYINPUT12), .ZN(n360) );
  XNOR2_X1 U417 ( .A(n361), .B(n360), .ZN(n379) );
  XOR2_X1 U418 ( .A(KEYINPUT79), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U419 ( .A(G8GAT), .B(G22GAT), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n367) );
  XOR2_X1 U421 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n365) );
  XNOR2_X1 U422 ( .A(G127GAT), .B(G155GAT), .ZN(n364) );
  XNOR2_X1 U423 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U424 ( .A(n367), .B(n366), .Z(n373) );
  XOR2_X1 U425 ( .A(G64GAT), .B(G71GAT), .Z(n369) );
  NAND2_X1 U426 ( .A1(G231GAT), .A2(G233GAT), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U428 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U429 ( .A(n373), .B(n372), .ZN(n374) );
  XOR2_X1 U430 ( .A(n374), .B(G211GAT), .Z(n377) );
  XNOR2_X1 U431 ( .A(G183GAT), .B(n375), .ZN(n376) );
  XNOR2_X1 U432 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U433 ( .A(n379), .B(n378), .Z(n569) );
  INV_X1 U434 ( .A(n569), .ZN(n482) );
  NAND2_X1 U435 ( .A1(n380), .A2(n482), .ZN(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT47), .B(n381), .ZN(n387) );
  XOR2_X1 U437 ( .A(KEYINPUT36), .B(n553), .Z(n574) );
  NOR2_X1 U438 ( .A1(n574), .A2(n482), .ZN(n383) );
  XNOR2_X1 U439 ( .A(KEYINPUT45), .B(KEYINPUT111), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n385) );
  XOR2_X1 U441 ( .A(KEYINPUT69), .B(n496), .Z(n452) );
  NAND2_X1 U442 ( .A1(n452), .A2(n564), .ZN(n384) );
  NOR2_X1 U443 ( .A1(n385), .A2(n384), .ZN(n386) );
  NOR2_X1 U444 ( .A1(n387), .A2(n386), .ZN(n389) );
  XOR2_X1 U445 ( .A(KEYINPUT21), .B(KEYINPUT88), .Z(n391) );
  XNOR2_X1 U446 ( .A(G197GAT), .B(G211GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n440) );
  XOR2_X1 U448 ( .A(n440), .B(n392), .Z(n394) );
  NAND2_X1 U449 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n396) );
  XOR2_X1 U451 ( .A(n396), .B(n395), .Z(n400) );
  XNOR2_X1 U452 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U453 ( .A(n400), .B(n399), .ZN(n511) );
  XNOR2_X1 U454 ( .A(n511), .B(KEYINPUT119), .ZN(n401) );
  NOR2_X1 U455 ( .A1(n519), .A2(n401), .ZN(n402) );
  XNOR2_X1 U456 ( .A(n402), .B(KEYINPUT54), .ZN(n428) );
  XOR2_X1 U457 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n404) );
  XNOR2_X1 U458 ( .A(KEYINPUT4), .B(KEYINPUT96), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U460 ( .A(G148GAT), .B(G57GAT), .Z(n406) );
  XNOR2_X1 U461 ( .A(G1GAT), .B(G120GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U463 ( .A(n408), .B(n407), .Z(n415) );
  INV_X1 U464 ( .A(n409), .ZN(n413) );
  XOR2_X1 U465 ( .A(KEYINPUT92), .B(KEYINPUT94), .Z(n411) );
  XNOR2_X1 U466 ( .A(G141GAT), .B(KEYINPUT93), .ZN(n410) );
  XNOR2_X1 U467 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U468 ( .A(n413), .B(n412), .Z(n414) );
  XNOR2_X1 U469 ( .A(n415), .B(n414), .ZN(n426) );
  XOR2_X1 U470 ( .A(KEYINPUT95), .B(KEYINPUT1), .Z(n417) );
  NAND2_X1 U471 ( .A1(G225GAT), .A2(G233GAT), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U473 ( .A(n418), .B(G85GAT), .Z(n424) );
  XNOR2_X1 U474 ( .A(KEYINPUT89), .B(KEYINPUT3), .ZN(n419) );
  XNOR2_X1 U475 ( .A(n419), .B(KEYINPUT90), .ZN(n420) );
  XOR2_X1 U476 ( .A(n420), .B(G155GAT), .Z(n422) );
  XNOR2_X1 U477 ( .A(KEYINPUT2), .B(G162GAT), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n422), .B(n421), .ZN(n445) );
  XNOR2_X1 U479 ( .A(G29GAT), .B(n445), .ZN(n423) );
  XNOR2_X1 U480 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U481 ( .A(n426), .B(n425), .ZN(n509) );
  INV_X1 U482 ( .A(n509), .ZN(n427) );
  NAND2_X1 U483 ( .A1(n428), .A2(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n429), .B(KEYINPUT64), .ZN(n558) );
  XOR2_X1 U485 ( .A(KEYINPUT23), .B(G218GAT), .Z(n431) );
  XNOR2_X1 U486 ( .A(G50GAT), .B(G204GAT), .ZN(n430) );
  XNOR2_X1 U487 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U488 ( .A(n433), .B(n432), .Z(n435) );
  NAND2_X1 U489 ( .A1(G228GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n435), .B(n434), .ZN(n439) );
  XOR2_X1 U491 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n437) );
  XNOR2_X1 U492 ( .A(KEYINPUT91), .B(KEYINPUT24), .ZN(n436) );
  XNOR2_X1 U493 ( .A(n437), .B(n436), .ZN(n438) );
  XOR2_X1 U494 ( .A(n439), .B(n438), .Z(n443) );
  XNOR2_X1 U495 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U496 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n458) );
  NOR2_X1 U498 ( .A1(n558), .A2(n458), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n446), .B(KEYINPUT55), .ZN(n447) );
  XNOR2_X1 U500 ( .A(n540), .B(KEYINPUT106), .ZN(n527) );
  NAND2_X1 U501 ( .A1(n554), .A2(n527), .ZN(n451) );
  XOR2_X1 U502 ( .A(G176GAT), .B(KEYINPUT56), .Z(n449) );
  XNOR2_X1 U503 ( .A(KEYINPUT120), .B(KEYINPUT57), .ZN(n448) );
  INV_X1 U504 ( .A(n452), .ZN(n549) );
  NAND2_X1 U505 ( .A1(n549), .A2(n564), .ZN(n485) );
  XNOR2_X1 U506 ( .A(KEYINPUT28), .B(n458), .ZN(n525) );
  XNOR2_X1 U507 ( .A(n511), .B(KEYINPUT27), .ZN(n461) );
  NAND2_X1 U508 ( .A1(n509), .A2(n461), .ZN(n520) );
  NOR2_X1 U509 ( .A1(n525), .A2(n520), .ZN(n453) );
  NAND2_X1 U510 ( .A1(n453), .A2(n457), .ZN(n454) );
  XNOR2_X1 U511 ( .A(n454), .B(KEYINPUT97), .ZN(n467) );
  AND2_X1 U512 ( .A1(n513), .A2(n511), .ZN(n455) );
  NOR2_X1 U513 ( .A1(n458), .A2(n455), .ZN(n456) );
  XNOR2_X1 U514 ( .A(n456), .B(KEYINPUT25), .ZN(n463) );
  NAND2_X1 U515 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT98), .ZN(n460) );
  XOR2_X1 U517 ( .A(KEYINPUT26), .B(n460), .Z(n537) );
  NAND2_X1 U518 ( .A1(n537), .A2(n461), .ZN(n462) );
  NAND2_X1 U519 ( .A1(n463), .A2(n462), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT99), .B(n464), .ZN(n465) );
  NOR2_X1 U521 ( .A1(n509), .A2(n465), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n480) );
  NOR2_X1 U523 ( .A1(n553), .A2(n482), .ZN(n468) );
  XOR2_X1 U524 ( .A(KEYINPUT16), .B(n468), .Z(n469) );
  OR2_X1 U525 ( .A1(n480), .A2(n469), .ZN(n497) );
  NOR2_X1 U526 ( .A1(n485), .A2(n497), .ZN(n477) );
  NAND2_X1 U527 ( .A1(n477), .A2(n509), .ZN(n470) );
  XNOR2_X1 U528 ( .A(KEYINPUT34), .B(n470), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G1GAT), .B(n471), .ZN(G1324GAT) );
  NAND2_X1 U530 ( .A1(n477), .A2(n511), .ZN(n472) );
  XNOR2_X1 U531 ( .A(n472), .B(KEYINPUT100), .ZN(n473) );
  XNOR2_X1 U532 ( .A(G8GAT), .B(n473), .ZN(G1325GAT) );
  XOR2_X1 U533 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n475) );
  NAND2_X1 U534 ( .A1(n477), .A2(n513), .ZN(n474) );
  XNOR2_X1 U535 ( .A(n475), .B(n474), .ZN(n476) );
  XOR2_X1 U536 ( .A(G15GAT), .B(n476), .Z(G1326GAT) );
  NAND2_X1 U537 ( .A1(n477), .A2(n525), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT102), .ZN(n479) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n479), .ZN(G1327GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT104), .B(KEYINPUT39), .Z(n488) );
  NOR2_X1 U541 ( .A1(n574), .A2(n480), .ZN(n481) );
  NAND2_X1 U542 ( .A1(n482), .A2(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n483), .B(KEYINPUT103), .ZN(n484) );
  XNOR2_X1 U544 ( .A(KEYINPUT37), .B(n484), .ZN(n508) );
  NOR2_X1 U545 ( .A1(n485), .A2(n508), .ZN(n486) );
  XNOR2_X1 U546 ( .A(n486), .B(KEYINPUT38), .ZN(n494) );
  NAND2_X1 U547 ( .A1(n494), .A2(n509), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(n489), .ZN(G1328GAT) );
  NAND2_X1 U550 ( .A1(n494), .A2(n511), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(G36GAT), .ZN(G1329GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n492) );
  NAND2_X1 U553 ( .A1(n513), .A2(n494), .ZN(n491) );
  XNOR2_X1 U554 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  NAND2_X1 U556 ( .A1(n494), .A2(n525), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n495), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U558 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  NAND2_X1 U559 ( .A1(n496), .A2(n527), .ZN(n507) );
  OR2_X1 U560 ( .A1(n497), .A2(n507), .ZN(n498) );
  XNOR2_X1 U561 ( .A(n498), .B(KEYINPUT107), .ZN(n503) );
  NAND2_X1 U562 ( .A1(n503), .A2(n509), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n500), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n511), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U566 ( .A1(n503), .A2(n513), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n502), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U569 ( .A1(n503), .A2(n525), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G78GAT), .B(n506), .ZN(G1335GAT) );
  NOR2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n515) );
  NAND2_X1 U573 ( .A1(n515), .A2(n509), .ZN(n510) );
  XNOR2_X1 U574 ( .A(G85GAT), .B(n510), .ZN(G1336GAT) );
  NAND2_X1 U575 ( .A1(n515), .A2(n511), .ZN(n512) );
  XNOR2_X1 U576 ( .A(n512), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n513), .ZN(n514) );
  XNOR2_X1 U578 ( .A(n514), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT44), .B(KEYINPUT109), .Z(n517) );
  NAND2_X1 U580 ( .A1(n515), .A2(n525), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U582 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U584 ( .A(n521), .B(KEYINPUT113), .ZN(n538) );
  NOR2_X1 U585 ( .A1(n522), .A2(n538), .ZN(n523) );
  XOR2_X1 U586 ( .A(KEYINPUT114), .B(n523), .Z(n524) );
  NOR2_X1 U587 ( .A1(n525), .A2(n524), .ZN(n532) );
  NAND2_X1 U588 ( .A1(n532), .A2(n549), .ZN(n526) );
  XNOR2_X1 U589 ( .A(n526), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U590 ( .A(G120GAT), .B(KEYINPUT49), .Z(n529) );
  NAND2_X1 U591 ( .A1(n532), .A2(n527), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(G1341GAT) );
  NAND2_X1 U593 ( .A1(n532), .A2(n569), .ZN(n530) );
  XNOR2_X1 U594 ( .A(n530), .B(KEYINPUT50), .ZN(n531) );
  XNOR2_X1 U595 ( .A(G127GAT), .B(n531), .ZN(G1342GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U597 ( .A1(n532), .A2(n553), .ZN(n533) );
  XNOR2_X1 U598 ( .A(n534), .B(n533), .ZN(n536) );
  XOR2_X1 U599 ( .A(G134GAT), .B(KEYINPUT115), .Z(n535) );
  XNOR2_X1 U600 ( .A(n536), .B(n535), .ZN(G1343GAT) );
  INV_X1 U601 ( .A(n537), .ZN(n557) );
  NOR2_X1 U602 ( .A1(n538), .A2(n557), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n559), .A2(n546), .ZN(n539) );
  XNOR2_X1 U604 ( .A(G141GAT), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT117), .B(KEYINPUT53), .Z(n542) );
  NAND2_X1 U606 ( .A1(n546), .A2(n540), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n544) );
  XOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT52), .Z(n543) );
  XNOR2_X1 U609 ( .A(n544), .B(n543), .ZN(G1345GAT) );
  NAND2_X1 U610 ( .A1(n546), .A2(n569), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U612 ( .A1(n546), .A2(n553), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n547), .B(KEYINPUT118), .ZN(n548) );
  XNOR2_X1 U614 ( .A(G162GAT), .B(n548), .ZN(G1347GAT) );
  NAND2_X1 U615 ( .A1(n554), .A2(n549), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U617 ( .A(G183GAT), .B(KEYINPUT121), .Z(n552) );
  NAND2_X1 U618 ( .A1(n554), .A2(n569), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(G1350GAT) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT58), .ZN(n556) );
  XNOR2_X1 U622 ( .A(G190GAT), .B(n556), .ZN(G1351GAT) );
  XNOR2_X1 U623 ( .A(KEYINPUT60), .B(KEYINPUT122), .ZN(n563) );
  XOR2_X1 U624 ( .A(G197GAT), .B(KEYINPUT59), .Z(n561) );
  NOR2_X1 U625 ( .A1(n558), .A2(n557), .ZN(n570) );
  NAND2_X1 U626 ( .A1(n570), .A2(n559), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U628 ( .A(n563), .B(n562), .ZN(G1352GAT) );
  INV_X1 U629 ( .A(n570), .ZN(n573) );
  NOR2_X1 U630 ( .A1(n573), .A2(n564), .ZN(n568) );
  XOR2_X1 U631 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n566) );
  XNOR2_X1 U632 ( .A(G204GAT), .B(KEYINPUT124), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(G1353GAT) );
  XOR2_X1 U635 ( .A(G211GAT), .B(KEYINPUT125), .Z(n572) );
  NAND2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1354GAT) );
  NOR2_X1 U638 ( .A1(n574), .A2(n573), .ZN(n576) );
  XNOR2_X1 U639 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(G218GAT), .B(n577), .Z(G1355GAT) );
endmodule

