

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768;

  XNOR2_X1 U382 ( .A(n481), .B(KEYINPUT10), .ZN(n753) );
  INV_X1 U383 ( .A(n632), .ZN(n359) );
  INV_X1 U384 ( .A(G953), .ZN(n762) );
  NOR2_X2 U385 ( .A1(n592), .A2(n591), .ZN(n614) );
  XNOR2_X2 U386 ( .A(n456), .B(n365), .ZN(n383) );
  XNOR2_X2 U387 ( .A(n479), .B(n432), .ZN(n505) );
  XNOR2_X2 U388 ( .A(n431), .B(G128), .ZN(n479) );
  INV_X1 U389 ( .A(n730), .ZN(n629) );
  NOR2_X1 U390 ( .A1(n360), .A2(n369), .ZN(n387) );
  XNOR2_X1 U391 ( .A(n587), .B(KEYINPUT45), .ZN(n632) );
  AND2_X1 U392 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U393 ( .A(n558), .B(n557), .ZN(n766) );
  NOR2_X1 U394 ( .A1(n556), .A2(n612), .ZN(n558) );
  INV_X1 U395 ( .A(n580), .ZN(n360) );
  XNOR2_X1 U396 ( .A(n492), .B(n491), .ZN(n547) );
  OR2_X1 U397 ( .A1(n655), .A2(G902), .ZN(n561) );
  XNOR2_X1 U398 ( .A(n505), .B(n433), .ZN(n755) );
  XNOR2_X1 U399 ( .A(n482), .B(G137), .ZN(n433) );
  XNOR2_X1 U400 ( .A(G146), .B(G125), .ZN(n481) );
  XNOR2_X1 U401 ( .A(KEYINPUT68), .B(KEYINPUT4), .ZN(n482) );
  XNOR2_X1 U402 ( .A(G113), .B(G104), .ZN(n515) );
  INV_X1 U403 ( .A(G134), .ZN(n432) );
  NOR2_X1 U404 ( .A1(n398), .A2(n584), .ZN(n585) );
  XNOR2_X1 U405 ( .A(n598), .B(n436), .ZN(n551) );
  NAND2_X1 U406 ( .A1(n418), .A2(n417), .ZN(n420) );
  NAND2_X1 U407 ( .A1(KEYINPUT44), .A2(KEYINPUT65), .ZN(n417) );
  AND2_X1 U408 ( .A1(n625), .A2(n692), .ZN(n380) );
  XNOR2_X1 U409 ( .A(n606), .B(n371), .ZN(n379) );
  XNOR2_X1 U410 ( .A(n394), .B(G131), .ZN(n514) );
  INV_X1 U411 ( .A(G140), .ZN(n394) );
  INV_X1 U412 ( .A(G143), .ZN(n431) );
  NOR2_X1 U413 ( .A1(n543), .A2(n542), .ZN(n595) );
  INV_X1 U414 ( .A(n547), .ZN(n412) );
  AND2_X1 U415 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U416 ( .A(n561), .B(n560), .ZN(n594) );
  XNOR2_X1 U417 ( .A(G472), .B(KEYINPUT106), .ZN(n560) );
  XNOR2_X1 U418 ( .A(n384), .B(n364), .ZN(n598) );
  OR2_X1 U419 ( .A1(n664), .A2(G902), .ZN(n384) );
  NAND2_X1 U420 ( .A1(n406), .A2(n404), .ZN(n403) );
  NAND2_X1 U421 ( .A1(n487), .A2(KEYINPUT64), .ZN(n406) );
  NAND2_X1 U422 ( .A1(n631), .A2(n405), .ZN(n404) );
  NAND2_X1 U423 ( .A1(KEYINPUT2), .A2(KEYINPUT64), .ZN(n405) );
  XNOR2_X1 U424 ( .A(n514), .B(n393), .ZN(n754) );
  INV_X1 U425 ( .A(KEYINPUT92), .ZN(n393) );
  XNOR2_X1 U426 ( .A(n755), .B(n434), .ZN(n465) );
  NAND2_X1 U427 ( .A1(n361), .A2(n359), .ZN(n410) );
  NAND2_X1 U428 ( .A1(n389), .A2(n386), .ZN(n694) );
  AND2_X1 U429 ( .A1(n391), .A2(n390), .ZN(n389) );
  NAND2_X1 U430 ( .A1(n388), .A2(n387), .ZN(n386) );
  NAND2_X1 U431 ( .A1(n392), .A2(n369), .ZN(n391) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n626) );
  INV_X1 U433 ( .A(KEYINPUT39), .ZN(n375) );
  AND2_X1 U434 ( .A1(n614), .A2(n696), .ZN(n376) );
  NOR2_X1 U435 ( .A1(n694), .A2(n567), .ZN(n554) );
  AND2_X1 U436 ( .A1(n762), .A2(G952), .ZN(n540) );
  XNOR2_X1 U437 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n478) );
  NAND2_X1 U438 ( .A1(n360), .A2(n369), .ZN(n390) );
  OR2_X1 U439 ( .A1(n640), .A2(n631), .ZN(n492) );
  XNOR2_X1 U440 ( .A(G113), .B(G131), .ZN(n457) );
  XNOR2_X1 U441 ( .A(G101), .B(G116), .ZN(n460) );
  NAND2_X1 U442 ( .A1(n377), .A2(n628), .ZN(n730) );
  XNOR2_X1 U443 ( .A(n378), .B(n370), .ZN(n377) );
  XNOR2_X1 U444 ( .A(KEYINPUT9), .B(KEYINPUT102), .ZN(n504) );
  XNOR2_X1 U445 ( .A(G122), .B(G116), .ZN(n470) );
  NAND2_X1 U446 ( .A1(n413), .A2(n411), .ZN(n608) );
  AND2_X1 U447 ( .A1(n416), .A2(n414), .ZN(n413) );
  NAND2_X1 U448 ( .A1(n412), .A2(n366), .ZN(n411) );
  OR2_X1 U449 ( .A1(n415), .A2(n695), .ZN(n414) );
  XNOR2_X1 U450 ( .A(n599), .B(KEYINPUT110), .ZN(n609) );
  AND2_X1 U451 ( .A1(n707), .A2(n422), .ZN(n421) );
  INV_X1 U452 ( .A(n594), .ZN(n422) );
  NOR2_X1 U453 ( .A1(n706), .A2(n598), .ZN(n382) );
  XNOR2_X1 U454 ( .A(n535), .B(n534), .ZN(n559) );
  NAND2_X1 U455 ( .A1(n368), .A2(n400), .ZN(n408) );
  NAND2_X1 U456 ( .A1(n401), .A2(n407), .ZN(n400) );
  XNOR2_X1 U457 ( .A(n385), .B(n465), .ZN(n664) );
  INV_X1 U458 ( .A(n410), .ZN(n381) );
  XNOR2_X1 U459 ( .A(n374), .B(n373), .ZN(n768) );
  INV_X1 U460 ( .A(KEYINPUT40), .ZN(n373) );
  XNOR2_X1 U461 ( .A(KEYINPUT36), .B(KEYINPUT89), .ZN(n621) );
  INV_X1 U462 ( .A(KEYINPUT35), .ZN(n557) );
  XOR2_X1 U463 ( .A(KEYINPUT107), .B(n593), .Z(n681) );
  AND2_X1 U464 ( .A1(n629), .A2(KEYINPUT2), .ZN(n361) );
  AND2_X1 U465 ( .A1(n661), .A2(n565), .ZN(n362) );
  AND2_X1 U466 ( .A1(n565), .A2(KEYINPUT44), .ZN(n363) );
  INV_X1 U467 ( .A(KEYINPUT64), .ZN(n409) );
  XOR2_X1 U468 ( .A(KEYINPUT70), .B(G469), .Z(n364) );
  XNOR2_X1 U469 ( .A(n455), .B(n454), .ZN(n365) );
  NAND2_X1 U470 ( .A1(n559), .A2(n707), .ZN(n579) );
  AND2_X1 U471 ( .A1(n695), .A2(n415), .ZN(n366) );
  AND2_X2 U472 ( .A1(n410), .A2(n408), .ZN(n662) );
  AND2_X1 U473 ( .A1(n412), .A2(n695), .ZN(n367) );
  OR2_X1 U474 ( .A1(n551), .A2(n706), .ZN(n392) );
  AND2_X1 U475 ( .A1(n402), .A2(n403), .ZN(n368) );
  XOR2_X1 U476 ( .A(KEYINPUT90), .B(KEYINPUT33), .Z(n369) );
  XOR2_X1 U477 ( .A(KEYINPUT86), .B(KEYINPUT48), .Z(n370) );
  XOR2_X1 U478 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n371) );
  AND2_X1 U479 ( .A1(n631), .A2(KEYINPUT64), .ZN(n372) );
  NAND2_X1 U480 ( .A1(n626), .A2(n593), .ZN(n374) );
  NAND2_X1 U481 ( .A1(n380), .A2(n379), .ZN(n378) );
  NOR2_X1 U482 ( .A1(n735), .A2(n381), .ZN(n738) );
  NAND2_X1 U483 ( .A1(n382), .A2(n588), .ZN(n592) );
  NAND2_X1 U484 ( .A1(n571), .A2(n382), .ZN(n572) );
  INV_X1 U485 ( .A(n383), .ZN(n712) );
  NAND2_X1 U486 ( .A1(n383), .A2(n588), .ZN(n542) );
  NAND2_X1 U487 ( .A1(n564), .A2(n383), .ZN(n661) );
  XNOR2_X1 U488 ( .A(n430), .B(n429), .ZN(n385) );
  INV_X1 U489 ( .A(n392), .ZN(n388) );
  XNOR2_X2 U490 ( .A(n715), .B(n466), .ZN(n580) );
  NAND2_X1 U491 ( .A1(n396), .A2(n395), .ZN(n398) );
  NAND2_X1 U492 ( .A1(n362), .A2(KEYINPUT65), .ZN(n395) );
  NAND2_X1 U493 ( .A1(n397), .A2(n362), .ZN(n396) );
  NOR2_X1 U494 ( .A1(n766), .A2(KEYINPUT44), .ZN(n397) );
  NAND2_X1 U495 ( .A1(n359), .A2(n629), .ZN(n401) );
  NAND2_X1 U496 ( .A1(n399), .A2(n359), .ZN(n402) );
  AND2_X1 U497 ( .A1(n629), .A2(n372), .ZN(n399) );
  AND2_X1 U498 ( .A1(n630), .A2(n409), .ZN(n407) );
  INV_X1 U499 ( .A(n495), .ZN(n415) );
  NAND2_X1 U500 ( .A1(n547), .A2(n495), .ZN(n416) );
  NAND2_X1 U501 ( .A1(n608), .A2(n500), .ZN(n501) );
  NAND2_X1 U502 ( .A1(n661), .A2(n363), .ZN(n418) );
  NAND2_X1 U503 ( .A1(n420), .A2(n419), .ZN(n566) );
  INV_X1 U504 ( .A(n766), .ZN(n419) );
  NAND2_X1 U505 ( .A1(n559), .A2(n421), .ZN(n563) );
  XNOR2_X1 U506 ( .A(n501), .B(KEYINPUT0), .ZN(n552) );
  XNOR2_X2 U507 ( .A(n561), .B(G472), .ZN(n715) );
  XNOR2_X1 U508 ( .A(KEYINPUT109), .B(KEYINPUT28), .ZN(n423) );
  AND2_X1 U509 ( .A1(n600), .A2(n550), .ZN(n424) );
  OR2_X1 U510 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n425) );
  XNOR2_X1 U511 ( .A(KEYINPUT23), .B(KEYINPUT93), .ZN(n437) );
  BUF_X1 U512 ( .A(n552), .Z(n567) );
  NOR2_X1 U513 ( .A1(n598), .A2(n597), .ZN(n599) );
  XNOR2_X1 U514 ( .A(n447), .B(n446), .ZN(n448) );
  NOR2_X1 U515 ( .A1(n575), .A2(n576), .ZN(n593) );
  XNOR2_X1 U516 ( .A(n622), .B(n621), .ZN(n624) );
  XOR2_X1 U517 ( .A(KEYINPUT79), .B(n754), .Z(n430) );
  NAND2_X1 U518 ( .A1(G227), .A2(n762), .ZN(n427) );
  XNOR2_X1 U519 ( .A(G107), .B(G104), .ZN(n426) );
  XNOR2_X1 U520 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U521 ( .A(G110), .B(G101), .ZN(n473) );
  XNOR2_X1 U522 ( .A(n428), .B(n473), .ZN(n429) );
  INV_X1 U523 ( .A(G146), .ZN(n434) );
  INV_X1 U524 ( .A(KEYINPUT67), .ZN(n435) );
  XNOR2_X1 U525 ( .A(n435), .B(KEYINPUT1), .ZN(n436) );
  INV_X1 U526 ( .A(n551), .ZN(n623) );
  INV_X1 U527 ( .A(n623), .ZN(n707) );
  XNOR2_X1 U528 ( .A(n753), .B(n437), .ZN(n439) );
  INV_X1 U529 ( .A(KEYINPUT78), .ZN(n438) );
  XNOR2_X1 U530 ( .A(n439), .B(n438), .ZN(n449) );
  NAND2_X1 U531 ( .A1(n762), .A2(G234), .ZN(n441) );
  XNOR2_X1 U532 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n440) );
  XNOR2_X1 U533 ( .A(n441), .B(n440), .ZN(n509) );
  NAND2_X1 U534 ( .A1(n509), .A2(G221), .ZN(n445) );
  XOR2_X1 U535 ( .A(KEYINPUT24), .B(G140), .Z(n443) );
  XNOR2_X1 U536 ( .A(G137), .B(G110), .ZN(n442) );
  XNOR2_X1 U537 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n447) );
  XNOR2_X1 U539 ( .A(G128), .B(G119), .ZN(n446) );
  XNOR2_X1 U540 ( .A(n449), .B(n448), .ZN(n634) );
  INV_X1 U541 ( .A(G902), .ZN(n527) );
  NAND2_X1 U542 ( .A1(n634), .A2(n527), .ZN(n456) );
  XOR2_X1 U543 ( .A(KEYINPUT94), .B(KEYINPUT77), .Z(n452) );
  XNOR2_X1 U544 ( .A(G902), .B(KEYINPUT15), .ZN(n487) );
  NAND2_X1 U545 ( .A1(G234), .A2(n487), .ZN(n450) );
  XNOR2_X1 U546 ( .A(KEYINPUT20), .B(n450), .ZN(n530) );
  NAND2_X1 U547 ( .A1(G217), .A2(n530), .ZN(n451) );
  XNOR2_X1 U548 ( .A(n452), .B(n451), .ZN(n455) );
  XOR2_X1 U549 ( .A(KEYINPUT95), .B(KEYINPUT76), .Z(n453) );
  XNOR2_X1 U550 ( .A(KEYINPUT25), .B(n453), .ZN(n454) );
  OR2_X1 U551 ( .A1(n707), .A2(n712), .ZN(n468) );
  XOR2_X1 U552 ( .A(KEYINPUT74), .B(KEYINPUT5), .Z(n458) );
  XNOR2_X1 U553 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U554 ( .A(KEYINPUT3), .B(G119), .ZN(n474) );
  XNOR2_X1 U555 ( .A(n459), .B(n474), .ZN(n463) );
  NOR2_X1 U556 ( .A1(G953), .A2(G237), .ZN(n518) );
  NAND2_X1 U557 ( .A1(n518), .A2(G210), .ZN(n461) );
  XNOR2_X1 U558 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U559 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U560 ( .A(n465), .B(n464), .ZN(n655) );
  INV_X1 U561 ( .A(KEYINPUT6), .ZN(n466) );
  XNOR2_X1 U562 ( .A(n580), .B(KEYINPUT80), .ZN(n467) );
  NOR2_X1 U563 ( .A1(n468), .A2(n467), .ZN(n536) );
  INV_X1 U564 ( .A(G107), .ZN(n469) );
  XNOR2_X1 U565 ( .A(n470), .B(n469), .ZN(n508) );
  INV_X1 U566 ( .A(n508), .ZN(n472) );
  XNOR2_X1 U567 ( .A(n515), .B(KEYINPUT16), .ZN(n471) );
  XNOR2_X1 U568 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U569 ( .A(n474), .B(n473), .ZN(n475) );
  XNOR2_X1 U570 ( .A(n476), .B(n475), .ZN(n742) );
  NAND2_X1 U571 ( .A1(n762), .A2(G224), .ZN(n477) );
  XNOR2_X1 U572 ( .A(n478), .B(n477), .ZN(n480) );
  XNOR2_X1 U573 ( .A(n480), .B(n479), .ZN(n485) );
  INV_X1 U574 ( .A(n481), .ZN(n483) );
  XNOR2_X1 U575 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U577 ( .A(n742), .B(n486), .ZN(n640) );
  INV_X1 U578 ( .A(n487), .ZN(n631) );
  INV_X1 U579 ( .A(G237), .ZN(n488) );
  NAND2_X1 U580 ( .A1(n527), .A2(n488), .ZN(n493) );
  NAND2_X1 U581 ( .A1(n493), .A2(G210), .ZN(n490) );
  INV_X1 U582 ( .A(KEYINPUT91), .ZN(n489) );
  XNOR2_X1 U583 ( .A(n490), .B(n489), .ZN(n491) );
  NAND2_X1 U584 ( .A1(n493), .A2(G214), .ZN(n695) );
  INV_X1 U585 ( .A(KEYINPUT75), .ZN(n494) );
  XNOR2_X1 U586 ( .A(n494), .B(KEYINPUT19), .ZN(n495) );
  NAND2_X1 U587 ( .A1(G234), .A2(G237), .ZN(n497) );
  INV_X1 U588 ( .A(KEYINPUT14), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n497), .B(n496), .ZN(n726) );
  NAND2_X1 U590 ( .A1(G953), .A2(G902), .ZN(n538) );
  NOR2_X1 U591 ( .A1(G898), .A2(n538), .ZN(n498) );
  NOR2_X1 U592 ( .A1(n498), .A2(n540), .ZN(n499) );
  NOR2_X1 U593 ( .A1(n726), .A2(n499), .ZN(n500) );
  INV_X1 U594 ( .A(n552), .ZN(n571) );
  XOR2_X1 U595 ( .A(KEYINPUT105), .B(KEYINPUT104), .Z(n503) );
  XNOR2_X1 U596 ( .A(KEYINPUT7), .B(KEYINPUT103), .ZN(n502) );
  XNOR2_X1 U597 ( .A(n503), .B(n502), .ZN(n507) );
  XNOR2_X1 U598 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U599 ( .A(n507), .B(n506), .Z(n512) );
  NAND2_X1 U600 ( .A1(G217), .A2(n509), .ZN(n510) );
  XNOR2_X1 U601 ( .A(n508), .B(n510), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n512), .B(n511), .ZN(n638) );
  NAND2_X1 U603 ( .A1(n638), .A2(n527), .ZN(n513) );
  XNOR2_X1 U604 ( .A(n513), .B(G478), .ZN(n576) );
  INV_X1 U605 ( .A(n514), .ZN(n516) );
  XNOR2_X1 U606 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U607 ( .A(n517), .B(n753), .ZN(n526) );
  XOR2_X1 U608 ( .A(KEYINPUT100), .B(KEYINPUT12), .Z(n520) );
  NAND2_X1 U609 ( .A1(G214), .A2(n518), .ZN(n519) );
  XNOR2_X1 U610 ( .A(n520), .B(n519), .ZN(n524) );
  XOR2_X1 U611 ( .A(KEYINPUT11), .B(KEYINPUT101), .Z(n522) );
  XNOR2_X1 U612 ( .A(G143), .B(G122), .ZN(n521) );
  XNOR2_X1 U613 ( .A(n522), .B(n521), .ZN(n523) );
  XOR2_X1 U614 ( .A(n524), .B(n523), .Z(n525) );
  XNOR2_X1 U615 ( .A(n526), .B(n525), .ZN(n649) );
  NAND2_X1 U616 ( .A1(n649), .A2(n527), .ZN(n529) );
  XNOR2_X1 U617 ( .A(KEYINPUT13), .B(G475), .ZN(n528) );
  XNOR2_X1 U618 ( .A(n529), .B(n528), .ZN(n575) );
  INV_X1 U619 ( .A(n575), .ZN(n555) );
  NOR2_X1 U620 ( .A1(n576), .A2(n555), .ZN(n600) );
  NAND2_X1 U621 ( .A1(n530), .A2(G221), .ZN(n532) );
  INV_X1 U622 ( .A(KEYINPUT21), .ZN(n531) );
  XNOR2_X1 U623 ( .A(n532), .B(n531), .ZN(n711) );
  XNOR2_X1 U624 ( .A(n711), .B(KEYINPUT96), .ZN(n550) );
  NAND2_X1 U625 ( .A1(n571), .A2(n424), .ZN(n535) );
  INV_X1 U626 ( .A(KEYINPUT72), .ZN(n533) );
  XNOR2_X1 U627 ( .A(n533), .B(KEYINPUT22), .ZN(n534) );
  NAND2_X1 U628 ( .A1(n536), .A2(n559), .ZN(n537) );
  XNOR2_X1 U629 ( .A(n537), .B(KEYINPUT32), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(G119), .ZN(G21) );
  INV_X1 U631 ( .A(n711), .ZN(n543) );
  NOR2_X1 U632 ( .A1(G900), .A2(n538), .ZN(n539) );
  NOR2_X1 U633 ( .A1(n540), .A2(n539), .ZN(n541) );
  NOR2_X1 U634 ( .A1(n541), .A2(n726), .ZN(n588) );
  NAND2_X1 U635 ( .A1(n595), .A2(n681), .ZN(n544) );
  NOR2_X1 U636 ( .A1(n360), .A2(n544), .ZN(n620) );
  NAND2_X1 U637 ( .A1(n620), .A2(n695), .ZN(n545) );
  NOR2_X1 U638 ( .A1(n623), .A2(n545), .ZN(n546) );
  XOR2_X1 U639 ( .A(n546), .B(KEYINPUT43), .Z(n549) );
  BUF_X1 U640 ( .A(n547), .Z(n548) );
  NAND2_X1 U641 ( .A1(n549), .A2(n548), .ZN(n627) );
  XNOR2_X1 U642 ( .A(n627), .B(G140), .ZN(G42) );
  NAND2_X1 U643 ( .A1(n550), .A2(n712), .ZN(n706) );
  XNOR2_X1 U644 ( .A(KEYINPUT71), .B(KEYINPUT34), .ZN(n553) );
  XNOR2_X1 U645 ( .A(n554), .B(n553), .ZN(n556) );
  NAND2_X1 U646 ( .A1(n576), .A2(n555), .ZN(n612) );
  INV_X1 U647 ( .A(KEYINPUT66), .ZN(n562) );
  XNOR2_X1 U648 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U649 ( .A1(n566), .A2(n425), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n388), .A2(n715), .ZN(n718) );
  NOR2_X1 U651 ( .A1(n718), .A2(n567), .ZN(n570) );
  XOR2_X1 U652 ( .A(KEYINPUT99), .B(KEYINPUT31), .Z(n568) );
  XNOR2_X1 U653 ( .A(KEYINPUT98), .B(n568), .ZN(n569) );
  XNOR2_X1 U654 ( .A(n570), .B(n569), .ZN(n689) );
  XNOR2_X1 U655 ( .A(KEYINPUT97), .B(n572), .ZN(n574) );
  INV_X1 U656 ( .A(n715), .ZN(n573) );
  NAND2_X1 U657 ( .A1(n574), .A2(n573), .ZN(n671) );
  NAND2_X1 U658 ( .A1(n689), .A2(n671), .ZN(n578) );
  AND2_X1 U659 ( .A1(n576), .A2(n575), .ZN(n676) );
  NOR2_X1 U660 ( .A1(n593), .A2(n676), .ZN(n701) );
  INV_X1 U661 ( .A(n701), .ZN(n577) );
  NAND2_X1 U662 ( .A1(n578), .A2(n577), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n579), .A2(n580), .ZN(n581) );
  XNOR2_X1 U664 ( .A(n581), .B(KEYINPUT88), .ZN(n582) );
  NAND2_X1 U665 ( .A1(n582), .A2(n712), .ZN(n669) );
  NAND2_X1 U666 ( .A1(n583), .A2(n669), .ZN(n584) );
  XOR2_X1 U667 ( .A(KEYINPUT30), .B(KEYINPUT108), .Z(n590) );
  NAND2_X1 U668 ( .A1(n695), .A2(n594), .ZN(n589) );
  XOR2_X1 U669 ( .A(n590), .B(n589), .Z(n591) );
  XNOR2_X1 U670 ( .A(n548), .B(KEYINPUT38), .ZN(n696) );
  XNOR2_X1 U671 ( .A(n596), .B(n423), .ZN(n597) );
  INV_X1 U672 ( .A(n609), .ZN(n603) );
  INV_X1 U673 ( .A(n600), .ZN(n699) );
  NAND2_X1 U674 ( .A1(n696), .A2(n695), .ZN(n700) );
  NOR2_X1 U675 ( .A1(n699), .A2(n700), .ZN(n602) );
  XOR2_X1 U676 ( .A(KEYINPUT41), .B(KEYINPUT111), .Z(n601) );
  XNOR2_X1 U677 ( .A(n602), .B(n601), .ZN(n736) );
  NOR2_X1 U678 ( .A1(n603), .A2(n736), .ZN(n605) );
  XNOR2_X1 U679 ( .A(KEYINPUT112), .B(KEYINPUT42), .ZN(n604) );
  XNOR2_X1 U680 ( .A(n605), .B(n604), .ZN(n767) );
  NOR2_X1 U681 ( .A1(n768), .A2(n767), .ZN(n606) );
  NAND2_X1 U682 ( .A1(n609), .A2(n608), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n607), .B(KEYINPUT47), .ZN(n611) );
  AND2_X1 U684 ( .A1(n609), .A2(n608), .ZN(n682) );
  NAND2_X1 U685 ( .A1(n682), .A2(n701), .ZN(n610) );
  NAND2_X1 U686 ( .A1(n611), .A2(n610), .ZN(n618) );
  NOR2_X1 U687 ( .A1(n612), .A2(n548), .ZN(n613) );
  AND2_X1 U688 ( .A1(n614), .A2(n613), .ZN(n679) );
  NAND2_X1 U689 ( .A1(KEYINPUT47), .A2(n701), .ZN(n615) );
  XNOR2_X1 U690 ( .A(KEYINPUT83), .B(n615), .ZN(n616) );
  NOR2_X1 U691 ( .A1(n679), .A2(n616), .ZN(n617) );
  NAND2_X1 U692 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U693 ( .A(n619), .B(KEYINPUT73), .ZN(n625) );
  NAND2_X1 U694 ( .A1(n620), .A2(n367), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n624), .A2(n623), .ZN(n692) );
  NAND2_X1 U696 ( .A1(n626), .A2(n676), .ZN(n693) );
  AND2_X1 U697 ( .A1(n627), .A2(n693), .ZN(n628) );
  INV_X1 U698 ( .A(KEYINPUT2), .ZN(n630) );
  NAND2_X1 U699 ( .A1(n662), .A2(G217), .ZN(n633) );
  XOR2_X1 U700 ( .A(n634), .B(n633), .Z(n636) );
  INV_X1 U701 ( .A(G952), .ZN(n635) );
  NAND2_X1 U702 ( .A1(n635), .A2(G953), .ZN(n658) );
  INV_X1 U703 ( .A(n658), .ZN(n667) );
  NOR2_X1 U704 ( .A1(n636), .A2(n667), .ZN(G66) );
  NAND2_X1 U705 ( .A1(n662), .A2(G478), .ZN(n637) );
  XOR2_X1 U706 ( .A(n638), .B(n637), .Z(n639) );
  NOR2_X1 U707 ( .A1(n639), .A2(n667), .ZN(G63) );
  NAND2_X1 U708 ( .A1(n662), .A2(G210), .ZN(n644) );
  XNOR2_X1 U709 ( .A(KEYINPUT82), .B(KEYINPUT54), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n641), .B(KEYINPUT55), .ZN(n642) );
  XNOR2_X1 U711 ( .A(n640), .B(n642), .ZN(n643) );
  XNOR2_X1 U712 ( .A(n644), .B(n643), .ZN(n645) );
  NAND2_X1 U713 ( .A1(n645), .A2(n658), .ZN(n647) );
  XNOR2_X1 U714 ( .A(KEYINPUT85), .B(KEYINPUT56), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n647), .B(n646), .ZN(G51) );
  NAND2_X1 U716 ( .A1(n662), .A2(G475), .ZN(n651) );
  XOR2_X1 U717 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n648) );
  XNOR2_X1 U718 ( .A(n649), .B(n648), .ZN(n650) );
  XNOR2_X1 U719 ( .A(n651), .B(n650), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n652), .A2(n658), .ZN(n654) );
  INV_X1 U721 ( .A(KEYINPUT60), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(G60) );
  NAND2_X1 U723 ( .A1(n662), .A2(G472), .ZN(n657) );
  XOR2_X1 U724 ( .A(KEYINPUT62), .B(n655), .Z(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(n659) );
  NAND2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(n660), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U728 ( .A(n661), .B(G110), .ZN(G12) );
  NAND2_X1 U729 ( .A1(n662), .A2(G469), .ZN(n666) );
  XOR2_X1 U730 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n663) );
  XNOR2_X1 U731 ( .A(n664), .B(n663), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n666), .B(n665), .ZN(n668) );
  NOR2_X1 U733 ( .A1(n668), .A2(n667), .ZN(G54) );
  XNOR2_X1 U734 ( .A(G101), .B(n669), .ZN(G3) );
  INV_X1 U735 ( .A(n681), .ZN(n686) );
  NOR2_X1 U736 ( .A1(n686), .A2(n671), .ZN(n670) );
  XOR2_X1 U737 ( .A(G104), .B(n670), .Z(G6) );
  INV_X1 U738 ( .A(n676), .ZN(n688) );
  NOR2_X1 U739 ( .A1(n671), .A2(n688), .ZN(n675) );
  XOR2_X1 U740 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n673) );
  XNOR2_X1 U741 ( .A(G107), .B(KEYINPUT113), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n673), .B(n672), .ZN(n674) );
  XNOR2_X1 U743 ( .A(n675), .B(n674), .ZN(G9) );
  XOR2_X1 U744 ( .A(G128), .B(KEYINPUT29), .Z(n678) );
  NAND2_X1 U745 ( .A1(n682), .A2(n676), .ZN(n677) );
  XNOR2_X1 U746 ( .A(n678), .B(n677), .ZN(G30) );
  XOR2_X1 U747 ( .A(G143), .B(n679), .Z(n680) );
  XNOR2_X1 U748 ( .A(KEYINPUT114), .B(n680), .ZN(G45) );
  XOR2_X1 U749 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n684) );
  NAND2_X1 U750 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U751 ( .A(n684), .B(n683), .ZN(n685) );
  XNOR2_X1 U752 ( .A(G146), .B(n685), .ZN(G48) );
  NOR2_X1 U753 ( .A1(n689), .A2(n686), .ZN(n687) );
  XOR2_X1 U754 ( .A(G113), .B(n687), .Z(G15) );
  NOR2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n690) );
  XOR2_X1 U756 ( .A(G116), .B(n690), .Z(G18) );
  XOR2_X1 U757 ( .A(G125), .B(KEYINPUT37), .Z(n691) );
  XNOR2_X1 U758 ( .A(n692), .B(n691), .ZN(G27) );
  XNOR2_X1 U759 ( .A(G134), .B(n693), .ZN(G36) );
  NOR2_X1 U760 ( .A1(n696), .A2(n695), .ZN(n697) );
  XOR2_X1 U761 ( .A(KEYINPUT119), .B(n697), .Z(n698) );
  NOR2_X1 U762 ( .A1(n699), .A2(n698), .ZN(n703) );
  NOR2_X1 U763 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U764 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n694), .A2(n704), .ZN(n705) );
  XNOR2_X1 U766 ( .A(n705), .B(KEYINPUT120), .ZN(n723) );
  XOR2_X1 U767 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n709) );
  NAND2_X1 U768 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U769 ( .A(n709), .B(n708), .ZN(n710) );
  XNOR2_X1 U770 ( .A(n710), .B(KEYINPUT117), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n712), .A2(n711), .ZN(n713) );
  XOR2_X1 U772 ( .A(KEYINPUT49), .B(n713), .Z(n714) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U774 ( .A1(n717), .A2(n716), .ZN(n719) );
  NAND2_X1 U775 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U776 ( .A(KEYINPUT51), .B(n720), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n736), .A2(n721), .ZN(n722) );
  NOR2_X1 U778 ( .A1(n723), .A2(n722), .ZN(n724) );
  XNOR2_X1 U779 ( .A(n724), .B(KEYINPUT52), .ZN(n725) );
  NOR2_X1 U780 ( .A1(n726), .A2(n725), .ZN(n727) );
  NAND2_X1 U781 ( .A1(n727), .A2(G952), .ZN(n728) );
  XNOR2_X1 U782 ( .A(KEYINPUT121), .B(n728), .ZN(n729) );
  NOR2_X1 U783 ( .A1(G953), .A2(n729), .ZN(n740) );
  NAND2_X1 U784 ( .A1(n632), .A2(n630), .ZN(n733) );
  NAND2_X1 U785 ( .A1(n730), .A2(n630), .ZN(n731) );
  XNOR2_X1 U786 ( .A(n731), .B(KEYINPUT84), .ZN(n732) );
  AND2_X1 U787 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U788 ( .A(KEYINPUT81), .B(n734), .ZN(n735) );
  NOR2_X1 U789 ( .A1(n694), .A2(n736), .ZN(n737) );
  NOR2_X1 U790 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U791 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U792 ( .A(KEYINPUT53), .B(n741), .Z(G75) );
  XNOR2_X1 U793 ( .A(n742), .B(KEYINPUT124), .ZN(n744) );
  NOR2_X1 U794 ( .A1(G898), .A2(n762), .ZN(n743) );
  NOR2_X1 U795 ( .A1(n744), .A2(n743), .ZN(n745) );
  XOR2_X1 U796 ( .A(KEYINPUT125), .B(n745), .Z(n752) );
  NAND2_X1 U797 ( .A1(n359), .A2(n762), .ZN(n750) );
  XOR2_X1 U798 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n747) );
  NAND2_X1 U799 ( .A1(G224), .A2(G953), .ZN(n746) );
  XNOR2_X1 U800 ( .A(n747), .B(n746), .ZN(n748) );
  NAND2_X1 U801 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U802 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U803 ( .A(n752), .B(n751), .ZN(G69) );
  XNOR2_X1 U804 ( .A(n753), .B(KEYINPUT126), .ZN(n757) );
  XNOR2_X1 U805 ( .A(n755), .B(n754), .ZN(n756) );
  XOR2_X1 U806 ( .A(n757), .B(n756), .Z(n760) );
  XNOR2_X1 U807 ( .A(G227), .B(n760), .ZN(n758) );
  NAND2_X1 U808 ( .A1(G900), .A2(n758), .ZN(n759) );
  NAND2_X1 U809 ( .A1(n759), .A2(G953), .ZN(n765) );
  XOR2_X1 U810 ( .A(n760), .B(n730), .Z(n761) );
  XNOR2_X1 U811 ( .A(n761), .B(KEYINPUT127), .ZN(n763) );
  NAND2_X1 U812 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U813 ( .A1(n765), .A2(n764), .ZN(G72) );
  XOR2_X1 U814 ( .A(G122), .B(n766), .Z(G24) );
  XOR2_X1 U815 ( .A(n767), .B(G137), .Z(G39) );
  XOR2_X1 U816 ( .A(n768), .B(G131), .Z(G33) );
endmodule

