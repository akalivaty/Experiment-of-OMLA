//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 1 1 0 1 1 1 0 1 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(KEYINPUT78), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT72), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G137), .ZN(new_n190));
  AND2_X1   g004(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n191));
  NOR2_X1   g005(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n190), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G131), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT64), .A2(KEYINPUT11), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n195), .A2(G134), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n193), .A2(new_n194), .A3(new_n198), .A4(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G131), .B1(new_n190), .B2(new_n199), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT70), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n201), .A2(KEYINPUT70), .A3(new_n202), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT66), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  AOI21_X1  g026(.A(G128), .B1(new_n210), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(KEYINPUT1), .A3(G146), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n208), .B1(new_n213), .B2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n214), .B(KEYINPUT66), .C1(new_n217), .C2(G128), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  AND4_X1   g034(.A1(new_n220), .A2(new_n210), .A3(new_n212), .A4(G128), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(KEYINPUT71), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT71), .ZN(new_n224));
  AOI211_X1 g038(.A(new_n224), .B(new_n221), .C1(new_n216), .C2(new_n218), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n207), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT30), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n199), .B1(new_n196), .B2(new_n197), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n194), .B1(new_n228), .B2(new_n193), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(new_n201), .ZN(new_n231));
  NAND2_X1  g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n217), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT0), .B(G128), .Z(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(new_n217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n227), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  OAI21_X1  g051(.A(new_n188), .B1(new_n226), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT2), .ZN(new_n239));
  INV_X1    g053(.A(G113), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n239), .A2(new_n240), .A3(KEYINPUT67), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT67), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n242), .B1(KEYINPUT2), .B2(G113), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n239), .A2(new_n240), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G116), .B(G119), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n245), .B1(new_n243), .B2(new_n241), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(KEYINPUT68), .ZN(new_n253));
  OAI21_X1  g067(.A(KEYINPUT69), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n250), .B1(new_n247), .B2(new_n248), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT69), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n252), .A2(KEYINPUT68), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n252), .A2(new_n250), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n201), .ZN(new_n261));
  OAI211_X1 g075(.A(KEYINPUT65), .B(new_n235), .C1(new_n261), .C2(new_n229), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n221), .B1(new_n216), .B2(new_n218), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n262), .B1(new_n263), .B2(new_n203), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT65), .B1(new_n231), .B2(new_n235), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n227), .B1(new_n264), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n219), .A2(new_n222), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n224), .ZN(new_n268));
  AND3_X1   g082(.A1(new_n201), .A2(KEYINPUT70), .A3(new_n202), .ZN(new_n269));
  AOI21_X1  g083(.A(KEYINPUT70), .B1(new_n201), .B2(new_n202), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n268), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n273), .A2(KEYINPUT72), .A3(new_n236), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n238), .A2(new_n260), .A3(new_n266), .A4(new_n274), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n254), .A2(new_n258), .A3(new_n259), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n231), .A2(new_n235), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n273), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n275), .A2(new_n278), .ZN(new_n279));
  XOR2_X1   g093(.A(KEYINPUT73), .B(G237), .Z(new_n280));
  AND2_X1   g094(.A1(KEYINPUT74), .A2(G953), .ZN(new_n281));
  NOR2_X1   g095(.A1(KEYINPUT74), .A2(G953), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(G210), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n284), .B(KEYINPUT27), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT26), .B(G101), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n285), .B(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n273), .A2(new_n276), .A3(KEYINPUT28), .A4(new_n277), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n260), .B1(new_n264), .B2(new_n265), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n278), .A2(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n294), .A2(KEYINPUT76), .A3(new_n287), .A4(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n296), .A2(new_n287), .A3(new_n292), .A4(new_n291), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT76), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n289), .A2(new_n290), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n261), .A2(new_n229), .ZN(new_n302));
  INV_X1    g116(.A(new_n235), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR3_X1   g118(.A1(new_n226), .A2(new_n260), .A3(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n276), .B1(new_n273), .B2(new_n277), .ZN(new_n306));
  OAI211_X1 g120(.A(KEYINPUT77), .B(KEYINPUT28), .C1(new_n305), .C2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT77), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n296), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(new_n260), .B1(new_n226), .B2(new_n304), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n295), .B1(new_n310), .B2(new_n278), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n307), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g126(.A1(new_n288), .A2(new_n290), .ZN(new_n313));
  AOI21_X1  g127(.A(G902), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n301), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G472), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT31), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n278), .A2(new_n287), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n275), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n223), .A2(new_n225), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n304), .B1(new_n320), .B2(new_n271), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT28), .B1(new_n321), .B2(new_n276), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n288), .B1(new_n293), .B2(new_n322), .ZN(new_n323));
  AND2_X1   g137(.A1(new_n319), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT75), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n275), .A2(new_n318), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(KEYINPUT31), .ZN(new_n327));
  AOI211_X1 g141(.A(KEYINPUT75), .B(new_n317), .C1(new_n275), .C2(new_n318), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n324), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(G472), .A2(G902), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT32), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n316), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(KEYINPUT32), .B1(new_n329), .B2(new_n330), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n187), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT9), .B(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT80), .ZN(new_n339));
  OAI21_X1  g153(.A(G221), .B1(new_n339), .B2(G902), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(G469), .ZN(new_n342));
  INV_X1    g156(.A(G902), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(G104), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n345), .A2(KEYINPUT3), .A3(G107), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(KEYINPUT81), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT81), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(G104), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(G107), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n346), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n347), .A2(new_n349), .A3(G107), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(KEYINPUT82), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT82), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n347), .A2(new_n349), .A3(new_n356), .A4(G107), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G101), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n358), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n358), .ZN(new_n361));
  AND2_X1   g175(.A1(KEYINPUT83), .A2(G101), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n360), .A2(KEYINPUT4), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(KEYINPUT4), .A3(new_n362), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n235), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n352), .B1(G104), .B2(new_n351), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G101), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n360), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n320), .A2(KEYINPUT10), .A3(new_n369), .ZN(new_n370));
  OR3_X1    g184(.A1(new_n221), .A2(new_n213), .A3(new_n215), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n360), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT10), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g188(.A1(new_n366), .A2(new_n370), .A3(new_n302), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n283), .A2(G227), .ZN(new_n376));
  XOR2_X1   g190(.A(G110), .B(G140), .Z(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n375), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n366), .A2(new_n370), .A3(new_n374), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(new_n231), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n302), .A2(KEYINPUT84), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n267), .B1(new_n360), .B2(new_n368), .ZN(new_n384));
  INV_X1    g198(.A(new_n372), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT12), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT12), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n388), .B(new_n383), .C1(new_n384), .C2(new_n385), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n375), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  AOI22_X1  g204(.A1(new_n380), .A2(new_n382), .B1(new_n390), .B2(new_n378), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n344), .B1(new_n391), .B2(G469), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n379), .B1(new_n382), .B2(new_n375), .ZN(new_n393));
  AND4_X1   g207(.A1(new_n375), .A2(new_n387), .A3(new_n379), .A4(new_n389), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n342), .B(new_n343), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n341), .B1(new_n392), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G122), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n363), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n276), .B1(new_n400), .B2(new_n364), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n402));
  INV_X1    g216(.A(G116), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n403), .A2(KEYINPUT5), .A3(G119), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(new_n240), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n252), .A2(new_n250), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n360), .A2(new_n406), .A3(new_n368), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT85), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT85), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n360), .A2(new_n406), .A3(new_n409), .A4(new_n368), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n399), .B1(new_n401), .B2(new_n411), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n260), .B1(new_n363), .B2(new_n365), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n413), .A2(new_n398), .A3(new_n408), .A4(new_n410), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(KEYINPUT6), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n235), .A2(G125), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n416), .B1(new_n263), .B2(G125), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT86), .B(G224), .ZN(new_n418));
  INV_X1    g232(.A(G953), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n417), .B(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT6), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n422), .B(new_n399), .C1(new_n401), .C2(new_n411), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n415), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT87), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n407), .A2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n360), .A2(new_n406), .A3(KEYINPUT87), .A4(new_n368), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n426), .B(new_n427), .C1(new_n369), .C2(new_n406), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n398), .B(KEYINPUT8), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n420), .A2(KEYINPUT7), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n417), .B(new_n431), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n414), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  AND2_X1   g247(.A1(new_n433), .A2(new_n343), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n424), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(G210), .B1(G237), .B2(G902), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n436), .B(KEYINPUT88), .Z(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n435), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(G234), .A2(G237), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(G952), .A3(new_n419), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT21), .B(G898), .Z(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT94), .ZN(new_n443));
  INV_X1    g257(.A(new_n283), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n444), .A2(G902), .A3(new_n440), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n441), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n424), .A2(new_n434), .A3(new_n437), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n439), .A2(new_n446), .A3(new_n447), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n280), .A2(G214), .A3(new_n283), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n211), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n280), .A2(G143), .A3(G214), .A4(new_n283), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n451), .A2(new_n194), .A3(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n194), .B1(new_n451), .B2(new_n452), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT91), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n451), .A2(new_n452), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT91), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(new_n459), .A3(new_n453), .ZN(new_n460));
  XNOR2_X1  g274(.A(G125), .B(G140), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT19), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n461), .A2(KEYINPUT19), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n209), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n461), .A2(KEYINPUT16), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT16), .ZN(new_n467));
  INV_X1    g281(.A(G140), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n466), .A2(G146), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT92), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n465), .A2(KEYINPUT92), .A3(new_n470), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n456), .A2(new_n460), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(KEYINPUT18), .A2(G131), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n451), .A2(new_n452), .A3(new_n476), .ZN(new_n477));
  XNOR2_X1  g291(.A(new_n461), .B(new_n209), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n476), .B1(new_n451), .B2(new_n452), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT90), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n480), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n478), .A4(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n475), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G113), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(new_n345), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n466), .A2(new_n469), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n209), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n470), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n493), .B1(new_n455), .B2(KEYINPUT17), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n458), .A2(new_n453), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n494), .B1(new_n495), .B2(KEYINPUT17), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n485), .A2(new_n496), .A3(new_n488), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n490), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(G475), .A2(G902), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n500), .A2(KEYINPUT93), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT20), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT93), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n499), .B2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n498), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n500), .B1(new_n490), .B2(new_n497), .ZN(new_n507));
  XNOR2_X1  g321(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n497), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n488), .B1(new_n485), .B2(new_n496), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n343), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G475), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n211), .A2(G128), .ZN(new_n514));
  INV_X1    g328(.A(G128), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(G143), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n514), .A2(new_n516), .A3(new_n189), .ZN(new_n517));
  INV_X1    g331(.A(G122), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G116), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n403), .A2(G122), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(G107), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n519), .A2(new_n520), .A3(new_n351), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n517), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n514), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n516), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n514), .A2(new_n525), .ZN(new_n528));
  OAI21_X1  g342(.A(G134), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n403), .A2(KEYINPUT14), .A3(G122), .ZN(new_n531));
  OAI211_X1 g345(.A(G107), .B(new_n531), .C1(new_n521), .C2(KEYINPUT14), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n189), .B1(new_n514), .B2(new_n516), .ZN(new_n533));
  OAI211_X1 g347(.A(new_n532), .B(new_n523), .C1(new_n517), .C2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(new_n339), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n536), .A2(G217), .A3(new_n419), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G217), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n339), .A2(new_n539), .A3(G953), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n540), .A2(new_n530), .A3(new_n534), .ZN(new_n541));
  AOI21_X1  g355(.A(G902), .B1(new_n538), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G478), .ZN(new_n543));
  OR2_X1    g357(.A1(new_n543), .A2(KEYINPUT15), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n542), .A2(new_n544), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n509), .A2(new_n513), .A3(new_n548), .ZN(new_n549));
  NOR3_X1   g363(.A1(new_n397), .A2(new_n449), .A3(new_n549), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n315), .A2(G472), .B1(new_n329), .B2(new_n333), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n319), .A2(new_n323), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n326), .A2(KEYINPUT31), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n326), .A2(new_n325), .A3(KEYINPUT31), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n332), .B1(new_n556), .B2(new_n331), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(KEYINPUT78), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(G119), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n559), .A2(G128), .ZN(new_n560));
  OR2_X1    g374(.A1(new_n560), .A2(KEYINPUT79), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(KEYINPUT79), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(G128), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(KEYINPUT24), .B(G110), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n515), .A2(KEYINPUT23), .A3(G119), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n563), .B(new_n567), .C1(new_n560), .C2(KEYINPUT23), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n566), .B1(G110), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n461), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n569), .B(new_n470), .C1(G146), .C2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n568), .A2(G110), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n493), .B(new_n572), .C1(new_n565), .C2(new_n564), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n283), .A2(G221), .A3(G234), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT22), .B(G137), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n571), .A2(new_n573), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n571), .B2(new_n573), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n539), .B1(G234), .B2(new_n343), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G902), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NOR3_X1   g396(.A1(new_n577), .A2(new_n578), .A3(G902), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n583), .B(KEYINPUT25), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n582), .B1(new_n584), .B2(new_n580), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n337), .A2(new_n550), .A3(new_n558), .A4(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  INV_X1    g401(.A(G472), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n588), .B1(new_n329), .B2(new_n343), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n590));
  OR2_X1    g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n589), .A2(new_n590), .B1(new_n330), .B2(new_n329), .ZN(new_n592));
  AND2_X1   g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n585), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n397), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n508), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n488), .B1(new_n475), .B2(new_n485), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n510), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n597), .B1(new_n599), .B2(new_n500), .ZN(new_n600));
  AOI22_X1  g414(.A1(new_n600), .A2(new_n506), .B1(G475), .B2(new_n512), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT33), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n538), .A2(new_n541), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n538), .B2(new_n541), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n543), .A2(G902), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT96), .B1(new_n606), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n610), .B(new_n607), .C1(new_n604), .C2(new_n605), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n542), .A2(G478), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(KEYINPUT97), .ZN(new_n614));
  AOI22_X1  g428(.A1(new_n609), .A2(new_n611), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n602), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n617), .A2(new_n449), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n596), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT98), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT34), .B(G104), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n620), .B(new_n621), .ZN(G6));
  AOI21_X1  g436(.A(new_n508), .B1(new_n498), .B2(new_n499), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n499), .B(new_n508), .C1(new_n510), .C2(new_n598), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n513), .B(new_n547), .C1(new_n623), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n449), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n596), .A2(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT35), .B(G107), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G9));
  NAND2_X1  g444(.A1(new_n584), .A2(new_n580), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n571), .A2(new_n573), .ZN(new_n632));
  INV_X1    g446(.A(new_n576), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n633), .A2(KEYINPUT36), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n632), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(new_n581), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n550), .A2(new_n591), .A3(new_n592), .A4(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  INV_X1    g454(.A(new_n637), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n439), .A2(new_n447), .A3(new_n448), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n397), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n441), .B(KEYINPUT99), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n644), .B1(new_n445), .B2(G900), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n626), .A2(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n337), .A2(new_n643), .A3(new_n558), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G128), .ZN(G30));
  XNOR2_X1  g463(.A(new_n645), .B(KEYINPUT39), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n396), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(new_n651), .B(KEYINPUT40), .Z(new_n652));
  NAND2_X1  g466(.A1(new_n439), .A2(new_n448), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT38), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n602), .A2(new_n447), .A3(new_n547), .ZN(new_n655));
  NOR3_X1   g469(.A1(new_n654), .A2(new_n637), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n288), .B1(new_n275), .B2(new_n278), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n310), .A2(new_n288), .A3(new_n278), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n658), .A2(new_n343), .ZN(new_n659));
  OAI21_X1  g473(.A(G472), .B1(new_n657), .B2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n557), .A2(new_n334), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n652), .A2(new_n656), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT100), .B(G143), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G45));
  AOI211_X1 g478(.A(new_n615), .B(new_n646), .C1(new_n509), .C2(new_n513), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n337), .A2(new_n643), .A3(new_n558), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  AND3_X1   g481(.A1(new_n551), .A2(KEYINPUT78), .A3(new_n557), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT78), .B1(new_n551), .B2(new_n557), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT101), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n343), .B1(new_n393), .B2(new_n394), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G469), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n673), .A2(new_n340), .A3(new_n395), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n674), .A2(new_n594), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n670), .A2(new_n671), .A3(new_n618), .A4(new_n675), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n337), .A2(new_n675), .A3(new_n558), .A4(new_n618), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT101), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT41), .B(G113), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NAND4_X1  g495(.A1(new_n337), .A2(new_n675), .A3(new_n558), .A4(new_n627), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G116), .ZN(G18));
  NAND4_X1  g497(.A1(new_n509), .A2(new_n446), .A3(new_n513), .A4(new_n548), .ZN(new_n684));
  NOR3_X1   g498(.A1(new_n642), .A2(new_n674), .A3(new_n684), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n337), .A2(new_n558), .A3(new_n637), .A4(new_n685), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G119), .ZN(G21));
  NOR2_X1   g501(.A1(new_n655), .A2(new_n653), .ZN(new_n688));
  XOR2_X1   g502(.A(new_n585), .B(KEYINPUT102), .Z(new_n689));
  AND2_X1   g503(.A1(new_n553), .A2(new_n319), .ZN(new_n690));
  OR2_X1    g504(.A1(new_n312), .A2(new_n287), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n331), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n589), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n446), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n674), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n688), .A2(new_n689), .A3(new_n693), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G122), .ZN(G24));
  NOR3_X1   g511(.A1(new_n589), .A2(new_n641), .A3(new_n692), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n642), .A2(new_n674), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n698), .A2(new_n665), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G125), .ZN(G27));
  INV_X1    g515(.A(new_n447), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n439), .B2(new_n448), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n703), .A2(new_n665), .A3(new_n396), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n551), .A2(new_n557), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n704), .A2(new_n705), .A3(new_n689), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT42), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n703), .A2(new_n665), .A3(new_n396), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(KEYINPUT42), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n337), .A3(new_n558), .A4(new_n585), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n194), .ZN(G33));
  AND3_X1   g526(.A1(new_n703), .A2(new_n647), .A3(new_n396), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n337), .A2(new_n558), .A3(new_n713), .A4(new_n585), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  NOR2_X1   g529(.A1(KEYINPUT105), .A2(KEYINPUT43), .ZN(new_n716));
  XOR2_X1   g530(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n717));
  NAND2_X1  g531(.A1(new_n601), .A2(new_n616), .ZN(new_n718));
  MUX2_X1   g532(.A(new_n716), .B(new_n717), .S(new_n718), .Z(new_n719));
  OR3_X1    g533(.A1(new_n593), .A2(new_n719), .A3(new_n641), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT44), .ZN(new_n721));
  OR2_X1    g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n703), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n395), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n380), .A2(new_n382), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n390), .A2(new_n378), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT45), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(KEYINPUT103), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n342), .B1(new_n729), .B2(new_n730), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n344), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n726), .B1(new_n734), .B2(KEYINPUT46), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  OAI211_X1 g552(.A(new_n737), .B(new_n738), .C1(KEYINPUT46), .C2(new_n734), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n340), .ZN(new_n740));
  INV_X1    g554(.A(new_n650), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n725), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT106), .B(G137), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G39));
  INV_X1    g558(.A(new_n670), .ZN(new_n745));
  AND3_X1   g559(.A1(new_n703), .A2(new_n665), .A3(new_n594), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT47), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n740), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n739), .A2(KEYINPUT47), .A3(new_n340), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n747), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(new_n468), .ZN(G42));
  NOR2_X1   g566(.A1(new_n723), .A2(new_n674), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  NOR4_X1   g568(.A1(new_n754), .A2(new_n661), .A3(new_n594), .A4(new_n441), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n602), .A2(new_n616), .ZN(new_n756));
  NOR3_X1   g570(.A1(new_n719), .A2(new_n754), .A3(new_n644), .ZN(new_n757));
  AOI22_X1  g571(.A1(new_n755), .A2(new_n756), .B1(new_n757), .B2(new_n698), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n719), .A2(new_n644), .ZN(new_n759));
  AND2_X1   g573(.A1(new_n689), .A2(new_n693), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n674), .A2(new_n447), .ZN(new_n761));
  AND4_X1   g575(.A1(new_n654), .A2(new_n759), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n762), .A2(KEYINPUT50), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(KEYINPUT50), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n763), .A2(KEYINPUT111), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(KEYINPUT111), .B1(new_n763), .B2(new_n764), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n758), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n673), .A2(new_n395), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n749), .B(new_n750), .C1(new_n340), .C2(new_n770), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n760), .A3(new_n703), .A4(new_n759), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n767), .A2(new_n768), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n769), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n549), .B1(new_n601), .B2(new_n616), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n449), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n595), .A2(new_n591), .A3(new_n592), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n586), .A2(new_n638), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT107), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n586), .A2(new_n638), .A3(new_n780), .A4(KEYINPUT107), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n682), .A2(new_n686), .A3(new_n696), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n786), .B1(new_n676), .B2(new_n678), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n513), .B1(new_n623), .B2(new_n625), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n548), .A2(new_n645), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n703), .A2(new_n396), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n337), .A2(new_n558), .A3(new_n637), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n704), .A2(new_n698), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n714), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n711), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n785), .A2(new_n787), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n648), .A2(new_n700), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT52), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n641), .A2(KEYINPUT109), .A3(new_n645), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT109), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n800), .B1(new_n637), .B2(new_n646), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n397), .B1(new_n799), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n661), .A3(new_n688), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n797), .A2(new_n798), .A3(new_n666), .A4(new_n803), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n648), .A2(new_n666), .A3(new_n803), .A4(new_n700), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n777), .B1(new_n796), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n648), .A2(new_n700), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT52), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n796), .A2(new_n807), .A3(new_n777), .A4(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT54), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n804), .A2(new_n806), .A3(new_n811), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n785), .A2(new_n787), .A3(new_n795), .A4(KEYINPUT108), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n707), .A2(new_n710), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n682), .A2(new_n686), .A3(new_n696), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n714), .A2(new_n792), .A3(new_n793), .ZN(new_n820));
  AND4_X1   g634(.A1(new_n679), .A2(new_n818), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT108), .B1(new_n821), .B2(new_n785), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n777), .B1(new_n817), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT110), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n825), .B(new_n777), .C1(new_n817), .C2(new_n822), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n796), .A2(new_n807), .A3(new_n777), .ZN(new_n827));
  INV_X1    g641(.A(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n824), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n814), .B1(new_n829), .B2(KEYINPUT54), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n689), .A2(new_n705), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n757), .A2(new_n831), .ZN(new_n832));
  XNOR2_X1  g646(.A(new_n832), .B(KEYINPUT48), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n759), .A2(new_n699), .A3(new_n760), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n419), .A2(G952), .ZN(new_n835));
  INV_X1    g649(.A(new_n617), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n835), .B1(new_n755), .B2(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n834), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n758), .A2(KEYINPUT51), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n839), .B1(new_n763), .B2(new_n764), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(new_n772), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n776), .A2(new_n830), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(G952), .A2(G953), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n689), .A2(new_n447), .A3(new_n340), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n770), .A2(KEYINPUT49), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n844), .A2(new_n718), .A3(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n846), .B(new_n654), .C1(KEYINPUT49), .C2(new_n770), .ZN(new_n847));
  OAI22_X1  g661(.A1(new_n842), .A2(new_n843), .B1(new_n661), .B2(new_n847), .ZN(G75));
  NOR2_X1   g662(.A1(new_n796), .A2(new_n807), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(KEYINPUT53), .A3(new_n811), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n343), .B1(new_n850), .B2(new_n808), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n437), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n415), .A2(new_n423), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(new_n421), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT55), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(KEYINPUT56), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n852), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n855), .B1(new_n852), .B2(new_n857), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n283), .A2(G952), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(G51));
  XNOR2_X1  g675(.A(new_n344), .B(KEYINPUT57), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n863), .B1(new_n850), .B2(new_n808), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n862), .B1(new_n814), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n865), .B1(new_n393), .B2(new_n394), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n851), .A2(new_n732), .A3(new_n733), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n860), .B1(new_n866), .B2(new_n867), .ZN(G54));
  INV_X1    g682(.A(new_n860), .ZN(new_n869));
  NAND2_X1  g683(.A1(KEYINPUT58), .A2(G475), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT114), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n851), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n869), .B1(new_n872), .B2(new_n599), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT115), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(new_n872), .B2(new_n599), .ZN(new_n875));
  AOI211_X1 g689(.A(KEYINPUT115), .B(new_n498), .C1(new_n851), .C2(new_n871), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n873), .A2(new_n875), .A3(new_n876), .ZN(G60));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND2_X1  g692(.A1(G478), .A2(G902), .ZN(new_n879));
  XOR2_X1   g693(.A(new_n879), .B(KEYINPUT59), .Z(new_n880));
  OAI211_X1 g694(.A(new_n878), .B(new_n606), .C1(new_n830), .C2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n880), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n827), .B1(new_n823), .B2(KEYINPUT110), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n863), .B1(new_n884), .B2(new_n826), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n883), .B1(new_n885), .B2(new_n814), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n878), .B1(new_n886), .B2(new_n606), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n606), .A2(new_n880), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n814), .B2(new_n864), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT116), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n869), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n890), .B1(new_n889), .B2(new_n869), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n882), .A2(new_n887), .A3(new_n893), .ZN(G63));
  NAND2_X1  g708(.A1(G217), .A2(G902), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT118), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT60), .Z(new_n897));
  AOI21_X1  g711(.A(new_n897), .B1(new_n850), .B2(new_n808), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(new_n635), .ZN(new_n899));
  NOR2_X1   g713(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n860), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g715(.A(new_n899), .B(new_n901), .C1(new_n579), .C2(new_n898), .ZN(new_n902));
  NAND2_X1  g716(.A1(KEYINPUT119), .A2(KEYINPUT61), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n902), .B(new_n903), .ZN(G66));
  AOI21_X1  g718(.A(new_n419), .B1(new_n443), .B2(new_n418), .ZN(new_n905));
  XOR2_X1   g719(.A(new_n905), .B(KEYINPUT121), .Z(new_n906));
  NAND2_X1  g720(.A1(new_n785), .A2(new_n787), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT120), .Z(new_n908));
  AOI21_X1  g722(.A(new_n906), .B1(new_n908), .B2(new_n283), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n853), .B1(G898), .B2(new_n283), .ZN(new_n910));
  XOR2_X1   g724(.A(new_n909), .B(new_n910), .Z(G69));
  AOI21_X1  g725(.A(new_n283), .B1(G227), .B2(G900), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT124), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n238), .A2(new_n266), .A3(new_n274), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n463), .A2(new_n464), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n916), .B(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n918), .A2(new_n444), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(new_n750), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT47), .B1(new_n739), .B2(new_n340), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n745), .B(new_n746), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n740), .A2(new_n741), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n924), .A2(new_n722), .A3(new_n724), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n723), .A2(new_n651), .A3(new_n778), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n670), .A2(new_n585), .A3(new_n926), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n923), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n797), .A2(new_n662), .A3(new_n666), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT62), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n920), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n283), .A2(G900), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n933), .B(KEYINPUT123), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n831), .A2(new_n688), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n924), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n818), .A2(new_n714), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n797), .A2(new_n666), .ZN(new_n939));
  NOR2_X1   g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n923), .A2(new_n925), .A3(new_n937), .A4(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n935), .B1(new_n941), .B2(new_n283), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n914), .B(new_n915), .C1(new_n932), .C2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n923), .A2(new_n925), .A3(new_n927), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n919), .B1(new_n945), .B2(new_n930), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n751), .A2(new_n742), .ZN(new_n947));
  AOI211_X1 g761(.A(new_n939), .B(new_n938), .C1(new_n924), .C2(new_n936), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n444), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n946), .B1(new_n949), .B2(new_n935), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n915), .B1(new_n950), .B2(new_n914), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n913), .B1(new_n944), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n914), .B1(new_n932), .B2(new_n942), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(new_n943), .A3(new_n912), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n941), .B2(new_n908), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n279), .A2(new_n287), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n860), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n947), .A2(new_n931), .A3(new_n927), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n958), .B1(new_n962), .B2(new_n908), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n963), .A2(KEYINPUT125), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n657), .B1(new_n963), .B2(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n289), .A2(KEYINPUT126), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n326), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n289), .A2(KEYINPUT126), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n958), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT127), .Z(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n884), .B2(new_n826), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n966), .A2(new_n972), .ZN(G57));
endmodule


