

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738;

  NOR2_X1 U367 ( .A1(n497), .A2(n563), .ZN(n636) );
  INV_X2 U368 ( .A(G953), .ZN(n730) );
  NOR2_X1 U369 ( .A1(n737), .A2(n738), .ZN(n573) );
  INV_X1 U370 ( .A(n630), .ZN(n392) );
  XNOR2_X1 U371 ( .A(n443), .B(n442), .ZN(n563) );
  NOR2_X2 U372 ( .A1(n388), .A2(n386), .ZN(n446) );
  XNOR2_X2 U373 ( .A(n481), .B(n404), .ZN(n441) );
  NOR2_X1 U374 ( .A1(n378), .A2(KEYINPUT80), .ZN(n377) );
  AND2_X1 U375 ( .A1(n531), .A2(n385), .ZN(n529) );
  XNOR2_X1 U376 ( .A(n496), .B(n495), .ZN(n385) );
  XNOR2_X1 U377 ( .A(KEYINPUT22), .B(n510), .ZN(n518) );
  OR2_X1 U378 ( .A1(n511), .A2(n630), .ZN(n497) );
  XOR2_X2 U379 ( .A(G122), .B(G107), .Z(n477) );
  NOR2_X1 U380 ( .A1(n377), .A2(n376), .ZN(n375) );
  AND2_X1 U381 ( .A1(n374), .A2(n534), .ZN(n373) );
  NOR2_X1 U382 ( .A1(n585), .A2(n584), .ZN(n586) );
  NOR2_X1 U383 ( .A1(n518), .A2(n512), .ZN(n514) );
  NOR2_X1 U384 ( .A1(n645), .A2(n648), .ZN(n562) );
  OR2_X1 U385 ( .A1(n511), .A2(n391), .ZN(n390) );
  NAND2_X1 U386 ( .A1(n393), .A2(n387), .ZN(n386) );
  BUF_X1 U387 ( .A(n536), .Z(n551) );
  XNOR2_X1 U388 ( .A(n485), .B(n484), .ZN(n505) );
  OR2_X1 U389 ( .A1(n610), .A2(G902), .ZN(n413) );
  INV_X1 U390 ( .A(KEYINPUT33), .ZN(n445) );
  AND2_X1 U391 ( .A1(n359), .A2(n360), .ZN(n345) );
  NAND2_X1 U392 ( .A1(n375), .A2(n373), .ZN(n535) );
  INV_X1 U393 ( .A(n645), .ZN(n507) );
  XNOR2_X1 U394 ( .A(n433), .B(n434), .ZN(n448) );
  XNOR2_X1 U395 ( .A(n432), .B(n431), .ZN(n433) );
  INV_X1 U396 ( .A(KEYINPUT84), .ZN(n431) );
  XNOR2_X1 U397 ( .A(n528), .B(KEYINPUT81), .ZN(n358) );
  XNOR2_X1 U398 ( .A(n402), .B(G131), .ZN(n486) );
  INV_X1 U399 ( .A(KEYINPUT69), .ZN(n402) );
  NAND2_X1 U400 ( .A1(n505), .A2(n506), .ZN(n645) );
  XNOR2_X1 U401 ( .A(KEYINPUT83), .B(G110), .ZN(n409) );
  XNOR2_X1 U402 ( .A(n712), .B(n396), .ZN(n704) );
  XNOR2_X1 U403 ( .A(n398), .B(n397), .ZN(n396) );
  XNOR2_X1 U404 ( .A(n457), .B(n453), .ZN(n398) );
  NOR2_X1 U405 ( .A1(n664), .A2(KEYINPUT122), .ZN(n363) );
  INV_X1 U406 ( .A(KEYINPUT0), .ZN(n468) );
  XNOR2_X1 U407 ( .A(n423), .B(n422), .ZN(n425) );
  XNOR2_X1 U408 ( .A(n348), .B(n421), .ZN(n422) );
  NAND2_X1 U409 ( .A1(n701), .A2(n702), .ZN(n384) );
  INV_X1 U410 ( .A(n544), .ZN(n393) );
  XNOR2_X1 U411 ( .A(G116), .B(KEYINPUT3), .ZN(n430) );
  XNOR2_X1 U412 ( .A(G113), .B(G119), .ZN(n432) );
  XNOR2_X1 U413 ( .A(n487), .B(n488), .ZN(n372) );
  XNOR2_X1 U414 ( .A(G113), .B(G104), .ZN(n487) );
  XNOR2_X1 U415 ( .A(G122), .B(G143), .ZN(n488) );
  INV_X1 U416 ( .A(n486), .ZN(n370) );
  XNOR2_X1 U417 ( .A(KEYINPUT4), .B(G137), .ZN(n403) );
  INV_X1 U418 ( .A(G128), .ZN(n400) );
  XOR2_X1 U419 ( .A(KEYINPUT38), .B(n551), .Z(n642) );
  OR2_X1 U420 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U421 ( .A(n459), .B(n458), .ZN(n536) );
  NOR2_X1 U422 ( .A1(n704), .A2(n700), .ZN(n459) );
  XNOR2_X1 U423 ( .A(n492), .B(n366), .ZN(n506) );
  XNOR2_X1 U424 ( .A(n367), .B(KEYINPUT13), .ZN(n366) );
  NOR2_X1 U425 ( .A1(G902), .A2(n602), .ZN(n492) );
  INV_X1 U426 ( .A(G475), .ZN(n367) );
  XNOR2_X1 U427 ( .A(G128), .B(G110), .ZN(n420) );
  XNOR2_X1 U428 ( .A(G119), .B(G137), .ZN(n419) );
  XOR2_X1 U429 ( .A(KEYINPUT8), .B(n418), .Z(n476) );
  XNOR2_X1 U430 ( .A(n722), .B(n368), .ZN(n602) );
  XNOR2_X1 U431 ( .A(n371), .B(n369), .ZN(n368) );
  XNOR2_X1 U432 ( .A(n370), .B(n491), .ZN(n369) );
  XNOR2_X1 U433 ( .A(n372), .B(n489), .ZN(n371) );
  XNOR2_X1 U434 ( .A(n441), .B(KEYINPUT88), .ZN(n724) );
  XNOR2_X1 U435 ( .A(G107), .B(G101), .ZN(n406) );
  AND2_X1 U436 ( .A1(n598), .A2(n597), .ZN(n728) );
  XNOR2_X1 U437 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U438 ( .A(KEYINPUT30), .B(KEYINPUT103), .ZN(n554) );
  INV_X1 U439 ( .A(KEYINPUT97), .ZN(n483) );
  XOR2_X1 U440 ( .A(KEYINPUT94), .B(n506), .Z(n502) );
  XNOR2_X1 U441 ( .A(n399), .B(n448), .ZN(n712) );
  XNOR2_X1 U442 ( .A(n450), .B(n447), .ZN(n399) );
  XNOR2_X1 U443 ( .A(n477), .B(n449), .ZN(n450) );
  NAND2_X1 U444 ( .A1(n701), .A2(n355), .ZN(n604) );
  AND2_X1 U445 ( .A1(n361), .A2(n730), .ZN(n360) );
  NOR2_X1 U446 ( .A1(n593), .A2(n590), .ZN(n548) );
  XNOR2_X1 U447 ( .A(n523), .B(n522), .ZN(n736) );
  NAND2_X1 U448 ( .A1(n524), .A2(n520), .ZN(n523) );
  INV_X1 U449 ( .A(KEYINPUT31), .ZN(n379) );
  NOR2_X1 U450 ( .A1(n576), .A2(n575), .ZN(n689) );
  AND2_X1 U451 ( .A1(n700), .A2(G217), .ZN(n395) );
  NAND2_X1 U452 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U453 ( .A(n384), .B(n354), .ZN(n383) );
  AND2_X1 U454 ( .A1(n701), .A2(n700), .ZN(n346) );
  AND2_X1 U455 ( .A1(n532), .A2(KEYINPUT80), .ZN(n347) );
  XOR2_X1 U456 ( .A(n419), .B(KEYINPUT23), .Z(n348) );
  OR2_X1 U457 ( .A1(n708), .A2(G902), .ZN(n349) );
  XNOR2_X1 U458 ( .A(KEYINPUT19), .B(KEYINPUT68), .ZN(n350) );
  XNOR2_X1 U459 ( .A(KEYINPUT85), .B(KEYINPUT74), .ZN(n351) );
  XOR2_X1 U460 ( .A(KEYINPUT24), .B(KEYINPUT89), .Z(n352) );
  XOR2_X1 U461 ( .A(KEYINPUT17), .B(KEYINPUT73), .Z(n353) );
  INV_X1 U462 ( .A(KEYINPUT100), .ZN(n394) );
  XOR2_X1 U463 ( .A(n704), .B(n703), .Z(n354) );
  AND2_X1 U464 ( .A1(n700), .A2(G475), .ZN(n355) );
  AND2_X1 U465 ( .A1(n700), .A2(G472), .ZN(n356) );
  XOR2_X1 U466 ( .A(KEYINPUT56), .B(KEYINPUT124), .Z(n357) );
  AND2_X1 U467 ( .A1(n605), .A2(G953), .ZN(n711) );
  INV_X1 U468 ( .A(n711), .ZN(n382) );
  NOR2_X1 U469 ( .A1(n538), .A2(n624), .ZN(n543) );
  XNOR2_X2 U470 ( .A(n349), .B(n426), .ZN(n538) );
  NAND2_X1 U471 ( .A1(n529), .A2(n358), .ZN(n378) );
  AND2_X1 U472 ( .A1(n358), .A2(n385), .ZN(n533) );
  NAND2_X1 U473 ( .A1(n345), .A2(n362), .ZN(n365) );
  NAND2_X1 U474 ( .A1(n665), .A2(KEYINPUT122), .ZN(n359) );
  NAND2_X1 U475 ( .A1(n664), .A2(KEYINPUT122), .ZN(n361) );
  NAND2_X1 U476 ( .A1(n364), .A2(n363), .ZN(n362) );
  INV_X1 U477 ( .A(n665), .ZN(n364) );
  XNOR2_X1 U478 ( .A(n365), .B(n666), .ZN(G75) );
  NAND2_X1 U479 ( .A1(n378), .A2(n347), .ZN(n374) );
  NOR2_X1 U480 ( .A1(n532), .A2(KEYINPUT80), .ZN(n376) );
  NAND2_X1 U481 ( .A1(n694), .A2(n676), .ZN(n503) );
  XNOR2_X2 U482 ( .A(n380), .B(n379), .ZN(n694) );
  NAND2_X1 U483 ( .A1(n636), .A2(n509), .ZN(n380) );
  XNOR2_X1 U484 ( .A(n381), .B(n357), .ZN(G51) );
  XNOR2_X1 U485 ( .A(n385), .B(G122), .ZN(G24) );
  NAND2_X1 U486 ( .A1(n630), .A2(KEYINPUT100), .ZN(n387) );
  NAND2_X1 U487 ( .A1(n390), .A2(n389), .ZN(n388) );
  NAND2_X1 U488 ( .A1(n511), .A2(KEYINPUT100), .ZN(n389) );
  NAND2_X1 U489 ( .A1(n392), .A2(n394), .ZN(n391) );
  XNOR2_X2 U490 ( .A(n498), .B(KEYINPUT1), .ZN(n511) );
  NAND2_X1 U491 ( .A1(n701), .A2(n395), .ZN(n709) );
  NAND2_X1 U492 ( .A1(n701), .A2(n356), .ZN(n669) );
  NAND2_X1 U493 ( .A1(n346), .A2(G478), .ZN(n706) );
  NAND2_X1 U494 ( .A1(n346), .A2(G469), .ZN(n612) );
  XNOR2_X1 U495 ( .A(n451), .B(n351), .ZN(n397) );
  BUF_X1 U496 ( .A(n511), .Z(n631) );
  XNOR2_X1 U497 ( .A(n461), .B(n350), .ZN(n574) );
  NOR2_X2 U498 ( .A1(n734), .A2(n588), .ZN(n589) );
  XNOR2_X1 U499 ( .A(n504), .B(KEYINPUT98), .ZN(n517) );
  BUF_X1 U500 ( .A(n498), .Z(n567) );
  BUF_X1 U501 ( .A(n653), .Z(n660) );
  NOR2_X2 U502 ( .A1(n517), .A2(n674), .ZN(n531) );
  NAND2_X1 U503 ( .A1(n574), .A2(n467), .ZN(n469) );
  XNOR2_X2 U504 ( .A(n535), .B(KEYINPUT45), .ZN(n714) );
  XNOR2_X1 U505 ( .A(KEYINPUT64), .B(KEYINPUT46), .ZN(n572) );
  XNOR2_X1 U506 ( .A(n573), .B(n572), .ZN(n587) );
  XNOR2_X1 U507 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U508 ( .A(n456), .ZN(n457) );
  XNOR2_X1 U509 ( .A(n448), .B(n439), .ZN(n440) );
  XNOR2_X1 U510 ( .A(n446), .B(n445), .ZN(n653) );
  XNOR2_X1 U511 ( .A(n441), .B(n440), .ZN(n667) );
  XNOR2_X1 U512 ( .A(n483), .B(G478), .ZN(n484) );
  XNOR2_X1 U513 ( .A(n521), .B(KEYINPUT75), .ZN(n522) );
  XNOR2_X2 U514 ( .A(KEYINPUT65), .B(G143), .ZN(n401) );
  XNOR2_X2 U515 ( .A(n401), .B(n400), .ZN(n451) );
  XNOR2_X2 U516 ( .A(n451), .B(G134), .ZN(n481) );
  XNOR2_X1 U517 ( .A(n486), .B(n403), .ZN(n404) );
  NAND2_X1 U518 ( .A1(n730), .A2(G227), .ZN(n405) );
  XNOR2_X1 U519 ( .A(n406), .B(n405), .ZN(n408) );
  XNOR2_X1 U520 ( .A(G146), .B(G140), .ZN(n407) );
  XNOR2_X1 U521 ( .A(n408), .B(n407), .ZN(n410) );
  XNOR2_X1 U522 ( .A(n409), .B(G104), .ZN(n447) );
  XNOR2_X1 U523 ( .A(n410), .B(n447), .ZN(n411) );
  XNOR2_X1 U524 ( .A(n724), .B(n411), .ZN(n610) );
  INV_X1 U525 ( .A(G469), .ZN(n412) );
  XNOR2_X2 U526 ( .A(n413), .B(n412), .ZN(n498) );
  XOR2_X1 U527 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n417) );
  INV_X1 U528 ( .A(KEYINPUT15), .ZN(n414) );
  XNOR2_X1 U529 ( .A(n414), .B(G902), .ZN(n700) );
  INV_X1 U530 ( .A(n700), .ZN(n600) );
  NAND2_X1 U531 ( .A1(G234), .A2(n600), .ZN(n415) );
  XNOR2_X1 U532 ( .A(KEYINPUT20), .B(n415), .ZN(n427) );
  NAND2_X1 U533 ( .A1(n427), .A2(G217), .ZN(n416) );
  XNOR2_X1 U534 ( .A(n417), .B(n416), .ZN(n426) );
  NAND2_X1 U535 ( .A1(G234), .A2(n730), .ZN(n418) );
  NAND2_X1 U536 ( .A1(G221), .A2(n476), .ZN(n423) );
  XNOR2_X1 U537 ( .A(n352), .B(n420), .ZN(n421) );
  XOR2_X2 U538 ( .A(G125), .B(G146), .Z(n455) );
  XNOR2_X1 U539 ( .A(n455), .B(KEYINPUT10), .ZN(n424) );
  XNOR2_X1 U540 ( .A(n424), .B(G140), .ZN(n722) );
  XNOR2_X1 U541 ( .A(n425), .B(n722), .ZN(n708) );
  NAND2_X1 U542 ( .A1(n427), .A2(G221), .ZN(n429) );
  INV_X1 U543 ( .A(KEYINPUT21), .ZN(n428) );
  XNOR2_X1 U544 ( .A(n429), .B(n428), .ZN(n537) );
  NAND2_X1 U545 ( .A1(n538), .A2(n537), .ZN(n630) );
  XNOR2_X1 U546 ( .A(n430), .B(G101), .ZN(n434) );
  XOR2_X1 U547 ( .A(KEYINPUT5), .B(KEYINPUT72), .Z(n436) );
  XNOR2_X1 U548 ( .A(G146), .B(KEYINPUT92), .ZN(n435) );
  XNOR2_X1 U549 ( .A(n436), .B(n435), .ZN(n438) );
  NOR2_X1 U550 ( .A1(G953), .A2(G237), .ZN(n490) );
  NAND2_X1 U551 ( .A1(G210), .A2(n490), .ZN(n437) );
  XNOR2_X1 U552 ( .A(n438), .B(n437), .ZN(n439) );
  NOR2_X1 U553 ( .A1(G902), .A2(n667), .ZN(n443) );
  XOR2_X1 U554 ( .A(KEYINPUT93), .B(G472), .Z(n442) );
  INV_X1 U555 ( .A(KEYINPUT6), .ZN(n444) );
  XNOR2_X1 U556 ( .A(n563), .B(n444), .ZN(n544) );
  XOR2_X1 U557 ( .A(KEYINPUT71), .B(KEYINPUT16), .Z(n449) );
  XNOR2_X1 U558 ( .A(KEYINPUT18), .B(KEYINPUT4), .ZN(n452) );
  XNOR2_X1 U559 ( .A(n353), .B(n452), .ZN(n453) );
  NAND2_X1 U560 ( .A1(G224), .A2(n730), .ZN(n454) );
  OR2_X1 U561 ( .A1(G902), .A2(G237), .ZN(n460) );
  NAND2_X1 U562 ( .A1(G210), .A2(n460), .ZN(n458) );
  NAND2_X1 U563 ( .A1(G214), .A2(n460), .ZN(n641) );
  NAND2_X1 U564 ( .A1(n536), .A2(n641), .ZN(n461) );
  OR2_X1 U565 ( .A1(G898), .A2(n730), .ZN(n713) );
  NAND2_X1 U566 ( .A1(G234), .A2(G237), .ZN(n462) );
  XNOR2_X1 U567 ( .A(n462), .B(KEYINPUT14), .ZN(n464) );
  NAND2_X1 U568 ( .A1(G902), .A2(n464), .ZN(n539) );
  OR2_X1 U569 ( .A1(n713), .A2(n539), .ZN(n463) );
  XOR2_X1 U570 ( .A(KEYINPUT87), .B(n463), .Z(n466) );
  NAND2_X1 U571 ( .A1(n464), .A2(G952), .ZN(n658) );
  NOR2_X1 U572 ( .A1(G953), .A2(n658), .ZN(n465) );
  XOR2_X1 U573 ( .A(KEYINPUT86), .B(n465), .Z(n542) );
  NAND2_X1 U574 ( .A1(n466), .A2(n542), .ZN(n467) );
  XNOR2_X2 U575 ( .A(n469), .B(n468), .ZN(n509) );
  NAND2_X1 U576 ( .A1(n653), .A2(n509), .ZN(n472) );
  INV_X1 U577 ( .A(KEYINPUT70), .ZN(n470) );
  XNOR2_X1 U578 ( .A(n470), .B(KEYINPUT34), .ZN(n471) );
  XNOR2_X1 U579 ( .A(n472), .B(n471), .ZN(n493) );
  XOR2_X1 U580 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n474) );
  XNOR2_X1 U581 ( .A(G116), .B(KEYINPUT95), .ZN(n473) );
  XNOR2_X1 U582 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U583 ( .A(n475), .B(KEYINPUT96), .Z(n480) );
  NAND2_X1 U584 ( .A1(n476), .A2(G217), .ZN(n478) );
  XNOR2_X1 U585 ( .A(n478), .B(n477), .ZN(n479) );
  XNOR2_X1 U586 ( .A(n480), .B(n479), .ZN(n482) );
  XNOR2_X1 U587 ( .A(n482), .B(n481), .ZN(n705) );
  NOR2_X1 U588 ( .A1(G902), .A2(n705), .ZN(n485) );
  XOR2_X1 U589 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n489) );
  NAND2_X1 U590 ( .A1(n490), .A2(G214), .ZN(n491) );
  NOR2_X1 U591 ( .A1(n505), .A2(n506), .ZN(n579) );
  NAND2_X1 U592 ( .A1(n493), .A2(n579), .ZN(n496) );
  INV_X1 U593 ( .A(KEYINPUT78), .ZN(n494) );
  XNOR2_X1 U594 ( .A(n494), .B(KEYINPUT35), .ZN(n495) );
  NOR2_X1 U595 ( .A1(n567), .A2(n630), .ZN(n499) );
  NAND2_X1 U596 ( .A1(n509), .A2(n499), .ZN(n500) );
  XNOR2_X1 U597 ( .A(n500), .B(KEYINPUT91), .ZN(n501) );
  NAND2_X1 U598 ( .A1(n501), .A2(n563), .ZN(n676) );
  NAND2_X1 U599 ( .A1(n505), .A2(n502), .ZN(n691) );
  NOR2_X1 U600 ( .A1(n505), .A2(n502), .ZN(n683) );
  INV_X1 U601 ( .A(n683), .ZN(n695) );
  NAND2_X1 U602 ( .A1(n691), .A2(n695), .ZN(n647) );
  AND2_X1 U603 ( .A1(n503), .A2(n647), .ZN(n504) );
  AND2_X1 U604 ( .A1(n507), .A2(n537), .ZN(n508) );
  NAND2_X1 U605 ( .A1(n509), .A2(n508), .ZN(n510) );
  NAND2_X1 U606 ( .A1(n544), .A2(n631), .ZN(n512) );
  INV_X1 U607 ( .A(KEYINPUT79), .ZN(n513) );
  XNOR2_X1 U608 ( .A(n514), .B(n513), .ZN(n516) );
  XNOR2_X1 U609 ( .A(n538), .B(KEYINPUT99), .ZN(n623) );
  INV_X1 U610 ( .A(n623), .ZN(n515) );
  AND2_X1 U611 ( .A1(n516), .A2(n515), .ZN(n674) );
  INV_X1 U612 ( .A(n518), .ZN(n524) );
  NAND2_X1 U613 ( .A1(n544), .A2(n623), .ZN(n519) );
  NOR2_X1 U614 ( .A1(n519), .A2(n631), .ZN(n520) );
  XOR2_X1 U615 ( .A(KEYINPUT32), .B(KEYINPUT66), .Z(n521) );
  INV_X1 U616 ( .A(n538), .ZN(n525) );
  AND2_X1 U617 ( .A1(n563), .A2(n525), .ZN(n526) );
  AND2_X1 U618 ( .A1(n631), .A2(n526), .ZN(n527) );
  NAND2_X1 U619 ( .A1(n524), .A2(n527), .ZN(n682) );
  NAND2_X1 U620 ( .A1(n736), .A2(n682), .ZN(n528) );
  INV_X1 U621 ( .A(KEYINPUT44), .ZN(n530) );
  NAND2_X1 U622 ( .A1(n531), .A2(n530), .ZN(n532) );
  NAND2_X1 U623 ( .A1(n533), .A2(n530), .ZN(n534) );
  INV_X1 U624 ( .A(n551), .ZN(n593) );
  INV_X1 U625 ( .A(n537), .ZN(n624) );
  NOR2_X1 U626 ( .A1(G900), .A2(n539), .ZN(n540) );
  NAND2_X1 U627 ( .A1(G953), .A2(n540), .ZN(n541) );
  NAND2_X1 U628 ( .A1(n542), .A2(n541), .ZN(n552) );
  NAND2_X1 U629 ( .A1(n543), .A2(n552), .ZN(n564) );
  NOR2_X1 U630 ( .A1(n544), .A2(n564), .ZN(n545) );
  XNOR2_X1 U631 ( .A(n545), .B(KEYINPUT101), .ZN(n546) );
  NOR2_X1 U632 ( .A1(n691), .A2(n546), .ZN(n547) );
  NAND2_X1 U633 ( .A1(n547), .A2(n641), .ZN(n590) );
  XOR2_X1 U634 ( .A(KEYINPUT36), .B(n548), .Z(n549) );
  NOR2_X1 U635 ( .A1(n549), .A2(n631), .ZN(n550) );
  XOR2_X1 U636 ( .A(KEYINPUT107), .B(n550), .Z(n734) );
  INV_X1 U637 ( .A(n691), .ZN(n688) );
  NAND2_X1 U638 ( .A1(n392), .A2(n552), .ZN(n553) );
  NOR2_X1 U639 ( .A1(n567), .A2(n553), .ZN(n557) );
  INV_X1 U640 ( .A(n563), .ZN(n628) );
  NAND2_X1 U641 ( .A1(n641), .A2(n628), .ZN(n555) );
  NAND2_X1 U642 ( .A1(n557), .A2(n556), .ZN(n577) );
  INV_X1 U643 ( .A(n577), .ZN(n558) );
  NAND2_X1 U644 ( .A1(n642), .A2(n558), .ZN(n559) );
  XNOR2_X1 U645 ( .A(KEYINPUT39), .B(n559), .ZN(n595) );
  AND2_X1 U646 ( .A1(n688), .A2(n595), .ZN(n560) );
  XNOR2_X1 U647 ( .A(KEYINPUT40), .B(n560), .ZN(n737) );
  NAND2_X1 U648 ( .A1(n642), .A2(n641), .ZN(n648) );
  XOR2_X1 U649 ( .A(KEYINPUT41), .B(KEYINPUT106), .Z(n561) );
  XNOR2_X1 U650 ( .A(n562), .B(n561), .ZN(n661) );
  INV_X1 U651 ( .A(n661), .ZN(n570) );
  XNOR2_X1 U652 ( .A(n565), .B(KEYINPUT28), .ZN(n566) );
  XNOR2_X1 U653 ( .A(KEYINPUT105), .B(n566), .ZN(n569) );
  INV_X1 U654 ( .A(n567), .ZN(n568) );
  NAND2_X1 U655 ( .A1(n569), .A2(n568), .ZN(n576) );
  NOR2_X1 U656 ( .A1(n570), .A2(n576), .ZN(n571) );
  XNOR2_X1 U657 ( .A(n571), .B(KEYINPUT42), .ZN(n738) );
  INV_X1 U658 ( .A(n574), .ZN(n575) );
  NAND2_X1 U659 ( .A1(n689), .A2(n647), .ZN(n583) );
  NAND2_X1 U660 ( .A1(n583), .A2(KEYINPUT47), .ZN(n581) );
  NOR2_X1 U661 ( .A1(n593), .A2(n577), .ZN(n578) );
  XNOR2_X1 U662 ( .A(KEYINPUT104), .B(n578), .ZN(n580) );
  NAND2_X1 U663 ( .A1(n580), .A2(n579), .ZN(n687) );
  NAND2_X1 U664 ( .A1(n581), .A2(n687), .ZN(n582) );
  XNOR2_X1 U665 ( .A(n582), .B(KEYINPUT76), .ZN(n585) );
  NOR2_X1 U666 ( .A1(KEYINPUT47), .A2(n583), .ZN(n584) );
  NAND2_X1 U667 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U668 ( .A(n589), .B(KEYINPUT48), .ZN(n598) );
  XOR2_X1 U669 ( .A(KEYINPUT102), .B(n590), .Z(n591) );
  NAND2_X1 U670 ( .A1(n591), .A2(n631), .ZN(n592) );
  XNOR2_X1 U671 ( .A(n592), .B(KEYINPUT43), .ZN(n594) );
  AND2_X1 U672 ( .A1(n594), .A2(n593), .ZN(n698) );
  NAND2_X1 U673 ( .A1(n683), .A2(n595), .ZN(n697) );
  INV_X1 U674 ( .A(n697), .ZN(n596) );
  NOR2_X1 U675 ( .A1(n698), .A2(n596), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n714), .A2(n728), .ZN(n617) );
  INV_X1 U677 ( .A(KEYINPUT2), .ZN(n615) );
  XNOR2_X1 U678 ( .A(n617), .B(n615), .ZN(n599) );
  INV_X2 U679 ( .A(n599), .ZN(n701) );
  XOR2_X1 U680 ( .A(KEYINPUT67), .B(KEYINPUT59), .Z(n601) );
  XNOR2_X1 U681 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U682 ( .A(n604), .B(n603), .ZN(n606) );
  INV_X1 U683 ( .A(G952), .ZN(n605) );
  NAND2_X1 U684 ( .A1(n606), .A2(n382), .ZN(n608) );
  INV_X1 U685 ( .A(KEYINPUT60), .ZN(n607) );
  XNOR2_X1 U686 ( .A(n608), .B(n607), .ZN(G60) );
  XOR2_X1 U687 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n609) );
  XNOR2_X1 U688 ( .A(n610), .B(n609), .ZN(n611) );
  XNOR2_X1 U689 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X1 U690 ( .A1(n613), .A2(n711), .ZN(G54) );
  XNOR2_X1 U691 ( .A(n714), .B(KEYINPUT77), .ZN(n614) );
  NOR2_X1 U692 ( .A1(n614), .A2(KEYINPUT2), .ZN(n619) );
  NOR2_X1 U693 ( .A1(n615), .A2(KEYINPUT77), .ZN(n616) );
  AND2_X1 U694 ( .A1(n617), .A2(n616), .ZN(n618) );
  NOR2_X1 U695 ( .A1(n619), .A2(n618), .ZN(n621) );
  NOR2_X1 U696 ( .A1(n728), .A2(KEYINPUT2), .ZN(n620) );
  NOR2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n665) );
  XOR2_X1 U698 ( .A(KEYINPUT114), .B(KEYINPUT49), .Z(n622) );
  XNOR2_X1 U699 ( .A(KEYINPUT115), .B(n622), .ZN(n626) );
  AND2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n625) );
  XOR2_X1 U701 ( .A(n626), .B(n625), .Z(n627) );
  NOR2_X1 U702 ( .A1(n628), .A2(n627), .ZN(n629) );
  XOR2_X1 U703 ( .A(KEYINPUT116), .B(n629), .Z(n634) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT50), .B(n632), .Z(n633) );
  NOR2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n635) );
  XOR2_X1 U707 ( .A(KEYINPUT117), .B(n635), .Z(n637) );
  NOR2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n638) );
  XNOR2_X1 U709 ( .A(KEYINPUT118), .B(n638), .ZN(n639) );
  XNOR2_X1 U710 ( .A(n639), .B(KEYINPUT51), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n640), .A2(n661), .ZN(n656) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U713 ( .A(KEYINPUT119), .B(n643), .Z(n644) );
  NOR2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U715 ( .A(KEYINPUT120), .B(n646), .ZN(n651) );
  INV_X1 U716 ( .A(n647), .ZN(n649) );
  NOR2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n652), .B(KEYINPUT121), .ZN(n654) );
  NAND2_X1 U720 ( .A1(n654), .A2(n660), .ZN(n655) );
  NAND2_X1 U721 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U722 ( .A(n657), .B(KEYINPUT52), .Z(n659) );
  OR2_X1 U723 ( .A1(n659), .A2(n658), .ZN(n663) );
  NAND2_X1 U724 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U725 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U726 ( .A(KEYINPUT123), .B(KEYINPUT53), .ZN(n666) );
  XNOR2_X1 U727 ( .A(n667), .B(KEYINPUT62), .ZN(n668) );
  XNOR2_X1 U728 ( .A(n669), .B(n668), .ZN(n670) );
  NOR2_X2 U729 ( .A1(n670), .A2(n711), .ZN(n673) );
  XOR2_X1 U730 ( .A(KEYINPUT82), .B(KEYINPUT108), .Z(n671) );
  XNOR2_X1 U731 ( .A(KEYINPUT63), .B(n671), .ZN(n672) );
  XNOR2_X1 U732 ( .A(n673), .B(n672), .ZN(G57) );
  XOR2_X1 U733 ( .A(G101), .B(n674), .Z(G3) );
  NOR2_X1 U734 ( .A1(n691), .A2(n676), .ZN(n675) );
  XOR2_X1 U735 ( .A(G104), .B(n675), .Z(G6) );
  NOR2_X1 U736 ( .A1(n695), .A2(n676), .ZN(n681) );
  XOR2_X1 U737 ( .A(KEYINPUT110), .B(KEYINPUT27), .Z(n678) );
  XNOR2_X1 U738 ( .A(G107), .B(KEYINPUT26), .ZN(n677) );
  XNOR2_X1 U739 ( .A(n678), .B(n677), .ZN(n679) );
  XNOR2_X1 U740 ( .A(KEYINPUT109), .B(n679), .ZN(n680) );
  XNOR2_X1 U741 ( .A(n681), .B(n680), .ZN(G9) );
  XNOR2_X1 U742 ( .A(G110), .B(n682), .ZN(G12) );
  XOR2_X1 U743 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U744 ( .A1(n689), .A2(n683), .ZN(n684) );
  XNOR2_X1 U745 ( .A(n685), .B(n684), .ZN(G30) );
  XOR2_X1 U746 ( .A(G143), .B(KEYINPUT111), .Z(n686) );
  XNOR2_X1 U747 ( .A(n687), .B(n686), .ZN(G45) );
  NAND2_X1 U748 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U749 ( .A(n690), .B(G146), .ZN(G48) );
  NOR2_X1 U750 ( .A1(n691), .A2(n694), .ZN(n692) );
  XOR2_X1 U751 ( .A(KEYINPUT112), .B(n692), .Z(n693) );
  XNOR2_X1 U752 ( .A(G113), .B(n693), .ZN(G15) );
  NOR2_X1 U753 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U754 ( .A(G116), .B(n696), .Z(G18) );
  XNOR2_X1 U755 ( .A(G134), .B(n697), .ZN(G36) );
  XNOR2_X1 U756 ( .A(G140), .B(n698), .ZN(n699) );
  XNOR2_X1 U757 ( .A(n699), .B(KEYINPUT113), .ZN(G42) );
  AND2_X1 U758 ( .A1(G210), .A2(n700), .ZN(n702) );
  XOR2_X1 U759 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n703) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n711), .A2(n707), .ZN(G63) );
  XNOR2_X1 U762 ( .A(n709), .B(n708), .ZN(n710) );
  NOR2_X1 U763 ( .A1(n711), .A2(n710), .ZN(G66) );
  NAND2_X1 U764 ( .A1(n713), .A2(n712), .ZN(n721) );
  NAND2_X1 U765 ( .A1(n714), .A2(n730), .ZN(n719) );
  NAND2_X1 U766 ( .A1(G953), .A2(G224), .ZN(n715) );
  XNOR2_X1 U767 ( .A(KEYINPUT61), .B(n715), .ZN(n716) );
  NAND2_X1 U768 ( .A1(n716), .A2(G898), .ZN(n717) );
  XOR2_X1 U769 ( .A(KEYINPUT125), .B(n717), .Z(n718) );
  NAND2_X1 U770 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U771 ( .A(n721), .B(n720), .Z(G69) );
  XOR2_X1 U772 ( .A(KEYINPUT126), .B(n722), .Z(n723) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(n729) );
  XNOR2_X1 U774 ( .A(KEYINPUT127), .B(n729), .ZN(n725) );
  XNOR2_X1 U775 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U776 ( .A1(n726), .A2(G900), .ZN(n727) );
  NAND2_X1 U777 ( .A1(n727), .A2(G953), .ZN(n733) );
  XNOR2_X1 U778 ( .A(n729), .B(n728), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n733), .A2(n732), .ZN(G72) );
  XNOR2_X1 U781 ( .A(G125), .B(n734), .ZN(n735) );
  XNOR2_X1 U782 ( .A(n735), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U783 ( .A(n736), .B(G119), .ZN(G21) );
  XOR2_X1 U784 ( .A(G131), .B(n737), .Z(G33) );
  XOR2_X1 U785 ( .A(G137), .B(n738), .Z(G39) );
endmodule

