

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723;

  NOR2_X1 U364 ( .A1(n656), .A2(n657), .ZN(n661) );
  INV_X2 U365 ( .A(G953), .ZN(n699) );
  NOR2_X1 U366 ( .A1(G953), .A2(G237), .ZN(n402) );
  XNOR2_X1 U367 ( .A(n426), .B(n425), .ZN(n698) );
  XNOR2_X1 U368 ( .A(n480), .B(KEYINPUT35), .ZN(n721) );
  AND2_X2 U369 ( .A1(n492), .A2(n575), .ZN(n496) );
  XNOR2_X2 U370 ( .A(n477), .B(n476), .ZN(n507) );
  NAND2_X1 U371 ( .A1(n354), .A2(n352), .ZN(n707) );
  NAND2_X1 U372 ( .A1(n661), .A2(n658), .ZN(n523) );
  XNOR2_X1 U373 ( .A(n541), .B(n441), .ZN(n556) );
  XNOR2_X1 U374 ( .A(n493), .B(KEYINPUT100), .ZN(n413) );
  INV_X2 U375 ( .A(G143), .ZN(n375) );
  NOR2_X1 U376 ( .A1(n610), .A2(n691), .ZN(n611) );
  NOR2_X1 U377 ( .A1(n593), .A2(n691), .ZN(n595) );
  NOR2_X1 U378 ( .A1(n603), .A2(n691), .ZN(n605) );
  NOR2_X1 U379 ( .A1(n617), .A2(n691), .ZN(n619) );
  XNOR2_X2 U380 ( .A(n548), .B(n518), .ZN(n657) );
  XNOR2_X2 U381 ( .A(n705), .B(G146), .ZN(n409) );
  XNOR2_X2 U382 ( .A(n423), .B(n351), .ZN(n705) );
  XNOR2_X2 U383 ( .A(n450), .B(n376), .ZN(n423) );
  NAND2_X1 U384 ( .A1(n363), .A2(n519), .ZN(n360) );
  XNOR2_X1 U385 ( .A(n488), .B(n487), .ZN(n492) );
  NAND2_X1 U386 ( .A1(n503), .A2(n343), .ZN(n488) );
  XOR2_X1 U387 ( .A(G140), .B(G113), .Z(n460) );
  XNOR2_X1 U388 ( .A(KEYINPUT88), .B(KEYINPUT48), .ZN(n570) );
  XOR2_X1 U389 ( .A(KEYINPUT10), .B(n420), .Z(n466) );
  XNOR2_X1 U390 ( .A(n377), .B(G131), .ZN(n351) );
  NOR2_X1 U391 ( .A1(n494), .A2(n598), .ZN(n495) );
  OR2_X1 U392 ( .A1(n649), .A2(n341), .ZN(n363) );
  NAND2_X1 U393 ( .A1(n361), .A2(n344), .ZN(n359) );
  XNOR2_X1 U394 ( .A(n466), .B(n393), .ZN(n704) );
  INV_X1 U395 ( .A(n392), .ZN(n393) );
  XNOR2_X1 U396 ( .A(n371), .B(KEYINPUT23), .ZN(n370) );
  INV_X1 U397 ( .A(KEYINPUT70), .ZN(n371) );
  XNOR2_X1 U398 ( .A(n475), .B(n474), .ZN(n476) );
  INV_X1 U399 ( .A(G475), .ZN(n474) );
  NAND2_X1 U400 ( .A1(n367), .A2(n347), .ZN(n366) );
  XNOR2_X1 U401 ( .A(n416), .B(n417), .ZN(n373) );
  INV_X1 U402 ( .A(KEYINPUT33), .ZN(n417) );
  INV_X1 U403 ( .A(G902), .ZN(n443) );
  INV_X1 U404 ( .A(G101), .ZN(n405) );
  XNOR2_X1 U405 ( .A(G137), .B(G116), .ZN(n406) );
  XNOR2_X1 U406 ( .A(n403), .B(G113), .ZN(n425) );
  XNOR2_X1 U407 ( .A(KEYINPUT3), .B(G119), .ZN(n403) );
  XNOR2_X1 U408 ( .A(n424), .B(G116), .ZN(n449) );
  XNOR2_X1 U409 ( .A(G104), .B(G122), .ZN(n467) );
  XNOR2_X1 U410 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U411 ( .A(G146), .ZN(n391) );
  XNOR2_X1 U412 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n419) );
  NOR2_X1 U413 ( .A1(n527), .A2(n526), .ZN(n538) );
  XNOR2_X1 U414 ( .A(n401), .B(KEYINPUT66), .ZN(n501) );
  NOR2_X1 U415 ( .A1(n481), .A2(n644), .ZN(n401) );
  XNOR2_X1 U416 ( .A(n409), .B(n348), .ZN(n589) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n348) );
  XNOR2_X1 U418 ( .A(n407), .B(n404), .ZN(n349) );
  XNOR2_X1 U419 ( .A(n408), .B(n425), .ZN(n350) );
  AND2_X1 U420 ( .A1(n597), .A2(n353), .ZN(n352) );
  XNOR2_X1 U421 ( .A(n355), .B(n570), .ZN(n354) );
  INV_X1 U422 ( .A(n642), .ZN(n353) );
  XNOR2_X1 U423 ( .A(G104), .B(G107), .ZN(n378) );
  XOR2_X1 U424 ( .A(G107), .B(G134), .Z(n455) );
  XNOR2_X1 U425 ( .A(n513), .B(KEYINPUT45), .ZN(n692) );
  XNOR2_X1 U426 ( .A(n522), .B(n521), .ZN(n571) );
  INV_X1 U427 ( .A(KEYINPUT39), .ZN(n521) );
  NOR2_X1 U428 ( .A1(n360), .A2(n359), .ZN(n520) );
  INV_X1 U429 ( .A(n359), .ZN(n358) );
  XNOR2_X1 U430 ( .A(n506), .B(n505), .ZN(n537) );
  INV_X1 U431 ( .A(KEYINPUT99), .ZN(n505) );
  XNOR2_X1 U432 ( .A(n390), .B(n369), .ZN(n368) );
  XNOR2_X1 U433 ( .A(n388), .B(n370), .ZN(n369) );
  AND2_X1 U434 ( .A1(n592), .A2(G953), .ZN(n691) );
  XNOR2_X1 U435 ( .A(n357), .B(n356), .ZN(n718) );
  XNOR2_X1 U436 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n356) );
  NOR2_X1 U437 ( .A1(n571), .A2(n537), .ZN(n357) );
  AND2_X1 U438 ( .A1(n479), .A2(n551), .ZN(n480) );
  AND2_X1 U439 ( .A1(n364), .A2(n345), .ZN(n598) );
  XNOR2_X1 U440 ( .A(n496), .B(n365), .ZN(n364) );
  INV_X1 U441 ( .A(KEYINPUT101), .ZN(n365) );
  OR2_X1 U442 ( .A1(n656), .A2(KEYINPUT30), .ZN(n341) );
  NOR2_X1 U443 ( .A1(n649), .A2(n499), .ZN(n342) );
  AND2_X1 U444 ( .A1(n658), .A2(n485), .ZN(n343) );
  AND2_X1 U445 ( .A1(n362), .A2(n517), .ZN(n344) );
  AND2_X1 U446 ( .A1(n643), .A2(n649), .ZN(n345) );
  AND2_X1 U447 ( .A1(n358), .A2(n363), .ZN(n346) );
  AND2_X1 U448 ( .A1(n516), .A2(n447), .ZN(n347) );
  XNOR2_X1 U449 ( .A(n704), .B(n368), .ZN(n686) );
  XNOR2_X2 U450 ( .A(n412), .B(n411), .ZN(n493) );
  XOR2_X2 U451 ( .A(KEYINPUT83), .B(n558), .Z(n633) );
  AND2_X2 U452 ( .A1(n569), .A2(n568), .ZN(n355) );
  NAND2_X1 U453 ( .A1(n649), .A2(KEYINPUT30), .ZN(n361) );
  NAND2_X1 U454 ( .A1(n656), .A2(KEYINPUT30), .ZN(n362) );
  XNOR2_X2 U455 ( .A(n366), .B(n448), .ZN(n503) );
  INV_X1 U456 ( .A(n556), .ZN(n367) );
  XNOR2_X1 U457 ( .A(n372), .B(n374), .ZN(n479) );
  NAND2_X1 U458 ( .A1(n675), .A2(n503), .ZN(n372) );
  XNOR2_X2 U459 ( .A(n415), .B(n373), .ZN(n675) );
  BUF_X1 U460 ( .A(n681), .Z(n685) );
  XNOR2_X1 U461 ( .A(n429), .B(n428), .ZN(n614) );
  XNOR2_X1 U462 ( .A(KEYINPUT73), .B(KEYINPUT34), .ZN(n374) );
  XNOR2_X1 U463 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U464 ( .A(KEYINPUT107), .ZN(n529) );
  XNOR2_X1 U465 ( .A(n529), .B(KEYINPUT28), .ZN(n530) );
  XNOR2_X1 U466 ( .A(n427), .B(n698), .ZN(n428) );
  XNOR2_X1 U467 ( .A(n531), .B(n530), .ZN(n533) );
  XNOR2_X1 U468 ( .A(n686), .B(n687), .ZN(n688) );
  XNOR2_X1 U469 ( .A(n537), .B(KEYINPUT104), .ZN(n636) );
  INV_X1 U470 ( .A(KEYINPUT63), .ZN(n594) );
  XNOR2_X1 U471 ( .A(n689), .B(n688), .ZN(n690) );
  XOR2_X1 U472 ( .A(KEYINPUT72), .B(KEYINPUT102), .Z(n416) );
  XNOR2_X2 U473 ( .A(n375), .B(G128), .ZN(n450) );
  INV_X1 U474 ( .A(KEYINPUT4), .ZN(n376) );
  XOR2_X1 U475 ( .A(G134), .B(KEYINPUT67), .Z(n377) );
  INV_X1 U476 ( .A(n378), .ZN(n380) );
  XNOR2_X1 U477 ( .A(G101), .B(G110), .ZN(n379) );
  XNOR2_X1 U478 ( .A(n380), .B(n379), .ZN(n697) );
  XNOR2_X1 U479 ( .A(n697), .B(KEYINPUT71), .ZN(n427) );
  XOR2_X1 U480 ( .A(G137), .B(G140), .Z(n392) );
  NAND2_X1 U481 ( .A1(G227), .A2(n699), .ZN(n381) );
  XNOR2_X1 U482 ( .A(n392), .B(n381), .ZN(n382) );
  XNOR2_X1 U483 ( .A(n427), .B(n382), .ZN(n383) );
  XNOR2_X1 U484 ( .A(n409), .B(n383), .ZN(n607) );
  OR2_X1 U485 ( .A1(n607), .A2(G902), .ZN(n385) );
  XNOR2_X1 U486 ( .A(KEYINPUT69), .B(G469), .ZN(n384) );
  XNOR2_X1 U487 ( .A(n385), .B(n384), .ZN(n502) );
  XNOR2_X1 U488 ( .A(n502), .B(KEYINPUT1), .ZN(n575) );
  INV_X1 U489 ( .A(n575), .ZN(n646) );
  XOR2_X1 U490 ( .A(KEYINPUT24), .B(G110), .Z(n387) );
  XNOR2_X1 U491 ( .A(G128), .B(G119), .ZN(n386) );
  XNOR2_X1 U492 ( .A(n387), .B(n386), .ZN(n388) );
  NAND2_X1 U493 ( .A1(n699), .A2(G234), .ZN(n389) );
  XOR2_X1 U494 ( .A(KEYINPUT8), .B(n389), .Z(n453) );
  NAND2_X1 U495 ( .A1(n453), .A2(G221), .ZN(n390) );
  XNOR2_X1 U496 ( .A(n391), .B(G125), .ZN(n420) );
  NOR2_X1 U497 ( .A1(n686), .A2(G902), .ZN(n397) );
  XNOR2_X2 U498 ( .A(KEYINPUT15), .B(G902), .ZN(n587) );
  NAND2_X1 U499 ( .A1(G234), .A2(n587), .ZN(n394) );
  XNOR2_X1 U500 ( .A(KEYINPUT20), .B(n394), .ZN(n398) );
  AND2_X1 U501 ( .A1(n398), .A2(G217), .ZN(n395) );
  XNOR2_X1 U502 ( .A(KEYINPUT25), .B(n395), .ZN(n396) );
  XNOR2_X1 U503 ( .A(n397), .B(n396), .ZN(n481) );
  AND2_X1 U504 ( .A1(n398), .A2(G221), .ZN(n400) );
  INV_X1 U505 ( .A(KEYINPUT21), .ZN(n399) );
  XNOR2_X1 U506 ( .A(n400), .B(n399), .ZN(n644) );
  NAND2_X1 U507 ( .A1(n646), .A2(n501), .ZN(n499) );
  INV_X1 U508 ( .A(KEYINPUT6), .ZN(n414) );
  XOR2_X1 U509 ( .A(KEYINPUT79), .B(n402), .Z(n469) );
  NAND2_X1 U510 ( .A1(n469), .A2(G210), .ZN(n408) );
  XNOR2_X1 U511 ( .A(KEYINPUT94), .B(KEYINPUT5), .ZN(n404) );
  NAND2_X1 U512 ( .A1(n589), .A2(n443), .ZN(n412) );
  INV_X1 U513 ( .A(KEYINPUT74), .ZN(n410) );
  XNOR2_X1 U514 ( .A(n410), .B(G472), .ZN(n411) );
  XNOR2_X2 U515 ( .A(n414), .B(n413), .ZN(n540) );
  OR2_X2 U516 ( .A1(n499), .A2(n540), .ZN(n415) );
  NAND2_X1 U517 ( .A1(n699), .A2(G224), .ZN(n418) );
  XNOR2_X1 U518 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U519 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U520 ( .A(n423), .B(n422), .ZN(n429) );
  INV_X1 U521 ( .A(G122), .ZN(n424) );
  XNOR2_X1 U522 ( .A(n449), .B(KEYINPUT16), .ZN(n426) );
  INV_X1 U523 ( .A(n587), .ZN(n430) );
  OR2_X2 U524 ( .A1(n614), .A2(n430), .ZN(n435) );
  INV_X1 U525 ( .A(G237), .ZN(n431) );
  NAND2_X1 U526 ( .A1(n443), .A2(n431), .ZN(n436) );
  NAND2_X1 U527 ( .A1(n436), .A2(G210), .ZN(n433) );
  INV_X1 U528 ( .A(KEYINPUT92), .ZN(n432) );
  XNOR2_X1 U529 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X2 U530 ( .A(n435), .B(n434), .ZN(n548) );
  NAND2_X1 U531 ( .A1(n436), .A2(G214), .ZN(n437) );
  XNOR2_X1 U532 ( .A(n437), .B(KEYINPUT93), .ZN(n656) );
  INV_X1 U533 ( .A(n656), .ZN(n438) );
  NAND2_X1 U534 ( .A1(n548), .A2(n438), .ZN(n541) );
  XNOR2_X1 U535 ( .A(KEYINPUT80), .B(KEYINPUT19), .ZN(n440) );
  INV_X1 U536 ( .A(KEYINPUT64), .ZN(n439) );
  XNOR2_X1 U537 ( .A(n440), .B(n439), .ZN(n441) );
  NAND2_X1 U538 ( .A1(G234), .A2(G237), .ZN(n442) );
  XNOR2_X1 U539 ( .A(n442), .B(KEYINPUT14), .ZN(n670) );
  INV_X1 U540 ( .A(G952), .ZN(n592) );
  NAND2_X1 U541 ( .A1(n699), .A2(n592), .ZN(n445) );
  NAND2_X1 U542 ( .A1(G953), .A2(n443), .ZN(n444) );
  AND2_X1 U543 ( .A1(n445), .A2(n444), .ZN(n446) );
  AND2_X1 U544 ( .A1(n670), .A2(n446), .ZN(n516) );
  NAND2_X1 U545 ( .A1(G953), .A2(G898), .ZN(n447) );
  INV_X1 U546 ( .A(KEYINPUT0), .ZN(n448) );
  XOR2_X1 U547 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n452) );
  XNOR2_X1 U548 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U549 ( .A(n452), .B(n451), .ZN(n457) );
  NAND2_X1 U550 ( .A1(G217), .A2(n453), .ZN(n454) );
  XNOR2_X1 U551 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U552 ( .A(n457), .B(n456), .ZN(n682) );
  NOR2_X1 U553 ( .A1(G902), .A2(n682), .ZN(n458) );
  XNOR2_X1 U554 ( .A(G478), .B(n458), .ZN(n508) );
  INV_X1 U555 ( .A(n508), .ZN(n484) );
  XNOR2_X1 U556 ( .A(G143), .B(G131), .ZN(n459) );
  XNOR2_X1 U557 ( .A(n460), .B(n459), .ZN(n464) );
  XOR2_X1 U558 ( .A(KEYINPUT95), .B(KEYINPUT12), .Z(n462) );
  XNOR2_X1 U559 ( .A(KEYINPUT98), .B(KEYINPUT96), .ZN(n461) );
  XNOR2_X1 U560 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U561 ( .A(n466), .B(n465), .ZN(n473) );
  XOR2_X1 U562 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n468) );
  XNOR2_X1 U563 ( .A(n468), .B(n467), .ZN(n471) );
  NAND2_X1 U564 ( .A1(G214), .A2(n469), .ZN(n470) );
  XNOR2_X1 U565 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U566 ( .A(n473), .B(n472), .ZN(n600) );
  NOR2_X1 U567 ( .A1(G902), .A2(n600), .ZN(n477) );
  INV_X1 U568 ( .A(KEYINPUT13), .ZN(n475) );
  NAND2_X1 U569 ( .A1(n484), .A2(n507), .ZN(n478) );
  XNOR2_X1 U570 ( .A(n478), .B(KEYINPUT103), .ZN(n551) );
  INV_X1 U571 ( .A(n481), .ZN(n527) );
  INV_X1 U572 ( .A(n527), .ZN(n643) );
  NAND2_X1 U573 ( .A1(n540), .A2(n643), .ZN(n482) );
  XOR2_X1 U574 ( .A(KEYINPUT91), .B(n575), .Z(n544) );
  NOR2_X1 U575 ( .A1(n482), .A2(n544), .ZN(n483) );
  XNOR2_X1 U576 ( .A(n483), .B(KEYINPUT82), .ZN(n489) );
  NOR2_X1 U577 ( .A1(n507), .A2(n484), .ZN(n658) );
  INV_X1 U578 ( .A(n644), .ZN(n485) );
  XNOR2_X1 U579 ( .A(KEYINPUT76), .B(KEYINPUT22), .ZN(n486) );
  XNOR2_X1 U580 ( .A(n486), .B(KEYINPUT75), .ZN(n487) );
  NAND2_X1 U581 ( .A1(n489), .A2(n492), .ZN(n491) );
  XOR2_X1 U582 ( .A(KEYINPUT81), .B(KEYINPUT32), .Z(n490) );
  XNOR2_X1 U583 ( .A(n491), .B(n490), .ZN(n596) );
  NAND2_X1 U584 ( .A1(n721), .A2(n596), .ZN(n494) );
  BUF_X2 U585 ( .A(n493), .Z(n649) );
  XNOR2_X1 U586 ( .A(n495), .B(KEYINPUT44), .ZN(n512) );
  NAND2_X1 U587 ( .A1(n496), .A2(n540), .ZN(n497) );
  XNOR2_X1 U588 ( .A(n497), .B(KEYINPUT89), .ZN(n498) );
  NAND2_X1 U589 ( .A1(n498), .A2(n527), .ZN(n621) );
  NAND2_X1 U590 ( .A1(n503), .A2(n342), .ZN(n500) );
  XOR2_X1 U591 ( .A(KEYINPUT31), .B(n500), .Z(n638) );
  INV_X1 U592 ( .A(n502), .ZN(n532) );
  NAND2_X1 U593 ( .A1(n501), .A2(n532), .ZN(n514) );
  INV_X1 U594 ( .A(n649), .ZN(n528) );
  NOR2_X1 U595 ( .A1(n514), .A2(n528), .ZN(n504) );
  NAND2_X1 U596 ( .A1(n504), .A2(n503), .ZN(n625) );
  NAND2_X1 U597 ( .A1(n638), .A2(n625), .ZN(n509) );
  NAND2_X1 U598 ( .A1(n508), .A2(n507), .ZN(n506) );
  NOR2_X1 U599 ( .A1(n508), .A2(n507), .ZN(n628) );
  INV_X1 U600 ( .A(n628), .ZN(n639) );
  NAND2_X1 U601 ( .A1(n537), .A2(n639), .ZN(n660) );
  NAND2_X1 U602 ( .A1(n509), .A2(n660), .ZN(n510) );
  AND2_X1 U603 ( .A1(n621), .A2(n510), .ZN(n511) );
  NAND2_X1 U604 ( .A1(n512), .A2(n511), .ZN(n513) );
  XNOR2_X1 U605 ( .A(n514), .B(KEYINPUT105), .ZN(n547) );
  NAND2_X1 U606 ( .A1(G953), .A2(G900), .ZN(n515) );
  NAND2_X1 U607 ( .A1(n516), .A2(n515), .ZN(n524) );
  INV_X1 U608 ( .A(n524), .ZN(n517) );
  XNOR2_X1 U609 ( .A(KEYINPUT78), .B(KEYINPUT38), .ZN(n518) );
  INV_X1 U610 ( .A(n657), .ZN(n519) );
  NAND2_X1 U611 ( .A1(n547), .A2(n520), .ZN(n522) );
  XOR2_X1 U612 ( .A(KEYINPUT41), .B(n523), .Z(n654) );
  NOR2_X1 U613 ( .A1(n644), .A2(n524), .ZN(n525) );
  XOR2_X1 U614 ( .A(KEYINPUT68), .B(n525), .Z(n526) );
  AND2_X1 U615 ( .A1(n528), .A2(n538), .ZN(n531) );
  NAND2_X1 U616 ( .A1(n533), .A2(n532), .ZN(n557) );
  NOR2_X1 U617 ( .A1(n654), .A2(n557), .ZN(n534) );
  XOR2_X1 U618 ( .A(KEYINPUT109), .B(n534), .Z(n535) );
  XNOR2_X1 U619 ( .A(KEYINPUT42), .B(n535), .ZN(n720) );
  NOR2_X1 U620 ( .A1(n718), .A2(n720), .ZN(n536) );
  XNOR2_X1 U621 ( .A(KEYINPUT46), .B(n536), .ZN(n569) );
  INV_X1 U622 ( .A(n636), .ZN(n632) );
  NAND2_X1 U623 ( .A1(n538), .A2(n632), .ZN(n539) );
  NOR2_X2 U624 ( .A1(n540), .A2(n539), .ZN(n572) );
  INV_X1 U625 ( .A(n541), .ZN(n542) );
  NAND2_X1 U626 ( .A1(n572), .A2(n542), .ZN(n543) );
  XNOR2_X1 U627 ( .A(n543), .B(KEYINPUT36), .ZN(n545) );
  NOR2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U629 ( .A(n546), .B(KEYINPUT110), .ZN(n722) );
  INV_X1 U630 ( .A(n660), .ZN(n561) );
  NAND2_X1 U631 ( .A1(KEYINPUT47), .A2(n561), .ZN(n553) );
  NAND2_X1 U632 ( .A1(n547), .A2(n346), .ZN(n549) );
  INV_X1 U633 ( .A(n548), .ZN(n577) );
  NOR2_X1 U634 ( .A1(n549), .A2(n577), .ZN(n550) );
  XNOR2_X1 U635 ( .A(n550), .B(KEYINPUT106), .ZN(n552) );
  NAND2_X1 U636 ( .A1(n552), .A2(n551), .ZN(n631) );
  NAND2_X1 U637 ( .A1(n553), .A2(n631), .ZN(n554) );
  XNOR2_X1 U638 ( .A(n554), .B(KEYINPUT84), .ZN(n555) );
  NOR2_X1 U639 ( .A1(n722), .A2(n555), .ZN(n567) );
  NOR2_X2 U640 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U641 ( .A(KEYINPUT47), .ZN(n559) );
  NOR2_X1 U642 ( .A1(n633), .A2(n559), .ZN(n560) );
  XOR2_X1 U643 ( .A(n560), .B(KEYINPUT86), .Z(n565) );
  NOR2_X1 U644 ( .A1(KEYINPUT47), .A2(n561), .ZN(n562) );
  XOR2_X1 U645 ( .A(KEYINPUT77), .B(n562), .Z(n563) );
  NAND2_X1 U646 ( .A1(n633), .A2(n563), .ZN(n564) );
  AND2_X1 U647 ( .A1(n565), .A2(n564), .ZN(n566) );
  AND2_X1 U648 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U649 ( .A1(n639), .A2(n571), .ZN(n642) );
  INV_X1 U650 ( .A(n572), .ZN(n573) );
  NOR2_X1 U651 ( .A1(n656), .A2(n573), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U653 ( .A(KEYINPUT43), .B(n576), .ZN(n578) );
  NAND2_X1 U654 ( .A1(n578), .A2(n577), .ZN(n597) );
  INV_X1 U655 ( .A(n707), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n692), .A2(n582), .ZN(n579) );
  OR2_X1 U657 ( .A1(KEYINPUT2), .A2(KEYINPUT87), .ZN(n580) );
  NAND2_X1 U658 ( .A1(n579), .A2(n580), .ZN(n584) );
  INV_X1 U659 ( .A(n580), .ZN(n581) );
  NAND2_X1 U660 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U661 ( .A1(n584), .A2(n583), .ZN(n586) );
  OR2_X1 U662 ( .A1(n692), .A2(KEYINPUT2), .ZN(n585) );
  NAND2_X1 U663 ( .A1(n586), .A2(n585), .ZN(n679) );
  NOR2_X4 U664 ( .A1(n679), .A2(n587), .ZN(n681) );
  NAND2_X1 U665 ( .A1(n681), .A2(G472), .ZN(n591) );
  XOR2_X1 U666 ( .A(KEYINPUT90), .B(KEYINPUT62), .Z(n588) );
  XNOR2_X1 U667 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U668 ( .A(n591), .B(n590), .ZN(n593) );
  XNOR2_X1 U669 ( .A(n595), .B(n594), .ZN(G57) );
  XNOR2_X1 U670 ( .A(n596), .B(G119), .ZN(G21) );
  XNOR2_X1 U671 ( .A(n597), .B(G140), .ZN(G42) );
  XOR2_X1 U672 ( .A(n598), .B(G110), .Z(G12) );
  NAND2_X1 U673 ( .A1(n681), .A2(G475), .ZN(n602) );
  XNOR2_X1 U674 ( .A(KEYINPUT119), .B(KEYINPUT59), .ZN(n599) );
  XNOR2_X1 U675 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U676 ( .A(n602), .B(n601), .ZN(n603) );
  XOR2_X1 U677 ( .A(KEYINPUT65), .B(KEYINPUT60), .Z(n604) );
  XNOR2_X1 U678 ( .A(n605), .B(n604), .ZN(G60) );
  NAND2_X1 U679 ( .A1(n681), .A2(G469), .ZN(n609) );
  XOR2_X1 U680 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n606) );
  XNOR2_X1 U681 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n609), .B(n608), .ZN(n610) );
  XNOR2_X1 U683 ( .A(n611), .B(KEYINPUT118), .ZN(G54) );
  NAND2_X1 U684 ( .A1(n681), .A2(G210), .ZN(n616) );
  XNOR2_X1 U685 ( .A(KEYINPUT85), .B(KEYINPUT54), .ZN(n612) );
  XNOR2_X1 U686 ( .A(n612), .B(KEYINPUT55), .ZN(n613) );
  XNOR2_X1 U687 ( .A(n614), .B(n613), .ZN(n615) );
  XNOR2_X1 U688 ( .A(n616), .B(n615), .ZN(n617) );
  XOR2_X1 U689 ( .A(KEYINPUT117), .B(KEYINPUT56), .Z(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(G51) );
  XOR2_X1 U691 ( .A(G101), .B(KEYINPUT111), .Z(n620) );
  XNOR2_X1 U692 ( .A(n621), .B(n620), .ZN(G3) );
  NOR2_X1 U693 ( .A1(n636), .A2(n625), .ZN(n622) );
  XOR2_X1 U694 ( .A(G104), .B(n622), .Z(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT112), .B(KEYINPUT26), .Z(n624) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT27), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(n627) );
  NOR2_X1 U698 ( .A1(n639), .A2(n625), .ZN(n626) );
  XOR2_X1 U699 ( .A(n627), .B(n626), .Z(G9) );
  XOR2_X1 U700 ( .A(G128), .B(KEYINPUT29), .Z(n630) );
  NAND2_X1 U701 ( .A1(n633), .A2(n628), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n630), .B(n629), .ZN(G30) );
  XNOR2_X1 U703 ( .A(G143), .B(n631), .ZN(G45) );
  XOR2_X1 U704 ( .A(G146), .B(KEYINPUT113), .Z(n635) );
  NAND2_X1 U705 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(G48) );
  NOR2_X1 U707 ( .A1(n636), .A2(n638), .ZN(n637) );
  XOR2_X1 U708 ( .A(G113), .B(n637), .Z(G15) );
  NOR2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U710 ( .A(KEYINPUT114), .B(n640), .Z(n641) );
  XNOR2_X1 U711 ( .A(G116), .B(n641), .ZN(G18) );
  XOR2_X1 U712 ( .A(G134), .B(n642), .Z(G36) );
  NAND2_X1 U713 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U714 ( .A(n645), .B(KEYINPUT49), .ZN(n651) );
  NOR2_X1 U715 ( .A1(n646), .A2(n501), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT50), .B(n647), .Z(n648) );
  NAND2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  NOR2_X1 U718 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U719 ( .A1(n342), .A2(n652), .ZN(n653) );
  XNOR2_X1 U720 ( .A(n653), .B(KEYINPUT51), .ZN(n655) );
  INV_X1 U721 ( .A(n654), .ZN(n674) );
  NAND2_X1 U722 ( .A1(n655), .A2(n674), .ZN(n668) );
  NAND2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n659) );
  NAND2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n664) );
  NAND2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n662) );
  XOR2_X1 U726 ( .A(KEYINPUT115), .B(n662), .Z(n663) );
  NAND2_X1 U727 ( .A1(n664), .A2(n663), .ZN(n665) );
  XNOR2_X1 U728 ( .A(KEYINPUT116), .B(n665), .ZN(n666) );
  NAND2_X1 U729 ( .A1(n666), .A2(n675), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U731 ( .A(KEYINPUT52), .B(n669), .Z(n672) );
  NAND2_X1 U732 ( .A1(G952), .A2(n670), .ZN(n671) );
  NOR2_X1 U733 ( .A1(n672), .A2(n671), .ZN(n673) );
  OR2_X1 U734 ( .A1(G953), .A2(n673), .ZN(n677) );
  AND2_X1 U735 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U736 ( .A1(n677), .A2(n676), .ZN(n678) );
  AND2_X1 U737 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U738 ( .A(KEYINPUT53), .B(n680), .ZN(G75) );
  NAND2_X1 U739 ( .A1(n685), .A2(G478), .ZN(n683) );
  XNOR2_X1 U740 ( .A(n683), .B(n682), .ZN(n684) );
  NOR2_X1 U741 ( .A1(n691), .A2(n684), .ZN(G63) );
  NAND2_X1 U742 ( .A1(n685), .A2(G217), .ZN(n689) );
  XOR2_X1 U743 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n687) );
  NOR2_X1 U744 ( .A1(n691), .A2(n690), .ZN(G66) );
  NAND2_X1 U745 ( .A1(n692), .A2(n699), .ZN(n696) );
  NAND2_X1 U746 ( .A1(G953), .A2(G224), .ZN(n693) );
  XNOR2_X1 U747 ( .A(KEYINPUT61), .B(n693), .ZN(n694) );
  NAND2_X1 U748 ( .A1(n694), .A2(G898), .ZN(n695) );
  NAND2_X1 U749 ( .A1(n696), .A2(n695), .ZN(n703) );
  XNOR2_X1 U750 ( .A(n698), .B(n697), .ZN(n701) );
  NOR2_X1 U751 ( .A1(n699), .A2(G898), .ZN(n700) );
  NOR2_X1 U752 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U753 ( .A(n703), .B(n702), .ZN(G69) );
  XNOR2_X1 U754 ( .A(n705), .B(n704), .ZN(n706) );
  XOR2_X1 U755 ( .A(n706), .B(KEYINPUT122), .Z(n711) );
  XOR2_X1 U756 ( .A(n707), .B(KEYINPUT87), .Z(n708) );
  XOR2_X1 U757 ( .A(n711), .B(n708), .Z(n709) );
  NOR2_X1 U758 ( .A1(G953), .A2(n709), .ZN(n710) );
  XNOR2_X1 U759 ( .A(n710), .B(KEYINPUT123), .ZN(n717) );
  XNOR2_X1 U760 ( .A(KEYINPUT124), .B(n711), .ZN(n712) );
  XNOR2_X1 U761 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U762 ( .A1(G900), .A2(n713), .ZN(n714) );
  XOR2_X1 U763 ( .A(KEYINPUT125), .B(n714), .Z(n715) );
  NAND2_X1 U764 ( .A1(n715), .A2(G953), .ZN(n716) );
  NAND2_X1 U765 ( .A1(n717), .A2(n716), .ZN(G72) );
  XOR2_X1 U766 ( .A(n718), .B(G131), .Z(G33) );
  XOR2_X1 U767 ( .A(G137), .B(KEYINPUT126), .Z(n719) );
  XNOR2_X1 U768 ( .A(n720), .B(n719), .ZN(G39) );
  XNOR2_X1 U769 ( .A(n721), .B(G122), .ZN(G24) );
  XNOR2_X1 U770 ( .A(G125), .B(KEYINPUT37), .ZN(n723) );
  XNOR2_X1 U771 ( .A(n723), .B(n722), .ZN(G27) );
endmodule

