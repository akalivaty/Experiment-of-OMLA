

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U553 ( .A1(n1001), .A2(n701), .ZN(n702) );
  NOR2_X1 U554 ( .A1(n696), .A2(n695), .ZN(n698) );
  INV_X1 U555 ( .A(KEYINPUT93), .ZN(n710) );
  NAND2_X1 U556 ( .A1(n765), .A2(n1016), .ZN(n767) );
  AND2_X1 U557 ( .A1(n1005), .A2(n519), .ZN(n771) );
  NOR2_X1 U558 ( .A1(n579), .A2(n578), .ZN(n581) );
  OR2_X1 U559 ( .A1(n770), .A2(n781), .ZN(n519) );
  OR2_X1 U560 ( .A1(n769), .A2(KEYINPUT33), .ZN(n520) );
  INV_X1 U561 ( .A(KEYINPUT26), .ZN(n697) );
  XNOR2_X1 U562 ( .A(KEYINPUT94), .B(KEYINPUT30), .ZN(n730) );
  INV_X1 U563 ( .A(KEYINPUT29), .ZN(n721) );
  NOR2_X1 U564 ( .A1(G1966), .A2(n781), .ZN(n755) );
  INV_X1 U565 ( .A(KEYINPUT103), .ZN(n766) );
  XNOR2_X1 U566 ( .A(n767), .B(n766), .ZN(n768) );
  AND2_X1 U567 ( .A1(n783), .A2(n782), .ZN(n694) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n784) );
  INV_X1 U569 ( .A(KEYINPUT13), .ZN(n576) );
  INV_X1 U570 ( .A(G2105), .ZN(n522) );
  AND2_X2 U571 ( .A1(G2105), .A2(G2104), .ZN(n892) );
  NOR2_X1 U572 ( .A1(n646), .A2(G651), .ZN(n656) );
  XNOR2_X1 U573 ( .A(n558), .B(KEYINPUT65), .ZN(n783) );
  NOR2_X1 U574 ( .A1(n835), .A2(n834), .ZN(n837) );
  NAND2_X1 U575 ( .A1(n581), .A2(n580), .ZN(n1001) );
  NOR2_X1 U576 ( .A1(n530), .A2(n529), .ZN(G164) );
  INV_X1 U577 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U578 ( .A1(G2104), .A2(n525), .ZN(n555) );
  NAND2_X1 U579 ( .A1(G126), .A2(n555), .ZN(n521) );
  XOR2_X1 U580 ( .A(KEYINPUT85), .B(n521), .Z(n524) );
  AND2_X4 U581 ( .A1(n522), .A2(G2104), .ZN(n887) );
  NAND2_X1 U582 ( .A1(n887), .A2(G102), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n524), .A2(n523), .ZN(n530) );
  NAND2_X1 U584 ( .A1(G114), .A2(n892), .ZN(n528) );
  NOR2_X1 U585 ( .A1(G2105), .A2(G2104), .ZN(n526) );
  XOR2_X1 U586 ( .A(KEYINPUT17), .B(n526), .Z(n618) );
  NAND2_X1 U587 ( .A1(G138), .A2(n618), .ZN(n527) );
  NAND2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U589 ( .A(KEYINPUT0), .B(G543), .Z(n646) );
  INV_X1 U590 ( .A(G651), .ZN(n537) );
  NOR2_X2 U591 ( .A1(n646), .A2(n537), .ZN(n653) );
  NAND2_X1 U592 ( .A1(G76), .A2(n653), .ZN(n534) );
  XOR2_X1 U593 ( .A(KEYINPUT69), .B(KEYINPUT4), .Z(n532) );
  NOR2_X1 U594 ( .A1(G543), .A2(G651), .ZN(n652) );
  NAND2_X1 U595 ( .A1(G89), .A2(n652), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  NAND2_X1 U597 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n535), .B(KEYINPUT70), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n536), .B(KEYINPUT5), .ZN(n544) );
  NOR2_X1 U600 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X2 U601 ( .A(KEYINPUT1), .B(n538), .Z(n658) );
  NAND2_X1 U602 ( .A1(n658), .A2(G63), .ZN(n539) );
  XOR2_X1 U603 ( .A(KEYINPUT71), .B(n539), .Z(n541) );
  NAND2_X1 U604 ( .A1(n656), .A2(G51), .ZN(n540) );
  NAND2_X1 U605 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U606 ( .A(KEYINPUT6), .B(n542), .Z(n543) );
  NAND2_X1 U607 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U608 ( .A(n545), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U609 ( .A(G168), .B(KEYINPUT8), .Z(n546) );
  XNOR2_X1 U610 ( .A(KEYINPUT72), .B(n546), .ZN(G286) );
  NAND2_X1 U611 ( .A1(G60), .A2(n658), .ZN(n548) );
  NAND2_X1 U612 ( .A1(G85), .A2(n652), .ZN(n547) );
  NAND2_X1 U613 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U614 ( .A1(G72), .A2(n653), .ZN(n550) );
  NAND2_X1 U615 ( .A1(G47), .A2(n656), .ZN(n549) );
  NAND2_X1 U616 ( .A1(n550), .A2(n549), .ZN(n551) );
  OR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(G290) );
  NAND2_X1 U618 ( .A1(G113), .A2(n892), .ZN(n553) );
  XNOR2_X1 U619 ( .A(KEYINPUT66), .B(n553), .ZN(n691) );
  NAND2_X1 U620 ( .A1(n887), .A2(G101), .ZN(n554) );
  XOR2_X1 U621 ( .A(n554), .B(KEYINPUT23), .Z(n557) );
  BUF_X2 U622 ( .A(n555), .Z(n891) );
  NAND2_X1 U623 ( .A1(n891), .A2(G125), .ZN(n556) );
  NAND2_X1 U624 ( .A1(n557), .A2(n556), .ZN(n558) );
  NAND2_X1 U625 ( .A1(G137), .A2(n618), .ZN(n693) );
  AND2_X1 U626 ( .A1(n783), .A2(n693), .ZN(n559) );
  AND2_X1 U627 ( .A1(n691), .A2(n559), .ZN(G160) );
  XOR2_X1 U628 ( .A(G2430), .B(G2451), .Z(n561) );
  XNOR2_X1 U629 ( .A(KEYINPUT107), .B(G2443), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n561), .B(n560), .ZN(n568) );
  XOR2_X1 U631 ( .A(G2435), .B(G2446), .Z(n563) );
  XNOR2_X1 U632 ( .A(G2427), .B(G2454), .ZN(n562) );
  XNOR2_X1 U633 ( .A(n563), .B(n562), .ZN(n564) );
  XOR2_X1 U634 ( .A(n564), .B(G2438), .Z(n566) );
  XNOR2_X1 U635 ( .A(G1341), .B(G1348), .ZN(n565) );
  XNOR2_X1 U636 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U637 ( .A(n568), .B(n567), .ZN(n569) );
  AND2_X1 U638 ( .A1(n569), .A2(G14), .ZN(G401) );
  AND2_X1 U639 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U640 ( .A(G57), .ZN(G237) );
  INV_X1 U641 ( .A(G132), .ZN(G219) );
  INV_X1 U642 ( .A(G82), .ZN(G220) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n570) );
  XNOR2_X1 U644 ( .A(n570), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n838) );
  NAND2_X1 U646 ( .A1(n838), .A2(G567), .ZN(n571) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n571), .Z(G234) );
  NAND2_X1 U648 ( .A1(G56), .A2(n658), .ZN(n572) );
  XOR2_X1 U649 ( .A(KEYINPUT14), .B(n572), .Z(n579) );
  NAND2_X1 U650 ( .A1(G68), .A2(n653), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n652), .A2(G81), .ZN(n573) );
  XNOR2_X1 U652 ( .A(n573), .B(KEYINPUT12), .ZN(n574) );
  NAND2_X1 U653 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U654 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n656), .A2(G43), .ZN(n580) );
  INV_X1 U656 ( .A(G860), .ZN(n608) );
  OR2_X1 U657 ( .A1(n1001), .A2(n608), .ZN(G153) );
  NAND2_X1 U658 ( .A1(G90), .A2(n652), .ZN(n583) );
  NAND2_X1 U659 ( .A1(G77), .A2(n653), .ZN(n582) );
  NAND2_X1 U660 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U661 ( .A(KEYINPUT9), .B(n584), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G64), .A2(n658), .ZN(n586) );
  NAND2_X1 U663 ( .A1(G52), .A2(n656), .ZN(n585) );
  NAND2_X1 U664 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U665 ( .A(KEYINPUT67), .B(n587), .ZN(n588) );
  NAND2_X1 U666 ( .A1(n589), .A2(n588), .ZN(G301) );
  NAND2_X1 U667 ( .A1(G868), .A2(G301), .ZN(n598) );
  NAND2_X1 U668 ( .A1(G79), .A2(n653), .ZN(n591) );
  NAND2_X1 U669 ( .A1(G54), .A2(n656), .ZN(n590) );
  NAND2_X1 U670 ( .A1(n591), .A2(n590), .ZN(n595) );
  NAND2_X1 U671 ( .A1(G66), .A2(n658), .ZN(n593) );
  NAND2_X1 U672 ( .A1(G92), .A2(n652), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n594) );
  NOR2_X1 U674 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U675 ( .A(n596), .B(KEYINPUT15), .ZN(n609) );
  INV_X1 U676 ( .A(G868), .ZN(n672) );
  NAND2_X1 U677 ( .A1(n609), .A2(n672), .ZN(n597) );
  NAND2_X1 U678 ( .A1(n598), .A2(n597), .ZN(G284) );
  NAND2_X1 U679 ( .A1(G65), .A2(n658), .ZN(n600) );
  NAND2_X1 U680 ( .A1(G53), .A2(n656), .ZN(n599) );
  NAND2_X1 U681 ( .A1(n600), .A2(n599), .ZN(n604) );
  NAND2_X1 U682 ( .A1(G91), .A2(n652), .ZN(n602) );
  NAND2_X1 U683 ( .A1(G78), .A2(n653), .ZN(n601) );
  NAND2_X1 U684 ( .A1(n602), .A2(n601), .ZN(n603) );
  NOR2_X1 U685 ( .A1(n604), .A2(n603), .ZN(n1015) );
  XOR2_X1 U686 ( .A(n1015), .B(KEYINPUT68), .Z(G299) );
  XNOR2_X1 U687 ( .A(KEYINPUT73), .B(G868), .ZN(n605) );
  NOR2_X1 U688 ( .A1(G286), .A2(n605), .ZN(n607) );
  NOR2_X1 U689 ( .A1(G299), .A2(G868), .ZN(n606) );
  NOR2_X1 U690 ( .A1(n607), .A2(n606), .ZN(G297) );
  NAND2_X1 U691 ( .A1(n608), .A2(G559), .ZN(n610) );
  INV_X1 U692 ( .A(n609), .ZN(n1008) );
  NAND2_X1 U693 ( .A1(n610), .A2(n1008), .ZN(n611) );
  XNOR2_X1 U694 ( .A(n611), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U695 ( .A1(n1008), .A2(G868), .ZN(n612) );
  NOR2_X1 U696 ( .A1(G559), .A2(n612), .ZN(n613) );
  XNOR2_X1 U697 ( .A(n613), .B(KEYINPUT74), .ZN(n615) );
  NOR2_X1 U698 ( .A1(n1001), .A2(G868), .ZN(n614) );
  NOR2_X1 U699 ( .A1(n615), .A2(n614), .ZN(G282) );
  NAND2_X1 U700 ( .A1(G99), .A2(n887), .ZN(n617) );
  NAND2_X1 U701 ( .A1(G111), .A2(n892), .ZN(n616) );
  NAND2_X1 U702 ( .A1(n617), .A2(n616), .ZN(n625) );
  BUF_X1 U703 ( .A(n618), .Z(n888) );
  NAND2_X1 U704 ( .A1(n888), .A2(G135), .ZN(n619) );
  XNOR2_X1 U705 ( .A(KEYINPUT75), .B(n619), .ZN(n622) );
  NAND2_X1 U706 ( .A1(n891), .A2(G123), .ZN(n620) );
  XOR2_X1 U707 ( .A(KEYINPUT18), .B(n620), .Z(n621) );
  NOR2_X1 U708 ( .A1(n622), .A2(n621), .ZN(n623) );
  XOR2_X1 U709 ( .A(KEYINPUT76), .B(n623), .Z(n624) );
  NOR2_X1 U710 ( .A1(n625), .A2(n624), .ZN(n935) );
  XNOR2_X1 U711 ( .A(n935), .B(G2096), .ZN(n627) );
  INV_X1 U712 ( .A(G2100), .ZN(n626) );
  NAND2_X1 U713 ( .A1(n627), .A2(n626), .ZN(G156) );
  NAND2_X1 U714 ( .A1(G67), .A2(n658), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G93), .A2(n652), .ZN(n628) );
  NAND2_X1 U716 ( .A1(n629), .A2(n628), .ZN(n632) );
  NAND2_X1 U717 ( .A1(G55), .A2(n656), .ZN(n630) );
  XNOR2_X1 U718 ( .A(KEYINPUT77), .B(n630), .ZN(n631) );
  NOR2_X1 U719 ( .A1(n632), .A2(n631), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n653), .A2(G80), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(n671) );
  NAND2_X1 U722 ( .A1(G559), .A2(n1008), .ZN(n635) );
  XNOR2_X1 U723 ( .A(n635), .B(n1001), .ZN(n669) );
  NOR2_X1 U724 ( .A1(G860), .A2(n669), .ZN(n636) );
  XOR2_X1 U725 ( .A(n671), .B(n636), .Z(G145) );
  XOR2_X1 U726 ( .A(KEYINPUT78), .B(KEYINPUT2), .Z(n638) );
  NAND2_X1 U727 ( .A1(G73), .A2(n653), .ZN(n637) );
  XNOR2_X1 U728 ( .A(n638), .B(n637), .ZN(n642) );
  NAND2_X1 U729 ( .A1(n652), .A2(G86), .ZN(n640) );
  NAND2_X1 U730 ( .A1(n658), .A2(G61), .ZN(n639) );
  NAND2_X1 U731 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U732 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U733 ( .A(KEYINPUT79), .B(n643), .Z(n645) );
  NAND2_X1 U734 ( .A1(n656), .A2(G48), .ZN(n644) );
  NAND2_X1 U735 ( .A1(n645), .A2(n644), .ZN(G305) );
  NAND2_X1 U736 ( .A1(G49), .A2(n656), .ZN(n648) );
  NAND2_X1 U737 ( .A1(G87), .A2(n646), .ZN(n647) );
  NAND2_X1 U738 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U739 ( .A1(n658), .A2(n649), .ZN(n651) );
  NAND2_X1 U740 ( .A1(G651), .A2(G74), .ZN(n650) );
  NAND2_X1 U741 ( .A1(n651), .A2(n650), .ZN(G288) );
  NAND2_X1 U742 ( .A1(G88), .A2(n652), .ZN(n655) );
  NAND2_X1 U743 ( .A1(G75), .A2(n653), .ZN(n654) );
  NAND2_X1 U744 ( .A1(n655), .A2(n654), .ZN(n662) );
  NAND2_X1 U745 ( .A1(G50), .A2(n656), .ZN(n657) );
  XNOR2_X1 U746 ( .A(n657), .B(KEYINPUT80), .ZN(n660) );
  NAND2_X1 U747 ( .A1(n658), .A2(G62), .ZN(n659) );
  NAND2_X1 U748 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U749 ( .A1(n662), .A2(n661), .ZN(G166) );
  INV_X1 U750 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U751 ( .A(G299), .B(G305), .ZN(n663) );
  XNOR2_X1 U752 ( .A(n663), .B(n671), .ZN(n664) );
  XNOR2_X1 U753 ( .A(KEYINPUT81), .B(n664), .ZN(n666) );
  XNOR2_X1 U754 ( .A(G288), .B(KEYINPUT19), .ZN(n665) );
  XNOR2_X1 U755 ( .A(n666), .B(n665), .ZN(n667) );
  XNOR2_X1 U756 ( .A(n667), .B(G303), .ZN(n668) );
  XNOR2_X1 U757 ( .A(n668), .B(G290), .ZN(n911) );
  XNOR2_X1 U758 ( .A(n669), .B(n911), .ZN(n670) );
  NAND2_X1 U759 ( .A1(n670), .A2(G868), .ZN(n674) );
  NAND2_X1 U760 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U761 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U762 ( .A1(G2084), .A2(G2078), .ZN(n675) );
  XOR2_X1 U763 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U764 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U765 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U766 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U767 ( .A(KEYINPUT82), .B(G44), .ZN(n679) );
  XNOR2_X1 U768 ( .A(n679), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U769 ( .A1(G220), .A2(G219), .ZN(n680) );
  XOR2_X1 U770 ( .A(KEYINPUT22), .B(n680), .Z(n681) );
  NOR2_X1 U771 ( .A1(G218), .A2(n681), .ZN(n682) );
  XOR2_X1 U772 ( .A(KEYINPUT83), .B(n682), .Z(n683) );
  NAND2_X1 U773 ( .A1(G96), .A2(n683), .ZN(n843) );
  NAND2_X1 U774 ( .A1(G2106), .A2(n843), .ZN(n687) );
  NAND2_X1 U775 ( .A1(G69), .A2(G120), .ZN(n684) );
  NOR2_X1 U776 ( .A1(G237), .A2(n684), .ZN(n685) );
  NAND2_X1 U777 ( .A1(G108), .A2(n685), .ZN(n844) );
  NAND2_X1 U778 ( .A1(G567), .A2(n844), .ZN(n686) );
  NAND2_X1 U779 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U780 ( .A(KEYINPUT84), .B(n688), .Z(G319) );
  INV_X1 U781 ( .A(G319), .ZN(n690) );
  NAND2_X1 U782 ( .A1(G661), .A2(G483), .ZN(n689) );
  NOR2_X1 U783 ( .A1(n690), .A2(n689), .ZN(n842) );
  NAND2_X1 U784 ( .A1(n842), .A2(G36), .ZN(G176) );
  INV_X1 U785 ( .A(G301), .ZN(G171) );
  AND2_X1 U786 ( .A1(G40), .A2(n691), .ZN(n692) );
  AND2_X1 U787 ( .A1(n693), .A2(n692), .ZN(n782) );
  NAND2_X1 U788 ( .A1(n694), .A2(n784), .ZN(n696) );
  BUF_X2 U789 ( .A(n696), .Z(n741) );
  NAND2_X1 U790 ( .A1(G8), .A2(n741), .ZN(n781) );
  NAND2_X1 U791 ( .A1(n741), .A2(G1341), .ZN(n700) );
  INV_X1 U792 ( .A(G1996), .ZN(n695) );
  XNOR2_X1 U793 ( .A(n698), .B(n697), .ZN(n699) );
  NAND2_X1 U794 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U795 ( .A(n702), .B(KEYINPUT64), .ZN(n707) );
  NAND2_X1 U796 ( .A1(n707), .A2(n1008), .ZN(n706) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n741), .ZN(n704) );
  INV_X1 U798 ( .A(n741), .ZN(n723) );
  NOR2_X1 U799 ( .A1(n723), .A2(G1348), .ZN(n703) );
  NOR2_X1 U800 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U801 ( .A1(n706), .A2(n705), .ZN(n709) );
  OR2_X1 U802 ( .A1(n707), .A2(n1008), .ZN(n708) );
  NAND2_X1 U803 ( .A1(n709), .A2(n708), .ZN(n711) );
  XNOR2_X1 U804 ( .A(n711), .B(n710), .ZN(n716) );
  NAND2_X1 U805 ( .A1(n723), .A2(G2072), .ZN(n712) );
  XNOR2_X1 U806 ( .A(n712), .B(KEYINPUT27), .ZN(n714) );
  AND2_X1 U807 ( .A1(G1956), .A2(n741), .ZN(n713) );
  NOR2_X1 U808 ( .A1(n714), .A2(n713), .ZN(n717) );
  NAND2_X1 U809 ( .A1(n717), .A2(n1015), .ZN(n715) );
  NAND2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n720) );
  NOR2_X1 U811 ( .A1(n717), .A2(n1015), .ZN(n718) );
  XOR2_X1 U812 ( .A(n718), .B(KEYINPUT28), .Z(n719) );
  NAND2_X1 U813 ( .A1(n720), .A2(n719), .ZN(n722) );
  XNOR2_X1 U814 ( .A(n722), .B(n721), .ZN(n728) );
  XNOR2_X1 U815 ( .A(KEYINPUT25), .B(G2078), .ZN(n955) );
  NAND2_X1 U816 ( .A1(n723), .A2(n955), .ZN(n724) );
  XNOR2_X1 U817 ( .A(n724), .B(KEYINPUT92), .ZN(n726) );
  INV_X1 U818 ( .A(G1961), .ZN(n973) );
  NAND2_X1 U819 ( .A1(n973), .A2(n741), .ZN(n725) );
  NAND2_X1 U820 ( .A1(n726), .A2(n725), .ZN(n734) );
  NAND2_X1 U821 ( .A1(n734), .A2(G171), .ZN(n727) );
  NAND2_X1 U822 ( .A1(n728), .A2(n727), .ZN(n740) );
  XNOR2_X1 U823 ( .A(KEYINPUT31), .B(KEYINPUT96), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G2084), .A2(n741), .ZN(n752) );
  NOR2_X1 U825 ( .A1(n752), .A2(n755), .ZN(n729) );
  NAND2_X1 U826 ( .A1(G8), .A2(n729), .ZN(n731) );
  XNOR2_X1 U827 ( .A(n731), .B(n730), .ZN(n732) );
  NOR2_X1 U828 ( .A1(G168), .A2(n732), .ZN(n733) );
  XNOR2_X1 U829 ( .A(n733), .B(KEYINPUT95), .ZN(n736) );
  OR2_X1 U830 ( .A1(n734), .A2(G171), .ZN(n735) );
  NAND2_X1 U831 ( .A1(n736), .A2(n735), .ZN(n737) );
  XNOR2_X1 U832 ( .A(n738), .B(n737), .ZN(n739) );
  NAND2_X1 U833 ( .A1(n740), .A2(n739), .ZN(n753) );
  NAND2_X1 U834 ( .A1(n753), .A2(G286), .ZN(n748) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n741), .ZN(n742) );
  XOR2_X1 U836 ( .A(KEYINPUT99), .B(n742), .Z(n745) );
  NOR2_X1 U837 ( .A1(G1971), .A2(n781), .ZN(n743) );
  XNOR2_X1 U838 ( .A(n743), .B(KEYINPUT98), .ZN(n744) );
  NOR2_X1 U839 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U840 ( .A1(n746), .A2(G303), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(n749) );
  XNOR2_X1 U842 ( .A(n749), .B(KEYINPUT100), .ZN(n750) );
  NAND2_X1 U843 ( .A1(n750), .A2(G8), .ZN(n751) );
  XNOR2_X1 U844 ( .A(n751), .B(KEYINPUT32), .ZN(n760) );
  NAND2_X1 U845 ( .A1(G8), .A2(n752), .ZN(n758) );
  INV_X1 U846 ( .A(n753), .ZN(n754) );
  NOR2_X1 U847 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U848 ( .A(KEYINPUT97), .B(n756), .Z(n757) );
  NAND2_X1 U849 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U850 ( .A1(n760), .A2(n759), .ZN(n772) );
  NOR2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n1023) );
  NOR2_X1 U852 ( .A1(G1971), .A2(G303), .ZN(n761) );
  XOR2_X1 U853 ( .A(n761), .B(KEYINPUT101), .Z(n762) );
  NOR2_X1 U854 ( .A1(n1023), .A2(n762), .ZN(n763) );
  XNOR2_X1 U855 ( .A(n763), .B(KEYINPUT102), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n772), .A2(n764), .ZN(n765) );
  NAND2_X1 U857 ( .A1(G1976), .A2(G288), .ZN(n1016) );
  NOR2_X1 U858 ( .A1(n781), .A2(n768), .ZN(n769) );
  XOR2_X1 U859 ( .A(G1981), .B(G305), .Z(n1005) );
  NAND2_X1 U860 ( .A1(n1023), .A2(KEYINPUT33), .ZN(n770) );
  NAND2_X1 U861 ( .A1(n520), .A2(n771), .ZN(n777) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n773) );
  NAND2_X1 U863 ( .A1(G8), .A2(n773), .ZN(n774) );
  NAND2_X1 U864 ( .A1(n772), .A2(n774), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n775), .A2(n781), .ZN(n776) );
  NAND2_X1 U866 ( .A1(n777), .A2(n776), .ZN(n778) );
  XNOR2_X1 U867 ( .A(n778), .B(KEYINPUT104), .ZN(n825) );
  NOR2_X1 U868 ( .A1(G1981), .A2(G305), .ZN(n779) );
  XOR2_X1 U869 ( .A(n779), .B(KEYINPUT24), .Z(n780) );
  NOR2_X1 U870 ( .A1(n781), .A2(n780), .ZN(n823) );
  NAND2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n785) );
  NOR2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n826) );
  NAND2_X1 U873 ( .A1(G105), .A2(n887), .ZN(n786) );
  XNOR2_X1 U874 ( .A(n786), .B(KEYINPUT38), .ZN(n793) );
  NAND2_X1 U875 ( .A1(G129), .A2(n891), .ZN(n788) );
  NAND2_X1 U876 ( .A1(G141), .A2(n888), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n788), .A2(n787), .ZN(n791) );
  NAND2_X1 U878 ( .A1(G117), .A2(n892), .ZN(n789) );
  XNOR2_X1 U879 ( .A(KEYINPUT91), .B(n789), .ZN(n790) );
  NOR2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n792) );
  NAND2_X1 U881 ( .A1(n793), .A2(n792), .ZN(n877) );
  NOR2_X1 U882 ( .A1(G1996), .A2(n877), .ZN(n933) );
  NAND2_X1 U883 ( .A1(n887), .A2(G95), .ZN(n794) );
  XNOR2_X1 U884 ( .A(n794), .B(KEYINPUT88), .ZN(n796) );
  NAND2_X1 U885 ( .A1(G131), .A2(n888), .ZN(n795) );
  NAND2_X1 U886 ( .A1(n796), .A2(n795), .ZN(n797) );
  XNOR2_X1 U887 ( .A(KEYINPUT89), .B(n797), .ZN(n801) );
  NAND2_X1 U888 ( .A1(n891), .A2(G119), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G107), .A2(n892), .ZN(n798) );
  AND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U891 ( .A1(n801), .A2(n800), .ZN(n874) );
  XNOR2_X1 U892 ( .A(KEYINPUT90), .B(G1991), .ZN(n951) );
  NAND2_X1 U893 ( .A1(n874), .A2(n951), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G1996), .A2(n877), .ZN(n802) );
  NAND2_X1 U895 ( .A1(n803), .A2(n802), .ZN(n926) );
  AND2_X1 U896 ( .A1(n826), .A2(n926), .ZN(n830) );
  NOR2_X1 U897 ( .A1(G1986), .A2(G290), .ZN(n804) );
  NOR2_X1 U898 ( .A1(n951), .A2(n874), .ZN(n936) );
  NOR2_X1 U899 ( .A1(n804), .A2(n936), .ZN(n805) );
  NOR2_X1 U900 ( .A1(n830), .A2(n805), .ZN(n806) );
  NOR2_X1 U901 ( .A1(n933), .A2(n806), .ZN(n807) );
  XNOR2_X1 U902 ( .A(n807), .B(KEYINPUT39), .ZN(n818) );
  XNOR2_X1 U903 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NAND2_X1 U904 ( .A1(G104), .A2(n887), .ZN(n809) );
  NAND2_X1 U905 ( .A1(G140), .A2(n888), .ZN(n808) );
  NAND2_X1 U906 ( .A1(n809), .A2(n808), .ZN(n811) );
  XOR2_X1 U907 ( .A(KEYINPUT87), .B(KEYINPUT34), .Z(n810) );
  XNOR2_X1 U908 ( .A(n811), .B(n810), .ZN(n816) );
  NAND2_X1 U909 ( .A1(G128), .A2(n891), .ZN(n813) );
  NAND2_X1 U910 ( .A1(G116), .A2(n892), .ZN(n812) );
  NAND2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  XOR2_X1 U912 ( .A(KEYINPUT35), .B(n814), .Z(n815) );
  NOR2_X1 U913 ( .A1(n816), .A2(n815), .ZN(n817) );
  XNOR2_X1 U914 ( .A(KEYINPUT36), .B(n817), .ZN(n904) );
  NOR2_X1 U915 ( .A1(n819), .A2(n904), .ZN(n929) );
  NAND2_X1 U916 ( .A1(n826), .A2(n929), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n818), .A2(n828), .ZN(n820) );
  NAND2_X1 U918 ( .A1(n819), .A2(n904), .ZN(n927) );
  NAND2_X1 U919 ( .A1(n820), .A2(n927), .ZN(n821) );
  XOR2_X1 U920 ( .A(KEYINPUT105), .B(n821), .Z(n822) );
  AND2_X1 U921 ( .A1(n826), .A2(n822), .ZN(n833) );
  OR2_X1 U922 ( .A1(n823), .A2(n833), .ZN(n824) );
  NOR2_X1 U923 ( .A1(n825), .A2(n824), .ZN(n835) );
  XNOR2_X1 U924 ( .A(G1986), .B(G290), .ZN(n1019) );
  NAND2_X1 U925 ( .A1(n1019), .A2(n826), .ZN(n827) );
  XNOR2_X1 U926 ( .A(n827), .B(KEYINPUT86), .ZN(n829) );
  NAND2_X1 U927 ( .A1(n829), .A2(n828), .ZN(n831) );
  NOR2_X1 U928 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U929 ( .A1(n833), .A2(n832), .ZN(n834) );
  XNOR2_X1 U930 ( .A(KEYINPUT106), .B(KEYINPUT40), .ZN(n836) );
  XNOR2_X1 U931 ( .A(n837), .B(n836), .ZN(G329) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n838), .ZN(G217) );
  NAND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n839) );
  XOR2_X1 U934 ( .A(KEYINPUT108), .B(n839), .Z(n840) );
  NAND2_X1 U935 ( .A1(G661), .A2(n840), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n841) );
  NAND2_X1 U937 ( .A1(n842), .A2(n841), .ZN(G188) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n844), .A2(n843), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  XOR2_X1 U944 ( .A(KEYINPUT110), .B(G1991), .Z(n846) );
  XNOR2_X1 U945 ( .A(G1956), .B(G1996), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U947 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U948 ( .A(G1981), .B(G1966), .ZN(n848) );
  XNOR2_X1 U949 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U950 ( .A(G1986), .B(G1976), .Z(n851) );
  XNOR2_X1 U951 ( .A(G1961), .B(G1971), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U953 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U954 ( .A(KEYINPUT41), .B(KEYINPUT111), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(G229) );
  XOR2_X1 U956 ( .A(G2678), .B(G2072), .Z(n857) );
  XNOR2_X1 U957 ( .A(G2090), .B(G2084), .ZN(n856) );
  XNOR2_X1 U958 ( .A(n857), .B(n856), .ZN(n858) );
  XOR2_X1 U959 ( .A(n858), .B(G2100), .Z(n860) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2067), .ZN(n859) );
  XNOR2_X1 U961 ( .A(n860), .B(n859), .ZN(n864) );
  XOR2_X1 U962 ( .A(G2096), .B(KEYINPUT109), .Z(n862) );
  XNOR2_X1 U963 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n861) );
  XNOR2_X1 U964 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U965 ( .A(n864), .B(n863), .Z(G227) );
  NAND2_X1 U966 ( .A1(n891), .A2(G124), .ZN(n865) );
  XNOR2_X1 U967 ( .A(n865), .B(KEYINPUT44), .ZN(n867) );
  NAND2_X1 U968 ( .A1(G136), .A2(n888), .ZN(n866) );
  NAND2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT112), .B(n868), .Z(n870) );
  NAND2_X1 U971 ( .A1(n887), .A2(G100), .ZN(n869) );
  NAND2_X1 U972 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U973 ( .A1(G112), .A2(n892), .ZN(n871) );
  XNOR2_X1 U974 ( .A(KEYINPUT113), .B(n871), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U976 ( .A(G162), .B(n874), .ZN(n907) );
  XOR2_X1 U977 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n876) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n875) );
  XNOR2_X1 U979 ( .A(n876), .B(n875), .ZN(n878) );
  XOR2_X1 U980 ( .A(n878), .B(n877), .Z(n902) );
  NAND2_X1 U981 ( .A1(G130), .A2(n891), .ZN(n880) );
  NAND2_X1 U982 ( .A1(G118), .A2(n892), .ZN(n879) );
  NAND2_X1 U983 ( .A1(n880), .A2(n879), .ZN(n886) );
  NAND2_X1 U984 ( .A1(n888), .A2(G142), .ZN(n881) );
  XNOR2_X1 U985 ( .A(n881), .B(KEYINPUT114), .ZN(n883) );
  NAND2_X1 U986 ( .A1(G106), .A2(n887), .ZN(n882) );
  NAND2_X1 U987 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U988 ( .A(KEYINPUT45), .B(n884), .Z(n885) );
  NOR2_X1 U989 ( .A1(n886), .A2(n885), .ZN(n900) );
  XNOR2_X1 U990 ( .A(G164), .B(n935), .ZN(n898) );
  NAND2_X1 U991 ( .A1(G103), .A2(n887), .ZN(n890) );
  NAND2_X1 U992 ( .A1(G139), .A2(n888), .ZN(n889) );
  NAND2_X1 U993 ( .A1(n890), .A2(n889), .ZN(n897) );
  NAND2_X1 U994 ( .A1(G127), .A2(n891), .ZN(n894) );
  NAND2_X1 U995 ( .A1(G115), .A2(n892), .ZN(n893) );
  NAND2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U997 ( .A(KEYINPUT47), .B(n895), .Z(n896) );
  NOR2_X1 U998 ( .A1(n897), .A2(n896), .ZN(n921) );
  XNOR2_X1 U999 ( .A(n898), .B(n921), .ZN(n899) );
  XOR2_X1 U1000 ( .A(n900), .B(n899), .Z(n901) );
  XNOR2_X1 U1001 ( .A(n902), .B(n901), .ZN(n903) );
  XNOR2_X1 U1002 ( .A(G160), .B(n903), .ZN(n905) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1005 ( .A1(G37), .A2(n908), .ZN(G395) );
  XNOR2_X1 U1006 ( .A(n1001), .B(KEYINPUT117), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(G171), .B(n1008), .ZN(n909) );
  XNOR2_X1 U1008 ( .A(n910), .B(n909), .ZN(n913) );
  XNOR2_X1 U1009 ( .A(G286), .B(n911), .ZN(n912) );
  XNOR2_X1 U1010 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n914), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n915) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n916), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n917), .ZN(n920) );
  NOR2_X1 U1016 ( .A1(G395), .A2(G397), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(n918), .B(KEYINPUT118), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XOR2_X1 U1021 ( .A(G2072), .B(n921), .Z(n923) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XOR2_X1 U1024 ( .A(KEYINPUT50), .B(n924), .Z(n944) );
  XOR2_X1 U1025 ( .A(G160), .B(G2084), .Z(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n931) );
  INV_X1 U1027 ( .A(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n941) );
  XOR2_X1 U1030 ( .A(G2090), .B(G162), .Z(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n934), .Z(n939) );
  NOR2_X1 U1033 ( .A1(n936), .A2(n935), .ZN(n937) );
  XOR2_X1 U1034 ( .A(KEYINPUT119), .B(n937), .Z(n938) );
  NAND2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1037 ( .A(KEYINPUT120), .B(n942), .Z(n943) );
  NOR2_X1 U1038 ( .A1(n944), .A2(n943), .ZN(n945) );
  XOR2_X1 U1039 ( .A(KEYINPUT52), .B(n945), .Z(n946) );
  NOR2_X1 U1040 ( .A1(KEYINPUT55), .A2(n946), .ZN(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n947), .ZN(n948) );
  NAND2_X1 U1042 ( .A1(n948), .A2(G29), .ZN(n1000) );
  XOR2_X1 U1043 ( .A(G2072), .B(G33), .Z(n950) );
  XOR2_X1 U1044 ( .A(G1996), .B(G32), .Z(n949) );
  NAND2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n953) );
  XNOR2_X1 U1046 ( .A(G25), .B(n951), .ZN(n952) );
  NOR2_X1 U1047 ( .A1(n953), .A2(n952), .ZN(n959) );
  XOR2_X1 U1048 ( .A(G2067), .B(G26), .Z(n954) );
  NAND2_X1 U1049 ( .A1(n954), .A2(G28), .ZN(n957) );
  XOR2_X1 U1050 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(KEYINPUT53), .B(n960), .ZN(n962) );
  XOR2_X1 U1054 ( .A(G2090), .B(G35), .Z(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n967) );
  XOR2_X1 U1056 ( .A(KEYINPUT122), .B(G34), .Z(n964) );
  XNOR2_X1 U1057 ( .A(KEYINPUT54), .B(KEYINPUT123), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n964), .B(n963), .ZN(n965) );
  XNOR2_X1 U1059 ( .A(n965), .B(G2084), .ZN(n966) );
  NOR2_X1 U1060 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT55), .B(n968), .ZN(n970) );
  INV_X1 U1062 ( .A(G29), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n971), .A2(G11), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT124), .ZN(n998) );
  XNOR2_X1 U1066 ( .A(G5), .B(n973), .ZN(n994) );
  XOR2_X1 U1067 ( .A(G1966), .B(G21), .Z(n984) );
  XNOR2_X1 U1068 ( .A(G1348), .B(KEYINPUT59), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(n974), .B(G4), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(G1956), .B(G20), .ZN(n976) );
  XNOR2_X1 U1071 ( .A(G19), .B(G1341), .ZN(n975) );
  NOR2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n981) );
  XNOR2_X1 U1074 ( .A(G6), .B(G1981), .ZN(n979) );
  XNOR2_X1 U1075 ( .A(KEYINPUT126), .B(n979), .ZN(n980) );
  NOR2_X1 U1076 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT60), .B(n982), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n992) );
  XNOR2_X1 U1079 ( .A(KEYINPUT58), .B(KEYINPUT127), .ZN(n990) );
  XOR2_X1 U1080 ( .A(G1976), .B(G23), .Z(n988) );
  XNOR2_X1 U1081 ( .A(G1971), .B(G22), .ZN(n986) );
  XNOR2_X1 U1082 ( .A(G24), .B(G1986), .ZN(n985) );
  NOR2_X1 U1083 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1084 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1085 ( .A(n990), .B(n989), .Z(n991) );
  NOR2_X1 U1086 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1087 ( .A1(n994), .A2(n993), .ZN(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT61), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n996), .A2(G16), .ZN(n997) );
  NOR2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1027) );
  XOR2_X1 U1092 ( .A(KEYINPUT56), .B(G16), .Z(n1025) );
  XNOR2_X1 U1093 ( .A(G1341), .B(KEYINPUT125), .ZN(n1002) );
  XNOR2_X1 U1094 ( .A(n1002), .B(n1001), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(G171), .B(G1961), .ZN(n1003) );
  NAND2_X1 U1096 ( .A1(n1004), .A2(n1003), .ZN(n1014) );
  XNOR2_X1 U1097 ( .A(G1966), .B(G168), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1099 ( .A(n1007), .B(KEYINPUT57), .ZN(n1012) );
  XOR2_X1 U1100 ( .A(n1008), .B(G1348), .Z(n1010) );
  XOR2_X1 U1101 ( .A(G166), .B(G1971), .Z(n1009) );
  NOR2_X1 U1102 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1021) );
  XNOR2_X1 U1105 ( .A(n1015), .B(G1956), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NOR2_X1 U1109 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NOR2_X1 U1111 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1112 ( .A(n1028), .B(KEYINPUT62), .ZN(G311) );
  INV_X1 U1113 ( .A(G311), .ZN(G150) );
endmodule

