//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n574, new_n575, new_n576,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n623,
    new_n624, new_n627, new_n629, new_n630, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n840, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1221, new_n1222, new_n1223, new_n1225;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  AND2_X1   g016(.A1(G2072), .A2(G2078), .ZN(new_n442));
  NAND3_X1  g017(.A1(new_n442), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT67), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT68), .Z(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n457), .A2(G567), .ZN(new_n460));
  INV_X1    g035(.A(G2106), .ZN(new_n461));
  OAI21_X1  g036(.A(new_n460), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  XNOR2_X1  g038(.A(KEYINPUT3), .B(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n464), .A2(G137), .A3(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G101), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n472), .B1(new_n464), .B2(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(KEYINPUT69), .B1(new_n473), .B2(new_n465), .ZN(new_n474));
  AND2_X1   g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NOR2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  OAI21_X1  g051(.A(G125), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(new_n471), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n470), .B1(new_n474), .B2(new_n480), .ZN(G160));
  NOR2_X1   g056(.A1(new_n475), .A2(new_n476), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n482), .A2(new_n465), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  INV_X1    g061(.A(G100), .ZN(new_n487));
  AND3_X1   g062(.A1(new_n487), .A2(new_n465), .A3(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g063(.A(KEYINPUT70), .B1(new_n487), .B2(new_n465), .ZN(new_n489));
  OAI221_X1 g064(.A(G2104), .B1(G112), .B2(new_n465), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n484), .A2(new_n486), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI21_X1  g067(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT71), .ZN(new_n495));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n495), .A2(new_n496), .A3(G2105), .ZN(new_n497));
  OAI21_X1  g072(.A(KEYINPUT71), .B1(new_n465), .B2(G114), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n494), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  OAI211_X1 g074(.A(G126), .B(G2105), .C1(new_n475), .C2(new_n476), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n464), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT4), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n503), .B(new_n506), .C1(new_n476), .C2(new_n475), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n501), .B1(new_n505), .B2(new_n507), .ZN(G164));
  XNOR2_X1  g083(.A(KEYINPUT5), .B(G543), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n509), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n509), .A2(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(G50), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(new_n511), .ZN(new_n516));
  NAND2_X1  g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n513), .A2(new_n514), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n512), .A2(new_n518), .ZN(G166));
  AND2_X1   g094(.A1(KEYINPUT6), .A2(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(KEYINPUT6), .A2(G651), .ZN(new_n521));
  OAI21_X1  g096(.A(KEYINPUT72), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT72), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n516), .A2(new_n523), .A3(new_n517), .ZN(new_n524));
  AND3_X1   g099(.A1(new_n522), .A2(new_n524), .A3(G543), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G51), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n509), .A2(G63), .A3(G651), .ZN(new_n529));
  AND2_X1   g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(G89), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n516), .A2(new_n517), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n532), .A2(new_n509), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n526), .B(new_n530), .C1(new_n531), .C2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(G168));
  AOI22_X1  g110(.A1(new_n509), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n511), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n525), .A2(G52), .ZN(new_n538));
  INV_X1    g113(.A(new_n533), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G90), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n537), .A2(new_n538), .A3(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n509), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n543), .A2(new_n511), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n525), .A2(G43), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n539), .A2(G81), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  XOR2_X1   g125(.A(KEYINPUT73), .B(KEYINPUT8), .Z(new_n551));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n551), .B(new_n552), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(new_n554));
  XOR2_X1   g129(.A(new_n554), .B(KEYINPUT74), .Z(G188));
  NAND3_X1  g130(.A1(new_n522), .A2(new_n524), .A3(G543), .ZN(new_n556));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n532), .B2(KEYINPUT72), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(new_n524), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n532), .A2(new_n509), .A3(G91), .ZN(new_n564));
  INV_X1    g139(.A(G78), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n565), .A2(new_n559), .ZN(new_n566));
  AOI21_X1  g141(.A(new_n566), .B1(new_n509), .B2(G65), .ZN(new_n567));
  OAI21_X1  g142(.A(new_n564), .B1(new_n567), .B2(new_n511), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n563), .A2(new_n569), .ZN(G299));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n534), .B(new_n571), .ZN(G286));
  INV_X1    g147(.A(G166), .ZN(G303));
  OAI21_X1  g148(.A(G651), .B1(new_n509), .B2(G74), .ZN(new_n574));
  INV_X1    g149(.A(G87), .ZN(new_n575));
  INV_X1    g150(.A(G49), .ZN(new_n576));
  OAI221_X1 g151(.A(new_n574), .B1(new_n533), .B2(new_n575), .C1(new_n556), .C2(new_n576), .ZN(G288));
  NAND2_X1  g152(.A1(G73), .A2(G543), .ZN(new_n578));
  NAND2_X1  g153(.A1(KEYINPUT5), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(KEYINPUT5), .A2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g159(.A1(G48), .A2(G543), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n584), .A2(G651), .B1(new_n532), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n532), .A2(new_n509), .A3(G86), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(G305));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  INV_X1    g164(.A(G60), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT5), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n591), .A2(new_n559), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n590), .B1(new_n592), .B2(new_n579), .ZN(new_n593));
  NAND2_X1  g168(.A1(G72), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(new_n594), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n589), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  OAI211_X1 g171(.A(KEYINPUT76), .B(new_n594), .C1(new_n582), .C2(new_n590), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n596), .A2(new_n597), .A3(G651), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT77), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT77), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n596), .A2(new_n597), .A3(new_n600), .A4(G651), .ZN(new_n601));
  INV_X1    g176(.A(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n556), .A2(new_n602), .B1(new_n603), .B2(new_n533), .ZN(new_n604));
  INV_X1    g179(.A(new_n604), .ZN(new_n605));
  AND4_X1   g180(.A1(KEYINPUT78), .A2(new_n599), .A3(new_n601), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n604), .B1(new_n598), .B2(KEYINPUT77), .ZN(new_n607));
  AOI21_X1  g182(.A(KEYINPUT78), .B1(new_n607), .B2(new_n601), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  NAND2_X1  g185(.A1(G301), .A2(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n525), .A2(G54), .ZN(new_n612));
  AOI22_X1  g187(.A1(new_n509), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n613));
  OR2_X1    g188(.A1(new_n613), .A2(new_n511), .ZN(new_n614));
  AOI21_X1  g189(.A(KEYINPUT10), .B1(new_n539), .B2(G92), .ZN(new_n615));
  AND4_X1   g190(.A1(KEYINPUT10), .A2(new_n532), .A3(new_n509), .A4(G92), .ZN(new_n616));
  OAI211_X1 g191(.A(new_n612), .B(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G868), .ZN(G284));
  OAI21_X1  g194(.A(new_n611), .B1(new_n618), .B2(G868), .ZN(G321));
  AOI21_X1  g195(.A(new_n568), .B1(new_n558), .B2(new_n562), .ZN(new_n621));
  INV_X1    g196(.A(G868), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G286), .B2(new_n622), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT79), .ZN(G297));
  XOR2_X1   g200(.A(new_n624), .B(KEYINPUT80), .Z(G280));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n618), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n547), .A2(new_n622), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n617), .A2(G559), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n629), .B1(new_n630), .B2(new_n622), .ZN(G323));
  XNOR2_X1  g206(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g207(.A1(new_n464), .A2(new_n468), .ZN(new_n633));
  XOR2_X1   g208(.A(KEYINPUT81), .B(KEYINPUT12), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(G2100), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n483), .A2(G135), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n485), .A2(G123), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n465), .A2(G111), .ZN(new_n642));
  OAI21_X1  g217(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n643));
  OAI211_X1 g218(.A(new_n640), .B(new_n641), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(G2096), .Z(new_n645));
  NAND3_X1  g220(.A1(new_n638), .A2(new_n639), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n646), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g222(.A(KEYINPUT15), .B(G2435), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2438), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2427), .B(G2430), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  AND2_X1   g227(.A1(new_n652), .A2(KEYINPUT83), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n652), .A2(KEYINPUT83), .ZN(new_n654));
  OAI22_X1  g229(.A1(new_n653), .A2(new_n654), .B1(new_n649), .B2(new_n650), .ZN(new_n655));
  XOR2_X1   g230(.A(G2443), .B(G2446), .Z(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n655), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g233(.A(G1341), .B(G1348), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  OR2_X1    g235(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n658), .A2(new_n660), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2451), .B(G2454), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT16), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n661), .A2(new_n665), .A3(new_n662), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(G14), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(G401));
  XNOR2_X1  g245(.A(G2067), .B(G2678), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT84), .ZN(new_n672));
  NOR2_X1   g247(.A1(G2072), .A2(G2078), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n442), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2084), .B(G2090), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT18), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n672), .A2(new_n674), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n674), .B(KEYINPUT17), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n678), .B(new_n675), .C1(new_n672), .C2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n675), .ZN(new_n681));
  NAND3_X1  g256(.A1(new_n679), .A2(new_n672), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n677), .A2(new_n680), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G2100), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT85), .B(G2096), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(new_n686), .ZN(G227));
  XNOR2_X1  g262(.A(G1956), .B(G2474), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1961), .B(G1966), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1971), .B(G1976), .ZN(new_n691));
  INV_X1    g266(.A(KEYINPUT19), .ZN(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n688), .A2(new_n689), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n690), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n695), .A2(KEYINPUT86), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n696), .B1(new_n693), .B2(new_n694), .ZN(new_n700));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1991), .B(G1996), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1981), .B(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(G229));
  XNOR2_X1  g284(.A(KEYINPUT30), .B(G28), .ZN(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  OR2_X1    g286(.A1(KEYINPUT31), .A2(G11), .ZN(new_n712));
  NAND2_X1  g287(.A1(KEYINPUT31), .A2(G11), .ZN(new_n713));
  AOI22_X1  g288(.A1(new_n710), .A2(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g289(.A(G16), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n715), .A2(G21), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(new_n534), .B2(G16), .ZN(new_n717));
  INV_X1    g292(.A(G1966), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n714), .B1(new_n711), .B2(new_n644), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(G171), .A2(new_n715), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G5), .B2(new_n715), .ZN(new_n721));
  INV_X1    g296(.A(G1961), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI211_X1 g298(.A(new_n719), .B(new_n723), .C1(new_n718), .C2(new_n717), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(KEYINPUT95), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n715), .A2(G20), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT23), .Z(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G299), .B2(G16), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(G1956), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n725), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n711), .A2(G33), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n465), .A2(G103), .A3(G2104), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n732), .B(KEYINPUT25), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n464), .A2(G127), .ZN(new_n734));
  NAND2_X1  g309(.A1(G115), .A2(G2104), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n465), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  AOI211_X1 g311(.A(new_n733), .B(new_n736), .C1(G139), .C2(new_n483), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n731), .B1(new_n737), .B2(new_n711), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(G2072), .ZN(new_n739));
  AND2_X1   g314(.A1(KEYINPUT24), .A2(G34), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n711), .B1(KEYINPUT24), .B2(G34), .ZN(new_n741));
  OAI22_X1  g316(.A1(G160), .A2(new_n711), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  XOR2_X1   g317(.A(KEYINPUT94), .B(G2084), .Z(new_n743));
  NOR2_X1   g318(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n711), .A2(G32), .ZN(new_n745));
  NAND3_X1  g320(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT26), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G129), .B2(new_n485), .ZN(new_n748));
  AOI22_X1  g323(.A1(new_n483), .A2(G141), .B1(G105), .B2(new_n468), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n711), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT27), .B(G1996), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NOR3_X1   g329(.A1(new_n739), .A2(new_n744), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n711), .A2(G26), .ZN(new_n756));
  XOR2_X1   g331(.A(new_n756), .B(KEYINPUT28), .Z(new_n757));
  NAND2_X1  g332(.A1(new_n483), .A2(G140), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT92), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n758), .B(new_n759), .ZN(new_n760));
  OAI21_X1  g335(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n761));
  INV_X1    g336(.A(G116), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n761), .B1(new_n762), .B2(G2105), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT93), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n485), .A2(G128), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n760), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n757), .B1(new_n766), .B2(G29), .ZN(new_n767));
  INV_X1    g342(.A(G2067), .ZN(new_n768));
  XNOR2_X1  g343(.A(new_n767), .B(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n742), .B2(new_n743), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n755), .B(new_n770), .C1(new_n724), .C2(KEYINPUT95), .ZN(new_n771));
  NOR2_X1   g346(.A1(G29), .A2(G35), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G162), .B2(G29), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT29), .ZN(new_n774));
  XOR2_X1   g349(.A(new_n774), .B(G2090), .Z(new_n775));
  NAND2_X1  g350(.A1(new_n715), .A2(G4), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(new_n618), .B2(new_n715), .ZN(new_n777));
  INV_X1    g352(.A(G1348), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n711), .A2(G27), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G164), .B2(new_n711), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(G2078), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n721), .B2(new_n722), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n715), .A2(G19), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n548), .B2(new_n715), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1341), .Z(new_n786));
  NAND4_X1  g361(.A1(new_n775), .A2(new_n779), .A3(new_n783), .A4(new_n786), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n730), .A2(new_n771), .A3(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n711), .A2(G25), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n485), .A2(G119), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT87), .Z(new_n792));
  NOR2_X1   g367(.A1(G95), .A2(G2105), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT88), .ZN(new_n794));
  INV_X1    g369(.A(G107), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n467), .B1(new_n795), .B2(G2105), .ZN(new_n796));
  AOI22_X1  g371(.A1(G131), .A2(new_n483), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(new_n798), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n790), .B1(new_n799), .B2(new_n711), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT35), .B(G1991), .Z(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n800), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n715), .A2(G22), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G166), .B2(new_n715), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(KEYINPUT91), .ZN(new_n808));
  OR2_X1    g383(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n807), .A2(new_n808), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n715), .A2(G23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n574), .B1(new_n533), .B2(new_n575), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G49), .B2(new_n525), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n811), .B1(new_n813), .B2(new_n715), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT33), .B(G1976), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  NAND3_X1  g391(.A1(new_n809), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  INV_X1    g392(.A(new_n817), .ZN(new_n818));
  MUX2_X1   g393(.A(G6), .B(G305), .S(G16), .Z(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT90), .Z(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT32), .B(G1981), .ZN(new_n821));
  OR2_X1    g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n821), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n818), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT34), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND4_X1  g401(.A1(new_n818), .A2(new_n822), .A3(KEYINPUT34), .A4(new_n823), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n803), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n715), .A2(G24), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n829), .B1(new_n609), .B2(new_n715), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT89), .Z(new_n831));
  INV_X1    g406(.A(G1986), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n828), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n835), .A2(KEYINPUT36), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT36), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n828), .A2(new_n837), .A3(new_n833), .A4(new_n834), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n789), .B1(new_n836), .B2(new_n838), .ZN(G311));
  NAND2_X1  g414(.A1(new_n836), .A2(new_n838), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n840), .A2(new_n788), .ZN(G150));
  NAND2_X1  g416(.A1(new_n525), .A2(G55), .ZN(new_n842));
  NAND2_X1  g417(.A1(G80), .A2(G543), .ZN(new_n843));
  INV_X1    g418(.A(G67), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n582), .B2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G651), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n539), .A2(G93), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT96), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT96), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n842), .A2(new_n846), .A3(new_n850), .A4(new_n847), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n849), .A2(new_n547), .A3(new_n851), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT97), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n548), .A2(new_n848), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n852), .B2(new_n854), .ZN(new_n857));
  OAI211_X1 g432(.A(G559), .B(new_n618), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n852), .A2(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT97), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n860), .B(new_n855), .C1(new_n627), .C2(new_n617), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n862));
  AND3_X1   g437(.A1(new_n858), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n858), .B2(new_n861), .ZN(new_n864));
  OR3_X1    g439(.A1(new_n863), .A2(new_n864), .A3(KEYINPUT39), .ZN(new_n865));
  XOR2_X1   g440(.A(KEYINPUT99), .B(G860), .Z(new_n866));
  OAI21_X1  g441(.A(KEYINPUT39), .B1(new_n863), .B2(new_n864), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n849), .A2(new_n851), .ZN(new_n869));
  INV_X1    g444(.A(new_n869), .ZN(new_n870));
  NOR2_X1   g445(.A1(new_n870), .A2(new_n866), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT37), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n868), .A2(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT100), .ZN(G145));
  NAND2_X1  g449(.A1(new_n483), .A2(G142), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n485), .A2(G130), .ZN(new_n876));
  OR2_X1    g451(.A1(G106), .A2(G2105), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n877), .B(G2104), .C1(G118), .C2(new_n465), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n875), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT101), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n635), .ZN(new_n881));
  AND2_X1   g456(.A1(new_n881), .A2(new_n799), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n881), .A2(new_n799), .ZN(new_n883));
  OR3_X1    g458(.A1(new_n882), .A2(new_n883), .A3(KEYINPUT102), .ZN(new_n884));
  OAI21_X1  g459(.A(KEYINPUT102), .B1(new_n882), .B2(new_n883), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n766), .B(G164), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n886), .A2(new_n737), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n737), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n750), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n750), .B1(new_n887), .B2(new_n888), .ZN(new_n891));
  OAI211_X1 g466(.A(new_n884), .B(new_n885), .C1(new_n890), .C2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  INV_X1    g468(.A(new_n885), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n893), .A2(new_n894), .A3(new_n889), .ZN(new_n895));
  XNOR2_X1  g470(.A(G162), .B(new_n644), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G160), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n892), .B2(new_n895), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT40), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT40), .ZN(new_n905));
  NOR3_X1   g480(.A1(new_n900), .A2(new_n905), .A3(new_n902), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n904), .A2(new_n906), .ZN(G395));
  XNOR2_X1  g482(.A(G305), .B(G166), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NOR3_X1   g484(.A1(new_n606), .A2(new_n608), .A3(G288), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n599), .A2(new_n601), .A3(new_n605), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT78), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n607), .A2(KEYINPUT78), .A3(new_n601), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n813), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n909), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT104), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(G288), .B1(new_n606), .B2(new_n608), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n913), .A2(new_n813), .A3(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n921), .A2(KEYINPUT104), .A3(new_n909), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n918), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n919), .A2(new_n920), .A3(new_n908), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT105), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT105), .ZN(new_n927));
  NAND4_X1  g502(.A1(new_n919), .A2(new_n927), .A3(new_n920), .A4(new_n908), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  AND3_X1   g504(.A1(new_n923), .A2(new_n924), .A3(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT103), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(new_n617), .B2(new_n621), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n617), .A2(new_n621), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(KEYINPUT41), .ZN(new_n935));
  INV_X1    g510(.A(new_n933), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n617), .A2(new_n621), .ZN(new_n937));
  AND2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n860), .A2(new_n630), .A3(new_n855), .ZN(new_n942));
  OAI22_X1  g517(.A1(new_n856), .A2(new_n857), .B1(G559), .B2(new_n617), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n943), .A2(new_n942), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n944), .B1(new_n945), .B2(new_n934), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n924), .B1(new_n923), .B2(new_n929), .ZN(new_n947));
  NOR3_X1   g522(.A1(new_n930), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n934), .B1(new_n943), .B2(new_n942), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(new_n945), .B2(new_n941), .ZN(new_n950));
  AOI21_X1  g525(.A(KEYINPUT104), .B1(new_n921), .B2(new_n909), .ZN(new_n951));
  AOI211_X1 g526(.A(new_n917), .B(new_n908), .C1(new_n919), .C2(new_n920), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n929), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n923), .A2(new_n924), .A3(new_n929), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n950), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(G868), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n870), .A2(G868), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(G295));
  INV_X1    g535(.A(KEYINPUT106), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n961), .B1(new_n957), .B2(new_n959), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n946), .B1(new_n930), .B2(new_n947), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n954), .A2(new_n950), .A3(new_n955), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n622), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NOR3_X1   g540(.A1(new_n965), .A2(KEYINPUT106), .A3(new_n958), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n962), .A2(new_n966), .ZN(G331));
  NOR2_X1   g542(.A1(G286), .A2(G301), .ZN(new_n968));
  NOR2_X1   g543(.A1(G168), .A2(G171), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n860), .B(new_n855), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  XNOR2_X1  g545(.A(new_n534), .B(KEYINPUT75), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n969), .B1(new_n971), .B2(G171), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n972), .B1(new_n856), .B2(new_n857), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n941), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n970), .A2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n934), .ZN(new_n976));
  AOI21_X1  g551(.A(G37), .B1(new_n976), .B2(new_n953), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT107), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n953), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n970), .A2(new_n973), .A3(KEYINPUT41), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n934), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n970), .A2(new_n973), .A3(KEYINPUT41), .A4(new_n938), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n923), .A2(KEYINPUT107), .A3(new_n929), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n979), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n977), .A2(new_n985), .A3(KEYINPUT43), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n975), .A2(new_n934), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n979), .A2(new_n987), .A3(new_n984), .A4(new_n974), .ZN(new_n988));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n988), .B2(new_n977), .ZN(new_n989));
  OAI21_X1  g564(.A(KEYINPUT44), .B1(new_n986), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT43), .ZN(new_n991));
  AND3_X1   g566(.A1(new_n977), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n991), .B1(new_n988), .B2(new_n977), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n990), .B1(new_n994), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g570(.A(KEYINPUT45), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G164), .B2(G1384), .ZN(new_n997));
  INV_X1    g572(.A(new_n470), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n479), .B1(new_n478), .B2(G2105), .ZN(new_n999));
  AOI211_X1 g574(.A(KEYINPUT69), .B(new_n465), .C1(new_n477), .C2(new_n471), .ZN(new_n1000));
  OAI211_X1 g575(.A(G40), .B(new_n998), .C1(new_n999), .C2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n1002), .A2(G1996), .A3(new_n750), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT109), .ZN(new_n1004));
  XNOR2_X1  g579(.A(new_n766), .B(G2067), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n750), .A2(G1996), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1004), .B1(new_n1007), .B2(new_n1002), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n799), .A2(new_n801), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n798), .A2(new_n802), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1002), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n609), .A2(new_n832), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT108), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1015), .B1(new_n832), .B2(new_n609), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1012), .B1(new_n1016), .B2(new_n1002), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT57), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT119), .B1(G299), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT119), .ZN(new_n1020));
  NOR3_X1   g595(.A1(new_n621), .A2(new_n1020), .A3(KEYINPUT57), .ZN(new_n1021));
  AND4_X1   g596(.A1(KEYINPUT120), .A2(new_n563), .A3(KEYINPUT57), .A4(new_n569), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT120), .B1(new_n621), .B2(KEYINPUT57), .ZN(new_n1023));
  OAI22_X1  g598(.A1(new_n1019), .A2(new_n1021), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(new_n507), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n506), .B1(new_n464), .B2(new_n503), .ZN(new_n1027));
  OAI211_X1 g602(.A(new_n500), .B(new_n499), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT50), .ZN(new_n1029));
  INV_X1    g604(.A(G1384), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(new_n1001), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1032), .B1(new_n1034), .B2(KEYINPUT116), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT116), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1036), .B1(new_n1033), .B2(new_n1001), .ZN(new_n1037));
  AOI21_X1  g612(.A(G1956), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1028), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT45), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1040));
  NOR3_X1   g615(.A1(new_n1039), .A2(new_n1040), .A3(new_n1001), .ZN(new_n1041));
  XNOR2_X1  g616(.A(KEYINPUT56), .B(G2072), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1041), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1025), .B1(new_n1038), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT110), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n1031), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(KEYINPUT110), .A3(KEYINPUT50), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1001), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g626(.A1(G160), .A2(G40), .A3(new_n1030), .A4(new_n1028), .ZN(new_n1052));
  OAI22_X1  g627(.A1(new_n1051), .A2(G1348), .B1(G2067), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1045), .B1(new_n1054), .B2(new_n617), .ZN(new_n1055));
  INV_X1    g630(.A(G40), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1056), .B(new_n470), .C1(new_n474), .C2(new_n480), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(new_n1046), .A3(KEYINPUT116), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(new_n1037), .A3(new_n1031), .ZN(new_n1059));
  INV_X1    g634(.A(G1956), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1061), .A2(new_n1043), .A3(new_n1024), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1055), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT59), .ZN(new_n1064));
  INV_X1    g639(.A(G1996), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1028), .A2(KEYINPUT45), .A3(new_n1030), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1057), .A2(new_n997), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  XOR2_X1   g642(.A(KEYINPUT58), .B(G1341), .Z(new_n1068));
  AOI22_X1  g643(.A1(new_n1067), .A2(KEYINPUT121), .B1(new_n1052), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT121), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(new_n1065), .A4(new_n1057), .ZN(new_n1072));
  AOI211_X1 g647(.A(new_n1064), .B(new_n547), .C1(new_n1069), .C2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1067), .A2(KEYINPUT121), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1052), .A2(new_n1068), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1072), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  AOI21_X1  g651(.A(KEYINPUT59), .B1(new_n1076), .B2(new_n548), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1073), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT61), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1024), .A2(new_n1043), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n1080), .A2(new_n1038), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1024), .B1(new_n1061), .B2(new_n1043), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1045), .A2(KEYINPUT61), .A3(new_n1062), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1078), .A2(new_n1083), .A3(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1054), .A2(KEYINPUT60), .A3(new_n617), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT60), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n618), .B1(new_n1053), .B2(new_n1087), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1086), .A2(new_n1088), .B1(new_n1087), .B2(new_n1053), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1063), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  INV_X1    g666(.A(G8), .ZN(new_n1092));
  NOR2_X1   g667(.A1(G168), .A2(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT122), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1091), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g670(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT117), .B(G2084), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n1001), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(G1966), .B2(new_n1041), .ZN(new_n1101));
  OAI211_X1 g676(.A(G8), .B(new_n1096), .C1(new_n1101), .C2(new_n534), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1093), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1093), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1057), .A2(new_n997), .A3(new_n1066), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1097), .A2(new_n1099), .B1(new_n718), .B2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1104), .B(new_n1095), .C1(new_n1106), .C2(new_n1092), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1102), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT123), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1102), .A2(KEYINPUT123), .A3(new_n1103), .A4(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1070), .A2(KEYINPUT53), .A3(new_n1113), .A4(new_n1057), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1057), .A2(new_n997), .A3(new_n1113), .A4(new_n1066), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT53), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  XOR2_X1   g692(.A(KEYINPUT124), .B(G1961), .Z(new_n1118));
  OAI211_X1 g693(.A(new_n1114), .B(new_n1117), .C1(new_n1051), .C2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT54), .B1(new_n1119), .B2(G171), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1113), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1121));
  AOI211_X1 g696(.A(new_n1121), .B(new_n470), .C1(G2105), .C2(new_n478), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1115), .A2(new_n1116), .B1(new_n1070), .B2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1051), .B2(new_n1118), .ZN(new_n1124));
  AOI21_X1  g699(.A(G301), .B1(new_n1124), .B2(KEYINPUT125), .ZN(new_n1125));
  OR2_X1    g700(.A1(new_n1051), .A2(new_n1118), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT125), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1126), .A2(new_n1127), .A3(new_n1123), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1120), .B1(new_n1125), .B2(new_n1128), .ZN(new_n1129));
  XOR2_X1   g704(.A(KEYINPUT111), .B(G2090), .Z(new_n1130));
  NAND3_X1  g705(.A1(new_n1097), .A2(new_n1057), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT112), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1105), .A2(new_n806), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1131), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1057), .A2(new_n1130), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1135), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1136));
  AOI21_X1  g711(.A(G1971), .B1(new_n1070), .B2(new_n1057), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT112), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(G303), .A2(G8), .ZN(new_n1139));
  XNOR2_X1  g714(.A(new_n1139), .B(KEYINPUT55), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1134), .A2(new_n1138), .A3(G8), .A4(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n813), .A2(G1976), .ZN(new_n1143));
  INV_X1    g718(.A(G1976), .ZN(new_n1144));
  AOI21_X1  g719(.A(KEYINPUT52), .B1(G288), .B2(new_n1144), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n1052), .A2(G8), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT113), .ZN(new_n1147));
  XNOR2_X1  g722(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1052), .A2(G8), .A3(new_n1143), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT52), .ZN(new_n1150));
  INV_X1    g725(.A(G1981), .ZN(new_n1151));
  XNOR2_X1  g726(.A(KEYINPUT115), .B(G86), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n539), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1151), .B1(new_n586), .B2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n583), .B1(new_n592), .B2(new_n579), .ZN(new_n1155));
  INV_X1    g730(.A(new_n578), .ZN(new_n1156));
  OAI21_X1  g731(.A(G651), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n532), .A2(new_n585), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1157), .A2(new_n1151), .A3(new_n587), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT114), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT114), .ZN(new_n1161));
  NAND4_X1  g736(.A1(new_n586), .A2(new_n1161), .A3(new_n1151), .A4(new_n587), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1154), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(G8), .B(new_n1052), .C1(new_n1163), .C2(KEYINPUT49), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT49), .ZN(new_n1165));
  AOI211_X1 g740(.A(new_n1165), .B(new_n1154), .C1(new_n1160), .C2(new_n1162), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1150), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1148), .A2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1058), .A2(new_n1037), .A3(new_n1031), .A4(new_n1130), .ZN(new_n1169));
  AND2_X1   g744(.A1(new_n1169), .A2(new_n1133), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1140), .B1(new_n1170), .B2(new_n1092), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1142), .A2(new_n1168), .A3(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1126), .A2(G301), .A3(new_n1123), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1119), .A2(G171), .ZN(new_n1174));
  AOI21_X1  g749(.A(KEYINPUT54), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NOR3_X1   g750(.A1(new_n1129), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1090), .A2(new_n1112), .A3(new_n1176), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1134), .A2(G8), .A3(new_n1138), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1178), .A2(new_n1140), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1100), .ZN(new_n1180));
  NOR2_X1   g755(.A1(new_n1041), .A2(G1966), .ZN(new_n1181));
  OAI211_X1 g756(.A(G8), .B(new_n971), .C1(new_n1180), .C2(new_n1181), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT63), .ZN(new_n1183));
  NOR2_X1   g758(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1179), .A2(new_n1184), .A3(new_n1142), .A4(new_n1168), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1185), .A2(KEYINPUT118), .ZN(new_n1186));
  AND2_X1   g761(.A1(new_n1142), .A2(new_n1168), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT118), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1187), .A2(new_n1188), .A3(new_n1179), .A4(new_n1184), .ZN(new_n1189));
  OAI21_X1  g764(.A(new_n1183), .B1(new_n1172), .B2(new_n1182), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1186), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1052), .A2(G8), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1144), .B(new_n813), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1162), .A2(new_n1160), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1192), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1142), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1195), .B1(new_n1196), .B2(new_n1168), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1177), .A2(new_n1191), .A3(new_n1197), .ZN(new_n1198));
  OR2_X1    g773(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT62), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1112), .A2(new_n1200), .ZN(new_n1201));
  NAND3_X1  g776(.A1(new_n1110), .A2(KEYINPUT62), .A3(new_n1111), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n1199), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1017), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g779(.A(KEYINPUT46), .B1(new_n1002), .B2(new_n1065), .ZN(new_n1205));
  XNOR2_X1  g780(.A(new_n1205), .B(KEYINPUT126), .ZN(new_n1206));
  AOI211_X1 g781(.A(new_n750), .B(new_n1005), .C1(KEYINPUT46), .C2(new_n1065), .ZN(new_n1207));
  INV_X1    g782(.A(new_n1002), .ZN(new_n1208));
  OAI21_X1  g783(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT47), .Z(new_n1210));
  INV_X1    g785(.A(KEYINPUT48), .ZN(new_n1211));
  NOR3_X1   g786(.A1(new_n1015), .A2(new_n1211), .A3(new_n1208), .ZN(new_n1212));
  AOI21_X1  g787(.A(KEYINPUT48), .B1(new_n1014), .B2(new_n1002), .ZN(new_n1213));
  NOR3_X1   g788(.A1(new_n1212), .A2(new_n1012), .A3(new_n1213), .ZN(new_n1214));
  NOR2_X1   g789(.A1(new_n766), .A2(G2067), .ZN(new_n1215));
  AOI21_X1  g790(.A(new_n1215), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1216));
  NOR2_X1   g791(.A1(new_n1216), .A2(new_n1208), .ZN(new_n1217));
  NOR3_X1   g792(.A1(new_n1210), .A2(new_n1214), .A3(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1204), .A2(new_n1218), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g794(.A1(new_n686), .A2(G319), .ZN(new_n1221));
  NOR2_X1   g795(.A1(G229), .A2(new_n1221), .ZN(new_n1222));
  OAI211_X1 g796(.A(new_n1222), .B(new_n669), .C1(new_n900), .C2(new_n902), .ZN(new_n1223));
  NOR2_X1   g797(.A1(new_n1223), .A2(new_n994), .ZN(G308));
  NOR3_X1   g798(.A1(G401), .A2(G229), .A3(new_n1221), .ZN(new_n1225));
  OAI221_X1 g799(.A(new_n1225), .B1(new_n902), .B2(new_n900), .C1(new_n993), .C2(new_n992), .ZN(G225));
endmodule


