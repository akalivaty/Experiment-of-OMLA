//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n768, new_n769, new_n770,
    new_n772, new_n773, new_n774, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n878, new_n879, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n957, new_n958, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1014,
    new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT101), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n203), .A2(G1gat), .ZN(new_n207));
  OAI21_X1  g006(.A(G8gat), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n203), .A2(new_n205), .ZN(new_n209));
  INV_X1    g008(.A(G8gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n209), .B(new_n210), .C1(G1gat), .C2(new_n203), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT21), .ZN(new_n214));
  XNOR2_X1  g013(.A(G71gat), .B(G78gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G71gat), .A2(G78gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT9), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G64gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(G57gat), .ZN(new_n222));
  INV_X1    g021(.A(G57gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(new_n223), .A2(G64gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n220), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n226), .A2(new_n218), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n216), .B1(new_n225), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g027(.A1(new_n226), .A2(new_n218), .ZN(new_n229));
  XOR2_X1   g028(.A(G57gat), .B(G64gat), .Z(new_n230));
  NAND4_X1  g029(.A1(new_n229), .A2(new_n230), .A3(new_n215), .A4(new_n220), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n213), .B1(new_n214), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(KEYINPUT96), .B(KEYINPUT97), .Z(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n237));
  AND2_X1   g036(.A1(new_n228), .A2(new_n231), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n237), .B1(new_n238), .B2(KEYINPUT21), .ZN(new_n239));
  NAND2_X1  g038(.A1(G231gat), .A2(G233gat), .ZN(new_n240));
  XOR2_X1   g039(.A(new_n240), .B(KEYINPUT95), .Z(new_n241));
  INV_X1    g040(.A(new_n237), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n232), .A2(new_n214), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n239), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G155gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n241), .ZN(new_n247));
  AOI21_X1  g046(.A(new_n242), .B1(new_n232), .B2(new_n214), .ZN(new_n248));
  AOI211_X1 g047(.A(KEYINPUT21), .B(new_n237), .C1(new_n228), .C2(new_n231), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n244), .A2(new_n246), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n246), .B1(new_n244), .B2(new_n250), .ZN(new_n253));
  XOR2_X1   g052(.A(G183gat), .B(G211gat), .Z(new_n254));
  NOR3_X1   g053(.A1(new_n252), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(new_n254), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n244), .A2(new_n250), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(new_n245), .ZN(new_n258));
  AOI21_X1  g057(.A(new_n256), .B1(new_n258), .B2(new_n251), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n236), .B1(new_n255), .B2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n254), .B1(new_n252), .B2(new_n253), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(new_n256), .A3(new_n251), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n261), .A2(new_n262), .A3(new_n235), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g063(.A1(G232gat), .A2(G233gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n265), .A2(KEYINPUT41), .ZN(new_n266));
  XNOR2_X1  g065(.A(G134gat), .B(G162gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(G99gat), .A2(G106gat), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT98), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(G99gat), .A3(G106gat), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n273), .A3(KEYINPUT8), .ZN(new_n274));
  OR2_X1    g073(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n275));
  INV_X1    g074(.A(G92gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(KEYINPUT99), .A2(G85gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n275), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(G85gat), .A2(G92gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT7), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT7), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(G85gat), .A3(G92gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n274), .A2(new_n278), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g083(.A1(G99gat), .A2(G106gat), .ZN(new_n285));
  NOR2_X1   g084(.A1(G99gat), .A2(G106gat), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n284), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n289), .A2(new_n274), .A3(new_n278), .A4(new_n283), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT100), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n288), .A2(new_n290), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT100), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G43gat), .B(G50gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT15), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT89), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT14), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n300), .B(new_n301), .C1(G29gat), .C2(G36gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(G29gat), .A2(G36gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n302), .B(new_n303), .C1(new_n297), .C2(KEYINPUT15), .ZN(new_n304));
  INV_X1    g103(.A(G29gat), .ZN(new_n305));
  INV_X1    g104(.A(G36gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n305), .A2(new_n306), .A3(KEYINPUT89), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n300), .B1(G29gat), .B2(G36gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT14), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n299), .B1(new_n304), .B2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G50gat), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G43gat), .ZN(new_n313));
  INV_X1    g112(.A(G43gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(G50gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT15), .ZN(new_n317));
  AOI22_X1  g116(.A1(new_n316), .A2(new_n317), .B1(G29gat), .B2(G36gat), .ZN(new_n318));
  NAND4_X1  g117(.A1(new_n318), .A2(new_n298), .A3(new_n309), .A4(new_n302), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n311), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n296), .A2(new_n320), .B1(KEYINPUT41), .B2(new_n265), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT17), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n311), .A2(new_n319), .A3(KEYINPUT17), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n292), .A2(new_n323), .A3(new_n324), .A4(new_n295), .ZN(new_n325));
  XOR2_X1   g124(.A(G190gat), .B(G218gat), .Z(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n321), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n327), .B1(new_n321), .B2(new_n325), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n269), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n330), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n332), .A2(new_n268), .A3(new_n328), .ZN(new_n333));
  AND2_X1   g132(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n202), .B1(new_n264), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n260), .A2(new_n263), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n331), .A2(new_n333), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n336), .A2(new_n337), .A3(KEYINPUT101), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G120gat), .B(G148gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n291), .A2(new_n238), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT103), .ZN(new_n345));
  AND3_X1   g144(.A1(new_n274), .A2(new_n278), .A3(new_n283), .ZN(new_n346));
  OR2_X1    g145(.A1(G99gat), .A2(G106gat), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT102), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n347), .A2(new_n348), .A3(new_n270), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT102), .B1(new_n285), .B2(new_n286), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n345), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n349), .A2(new_n350), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(new_n284), .A3(KEYINPUT103), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n228), .A2(new_n290), .A3(new_n231), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT104), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(new_n356), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT104), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n352), .A4(new_n354), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n344), .B1(new_n357), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT105), .ZN(new_n363));
  NAND2_X1  g162(.A1(G230gat), .A2(G233gat), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n362), .A2(new_n363), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g165(.A(KEYINPUT105), .B1(new_n361), .B2(new_n364), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n369));
  INV_X1    g168(.A(new_n344), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n353), .A2(new_n284), .A3(KEYINPUT103), .ZN(new_n371));
  AOI21_X1  g170(.A(KEYINPUT103), .B1(new_n353), .B2(new_n284), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n359), .B1(new_n373), .B2(new_n358), .ZN(new_n374));
  NOR4_X1   g173(.A1(new_n356), .A2(new_n371), .A3(new_n372), .A4(KEYINPUT104), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n369), .B(new_n370), .C1(new_n374), .C2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n232), .A2(new_n369), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n296), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n365), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n343), .B1(new_n368), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g179(.A(KEYINPUT10), .B(new_n344), .C1(new_n357), .C2(new_n360), .ZN(new_n381));
  AND2_X1   g180(.A1(new_n296), .A2(new_n377), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n364), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  NAND4_X1  g182(.A1(new_n383), .A2(new_n366), .A3(new_n342), .A4(new_n367), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NOR2_X1   g184(.A1(new_n339), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT64), .ZN(new_n388));
  NOR2_X1   g187(.A1(G169gat), .A2(G176gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n388), .B1(new_n389), .B2(KEYINPUT23), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT23), .ZN(new_n391));
  OAI211_X1 g190(.A(new_n391), .B(KEYINPUT64), .C1(G169gat), .C2(G176gat), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n390), .A2(new_n392), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n389), .B(KEYINPUT65), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n393), .B1(new_n391), .B2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(G183gat), .A2(G190gat), .ZN(new_n396));
  AOI21_X1  g195(.A(KEYINPUT24), .B1(new_n396), .B2(KEYINPUT66), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(KEYINPUT66), .B2(new_n396), .ZN(new_n398));
  NAND3_X1  g197(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(G183gat), .B2(G190gat), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT67), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n399), .A2(KEYINPUT67), .ZN(new_n403));
  AND3_X1   g202(.A1(new_n398), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT25), .B1(new_n395), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(KEYINPUT25), .B1(new_n389), .B2(KEYINPUT23), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n407));
  OAI211_X1 g206(.A(new_n393), .B(new_n406), .C1(new_n400), .C2(new_n407), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n410));
  INV_X1    g209(.A(G169gat), .ZN(new_n411));
  INV_X1    g210(.A(G176gat), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n410), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(KEYINPUT70), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n414), .B(new_n415), .C1(KEYINPUT26), .C2(new_n394), .ZN(new_n416));
  XNOR2_X1  g215(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n417));
  XOR2_X1   g216(.A(KEYINPUT27), .B(G183gat), .Z(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n419), .A2(KEYINPUT68), .ZN(new_n420));
  INV_X1    g219(.A(G183gat), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n421), .A2(KEYINPUT27), .ZN(new_n422));
  AOI21_X1  g221(.A(G190gat), .B1(new_n422), .B2(KEYINPUT68), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n417), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(G190gat), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n419), .A2(KEYINPUT28), .A3(new_n425), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n396), .B(new_n416), .C1(new_n424), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g227(.A(G127gat), .B(G134gat), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT71), .ZN(new_n430));
  INV_X1    g229(.A(G113gat), .ZN(new_n431));
  INV_X1    g230(.A(G120gat), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT1), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n433), .B1(new_n431), .B2(new_n432), .ZN(new_n434));
  INV_X1    g233(.A(G127gat), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(G134gat), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n430), .B(new_n434), .C1(KEYINPUT71), .C2(new_n436), .ZN(new_n437));
  XOR2_X1   g236(.A(KEYINPUT72), .B(G120gat), .Z(new_n438));
  OAI211_X1 g237(.A(new_n433), .B(new_n429), .C1(new_n438), .C2(new_n431), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n428), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(G227gat), .ZN(new_n442));
  INV_X1    g241(.A(G233gat), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n437), .A2(new_n439), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n409), .A2(new_n427), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n441), .A2(new_n444), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT32), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G15gat), .B(G43gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n453), .ZN(new_n455));
  OAI211_X1 g254(.A(new_n447), .B(KEYINPUT32), .C1(new_n449), .C2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n454), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT34), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n446), .ZN(new_n459));
  INV_X1    g258(.A(new_n444), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n461), .ZN(new_n462));
  AOI211_X1 g261(.A(KEYINPUT34), .B(new_n444), .C1(new_n441), .C2(new_n446), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n464), .A3(KEYINPUT74), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT74), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n466), .B1(new_n461), .B2(new_n463), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n457), .A2(new_n465), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n462), .A2(new_n464), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n469), .A2(new_n466), .A3(new_n454), .A4(new_n456), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G228gat), .A2(G233gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n472), .B(G22gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(KEYINPUT31), .B(G50gat), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n473), .B(new_n474), .Z(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT3), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT22), .ZN(new_n478));
  AOI22_X1  g277(.A1(new_n478), .A2(KEYINPUT75), .B1(G211gat), .B2(G218gat), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(KEYINPUT75), .B2(new_n478), .ZN(new_n480));
  XNOR2_X1  g279(.A(G197gat), .B(G204gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT76), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n482), .B(new_n483), .ZN(new_n484));
  XOR2_X1   g283(.A(G211gat), .B(G218gat), .Z(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n484), .B(new_n486), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n477), .B1(new_n487), .B2(KEYINPUT29), .ZN(new_n488));
  XOR2_X1   g287(.A(G141gat), .B(G148gat), .Z(new_n489));
  INV_X1    g288(.A(G155gat), .ZN(new_n490));
  INV_X1    g289(.A(G162gat), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT2), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  XOR2_X1   g292(.A(G155gat), .B(G162gat), .Z(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n488), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(new_n494), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n493), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n477), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT29), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n487), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G78gat), .B(G106gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n496), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n504), .B1(new_n496), .B2(new_n502), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n476), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n507), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n509), .A2(new_n505), .A3(new_n475), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  XOR2_X1   g311(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n513));
  NAND3_X1  g312(.A1(new_n471), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT87), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n440), .A2(new_n498), .ZN(new_n517));
  AOI21_X1  g316(.A(KEYINPUT81), .B1(new_n517), .B2(KEYINPUT4), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n495), .A2(new_n445), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT4), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n518), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(G225gat), .A2(G233gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT80), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n495), .A2(KEYINPUT3), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n499), .A2(new_n526), .A3(new_n445), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n519), .A2(KEYINPUT81), .A3(new_n520), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n522), .A2(new_n525), .A3(new_n527), .A4(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT5), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n495), .A2(new_n445), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n517), .A2(new_n531), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n532), .B2(new_n524), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT83), .B1(new_n517), .B2(KEYINPUT4), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT83), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n535), .A3(new_n520), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n517), .A2(KEYINPUT84), .A3(KEYINPUT4), .ZN(new_n537));
  AOI21_X1  g336(.A(KEYINPUT84), .B1(new_n517), .B2(KEYINPUT4), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n534), .B(new_n536), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n527), .A2(new_n530), .A3(new_n525), .ZN(new_n540));
  AOI22_X1  g339(.A1(new_n529), .A2(new_n533), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  XOR2_X1   g340(.A(G1gat), .B(G29gat), .Z(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(G57gat), .B(G85gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n541), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT85), .B1(new_n547), .B2(KEYINPUT6), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT6), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n541), .A2(new_n550), .A3(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n529), .A2(new_n533), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n539), .A2(new_n540), .ZN(new_n553));
  AND3_X1   g352(.A1(new_n552), .A2(new_n546), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n553), .ZN(new_n556));
  INV_X1    g355(.A(new_n546), .ZN(new_n557));
  AOI21_X1  g356(.A(KEYINPUT6), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n551), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT85), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n549), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(G226gat), .A2(G233gat), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n563), .B1(new_n428), .B2(new_n500), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n562), .B1(new_n409), .B2(new_n427), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n487), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n428), .A2(new_n563), .ZN(new_n567));
  INV_X1    g366(.A(new_n487), .ZN(new_n568));
  AOI21_X1  g367(.A(KEYINPUT29), .B1(new_n409), .B2(new_n427), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n567), .B(new_n568), .C1(new_n563), .C2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G8gat), .B(G36gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(G64gat), .B(G92gat), .ZN(new_n572));
  XOR2_X1   g371(.A(new_n571), .B(new_n572), .Z(new_n573));
  NAND3_X1  g372(.A1(new_n566), .A2(new_n570), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT78), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT78), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n566), .A2(new_n576), .A3(new_n570), .A4(new_n573), .ZN(new_n577));
  XNOR2_X1  g376(.A(KEYINPUT79), .B(KEYINPUT30), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n566), .A2(KEYINPUT30), .A3(new_n570), .A4(new_n573), .ZN(new_n580));
  INV_X1    g379(.A(new_n573), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n570), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT77), .B1(new_n566), .B2(new_n570), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n581), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g383(.A1(new_n579), .A2(new_n580), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n516), .B1(new_n561), .B2(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n556), .A2(KEYINPUT6), .A3(new_n557), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n550), .B1(new_n541), .B2(new_n546), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n587), .B1(new_n588), .B2(new_n554), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n548), .B1(new_n589), .B2(KEYINPUT85), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n579), .A2(new_n584), .A3(new_n580), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT87), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n515), .B1(new_n586), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT35), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT73), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n457), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n469), .ZN(new_n597));
  NAND4_X1  g396(.A1(new_n457), .A2(new_n595), .A3(new_n462), .A4(new_n464), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n511), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND4_X1  g398(.A1(new_n579), .A2(new_n589), .A3(new_n584), .A4(new_n580), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n594), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n525), .B1(new_n539), .B2(new_n527), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT39), .B1(new_n532), .B2(new_n524), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT39), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n557), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n606), .A2(new_n608), .A3(KEYINPUT40), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT40), .B1(new_n606), .B2(new_n608), .ZN(new_n610));
  NOR3_X1   g409(.A1(new_n609), .A2(new_n610), .A3(new_n547), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n511), .B1(new_n611), .B2(new_n591), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n575), .A2(new_n577), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT37), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n566), .A2(new_n614), .A3(new_n570), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(new_n581), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n566), .A2(new_n570), .ZN(new_n618));
  AOI21_X1  g417(.A(KEYINPUT38), .B1(new_n618), .B2(KEYINPUT37), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n613), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT38), .ZN(new_n621));
  OAI21_X1  g420(.A(KEYINPUT37), .B1(new_n582), .B2(new_n583), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n621), .B1(new_n622), .B2(new_n617), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n620), .B(new_n590), .C1(new_n623), .C2(KEYINPUT86), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT77), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n618), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n566), .A2(KEYINPUT77), .A3(new_n570), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n614), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  OAI21_X1  g427(.A(KEYINPUT38), .B1(new_n628), .B2(new_n616), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT86), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n612), .B1(new_n624), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n600), .A2(new_n511), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n471), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n597), .A2(KEYINPUT36), .A3(new_n598), .ZN(new_n636));
  AND3_X1   g435(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  AOI22_X1  g436(.A1(new_n593), .A2(new_n603), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT90), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n323), .A2(new_n639), .A3(new_n213), .A4(new_n324), .ZN(new_n640));
  AND3_X1   g439(.A1(new_n311), .A2(new_n319), .A3(KEYINPUT17), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT17), .B1(new_n311), .B2(new_n319), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n641), .A2(new_n642), .A3(new_n212), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n639), .B1(new_n320), .B2(new_n212), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n640), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G229gat), .A2(G233gat), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT18), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n647), .B(KEYINPUT13), .Z(new_n650));
  OAI21_X1  g449(.A(KEYINPUT92), .B1(new_n320), .B2(new_n212), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n320), .A2(new_n212), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n651), .B(new_n652), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n648), .A2(new_n649), .B1(new_n650), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G113gat), .B(G141gat), .ZN(new_n655));
  INV_X1    g454(.A(G197gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g456(.A(KEYINPUT11), .B(G169gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT12), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n646), .A2(KEYINPUT18), .A3(new_n647), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT91), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n647), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n323), .A2(new_n213), .A3(new_n324), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n644), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n666), .B2(new_n640), .ZN(new_n667));
  AOI21_X1  g466(.A(KEYINPUT91), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n654), .B(new_n660), .C1(new_n663), .C2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n661), .A2(new_n662), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n667), .A2(KEYINPUT91), .A3(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n660), .B1(new_n673), .B2(new_n654), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT93), .B1(new_n638), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT93), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n654), .B1(new_n663), .B2(new_n668), .ZN(new_n678));
  INV_X1    g477(.A(new_n660), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(new_n669), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n561), .A2(new_n585), .A3(new_n516), .ZN(new_n682));
  OAI21_X1  g481(.A(KEYINPUT87), .B1(new_n590), .B2(new_n591), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n514), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n602), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n629), .A2(new_n630), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n687), .A2(new_n688), .A3(new_n590), .A4(new_n620), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n686), .B1(new_n689), .B2(new_n612), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n677), .B(new_n681), .C1(new_n685), .C2(new_n690), .ZN(new_n691));
  AOI21_X1  g490(.A(new_n387), .B1(new_n676), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n559), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT106), .B(G1gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1324gat));
  NAND2_X1  g494(.A1(new_n676), .A2(new_n691), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  AND4_X1   g496(.A1(new_n591), .A2(new_n696), .A3(new_n386), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n210), .B1(new_n692), .B2(new_n591), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n692), .A2(new_n591), .A3(new_n697), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(G1325gat));
  INV_X1    g503(.A(new_n692), .ZN(new_n705));
  INV_X1    g504(.A(new_n471), .ZN(new_n706));
  OR3_X1    g505(.A1(new_n705), .A2(G15gat), .A3(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n635), .A2(new_n636), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G15gat), .B1(new_n705), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n707), .A2(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n692), .A2(new_n511), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(KEYINPUT45), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n385), .A2(new_n336), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n717), .A2(new_n337), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n696), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n589), .A2(G29gat), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n715), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n696), .A2(KEYINPUT45), .A3(new_n718), .A4(new_n720), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(new_n638), .B2(new_n337), .ZN(new_n725));
  OAI211_X1 g524(.A(KEYINPUT44), .B(new_n334), .C1(new_n685), .C2(new_n690), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n717), .A2(new_n675), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n725), .A2(new_n559), .A3(new_n726), .A4(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n730), .A2(G29gat), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n728), .A2(new_n729), .ZN(new_n732));
  OAI211_X1 g531(.A(new_n722), .B(new_n723), .C1(new_n731), .C2(new_n732), .ZN(G1328gat));
  NAND2_X1  g532(.A1(new_n591), .A2(new_n306), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n719), .A2(KEYINPUT46), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n725), .A2(new_n726), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(new_n591), .A3(new_n727), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(G36gat), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT46), .B1(new_n719), .B2(new_n734), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n735), .A2(new_n738), .A3(new_n739), .ZN(G1329gat));
  NOR2_X1   g539(.A1(new_n706), .A2(G43gat), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n696), .A2(new_n718), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT47), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n725), .A2(new_n708), .A3(new_n726), .A4(new_n727), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G43gat), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n744), .A2(new_n747), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n746), .B(new_n742), .C1(new_n743), .C2(KEYINPUT47), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1330gat));
  NOR2_X1   g549(.A1(new_n512), .A2(G50gat), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n696), .A2(new_n718), .A3(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT109), .ZN(new_n753));
  AOI21_X1  g552(.A(KEYINPUT48), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n725), .A2(new_n511), .A3(new_n726), .A4(new_n727), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(G50gat), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(new_n752), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n756), .B(new_n752), .C1(new_n753), .C2(KEYINPUT48), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(G1331gat));
  NAND2_X1  g559(.A1(new_n632), .A2(new_n637), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n602), .B2(new_n684), .ZN(new_n762));
  INV_X1    g561(.A(new_n385), .ZN(new_n763));
  NOR3_X1   g562(.A1(new_n339), .A2(new_n681), .A3(new_n763), .ZN(new_n764));
  AND2_X1   g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n559), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n591), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n769));
  XOR2_X1   g568(.A(KEYINPUT49), .B(G64gat), .Z(new_n770));
  OAI21_X1  g569(.A(new_n769), .B1(new_n768), .B2(new_n770), .ZN(G1333gat));
  NAND3_X1  g570(.A1(new_n762), .A2(new_n471), .A3(new_n764), .ZN(new_n772));
  INV_X1    g571(.A(G71gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n709), .A2(new_n773), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n762), .A2(new_n764), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n780), .B(new_n781), .ZN(G1334gat));
  NAND2_X1  g581(.A1(new_n765), .A2(new_n511), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g583(.A1(new_n275), .A2(new_n277), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n589), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n675), .A2(new_n264), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT112), .ZN(new_n788));
  OAI211_X1 g587(.A(new_n334), .B(new_n788), .C1(new_n685), .C2(new_n690), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n789), .A2(new_n790), .ZN(new_n792));
  OAI211_X1 g591(.A(new_n385), .B(new_n786), .C1(new_n791), .C2(new_n792), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n788), .A2(new_n385), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n725), .A2(new_n559), .A3(new_n726), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(KEYINPUT113), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n796), .A2(new_n785), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n795), .A2(KEYINPUT113), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n793), .B1(new_n797), .B2(new_n798), .ZN(G1336gat));
  NOR3_X1   g598(.A1(new_n585), .A2(G92gat), .A3(new_n763), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n791), .B2(new_n792), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n725), .A2(new_n591), .A3(new_n726), .A4(new_n794), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  XNOR2_X1  g602(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n801), .A2(new_n803), .A3(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT114), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n789), .A2(new_n806), .A3(KEYINPUT51), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT51), .B1(new_n789), .B2(new_n806), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI22_X1  g608(.A1(new_n809), .A2(new_n800), .B1(G92gat), .B2(new_n802), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n805), .B1(new_n810), .B2(new_n811), .ZN(G1337gat));
  NAND3_X1  g611(.A1(new_n736), .A2(new_n708), .A3(new_n794), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n813), .A2(G99gat), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n706), .A2(G99gat), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n385), .B(new_n815), .C1(new_n791), .C2(new_n792), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n814), .A2(new_n816), .ZN(G1338gat));
  NOR3_X1   g616(.A1(new_n512), .A2(G106gat), .A3(new_n763), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n791), .B2(new_n792), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n725), .A2(new_n511), .A3(new_n726), .A4(new_n794), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(G106gat), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT53), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n819), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  XOR2_X1   g622(.A(new_n818), .B(KEYINPUT116), .Z(new_n824));
  AOI22_X1  g623(.A1(new_n809), .A2(new_n824), .B1(G106gat), .B2(new_n820), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n823), .B1(new_n825), .B2(new_n822), .ZN(G1339gat));
  OAI22_X1  g625(.A1(new_n650), .A2(new_n653), .B1(new_n646), .B2(new_n647), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n659), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n385), .A2(new_n669), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n830), .B(new_n364), .C1(new_n381), .C2(new_n382), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n378), .A2(new_n365), .ZN(new_n832));
  OAI21_X1  g631(.A(KEYINPUT54), .B1(new_n381), .B2(new_n832), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n831), .B(new_n343), .C1(new_n833), .C2(new_n379), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT55), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n376), .A2(new_n378), .A3(new_n365), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n382), .B1(new_n361), .B2(new_n369), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n837), .B(KEYINPUT54), .C1(new_n838), .C2(new_n365), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n342), .B1(new_n379), .B2(new_n830), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n840), .A3(KEYINPUT55), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n836), .A2(new_n384), .A3(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n829), .B1(new_n675), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n337), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT55), .B1(new_n833), .B2(new_n379), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n831), .A2(new_n343), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n384), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(KEYINPUT55), .B1(new_n839), .B2(new_n840), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n653), .A2(new_n650), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n850), .B1(new_n667), .B2(KEYINPUT18), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n851), .B1(new_n671), .B2(new_n672), .ZN(new_n852));
  AOI22_X1  g651(.A1(new_n852), .A2(new_n660), .B1(new_n659), .B2(new_n827), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(new_n334), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n844), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(new_n338), .ZN(new_n856));
  AOI21_X1  g655(.A(KEYINPUT101), .B1(new_n336), .B2(new_n337), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT117), .ZN(new_n859));
  NAND4_X1  g658(.A1(new_n858), .A2(new_n859), .A3(new_n675), .A4(new_n763), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n335), .A2(new_n675), .A3(new_n338), .A4(new_n763), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n855), .A2(new_n264), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n863), .A2(new_n511), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n591), .A2(new_n589), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n864), .A2(new_n471), .A3(new_n865), .ZN(new_n866));
  NOR3_X1   g665(.A1(new_n866), .A2(new_n431), .A3(new_n675), .ZN(new_n867));
  INV_X1    g666(.A(new_n599), .ZN(new_n868));
  NOR4_X1   g667(.A1(new_n863), .A2(new_n589), .A3(new_n591), .A4(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(G113gat), .B1(new_n869), .B2(new_n681), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n867), .A2(new_n870), .ZN(G1340gat));
  NAND3_X1  g670(.A1(new_n869), .A2(new_n438), .A3(new_n385), .ZN(new_n872));
  OAI21_X1  g671(.A(G120gat), .B1(new_n866), .B2(new_n763), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT118), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1341gat));
  OAI21_X1  g676(.A(G127gat), .B1(new_n866), .B2(new_n264), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n869), .A2(new_n435), .A3(new_n336), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(G1342gat));
  INV_X1    g679(.A(G134gat), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n869), .A2(new_n881), .A3(new_n334), .ZN(new_n882));
  OR2_X1    g681(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n866), .B2(new_n337), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n882), .A2(KEYINPUT56), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  NAND2_X1  g685(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT122), .Z(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n860), .A2(new_n862), .ZN(new_n890));
  INV_X1    g689(.A(new_n854), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n891), .B1(new_n337), .B2(new_n843), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n890), .B1(new_n892), .B2(new_n336), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n708), .A2(new_n591), .A3(new_n512), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n893), .A2(new_n559), .A3(new_n681), .A4(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(G141gat), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g696(.A1(KEYINPUT121), .A2(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n709), .A2(new_n865), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n512), .A2(new_n902), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n849), .A2(new_n681), .B1(new_n853), .B2(new_n385), .ZN(new_n904));
  OAI21_X1  g703(.A(KEYINPUT119), .B1(new_n904), .B2(new_n334), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n843), .A2(new_n906), .A3(new_n337), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n905), .A2(new_n907), .A3(new_n854), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n908), .A2(new_n909), .A3(new_n264), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(new_n890), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n909), .B1(new_n908), .B2(new_n264), .ZN(new_n912));
  OAI21_X1  g711(.A(new_n903), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n893), .B2(new_n511), .ZN(new_n914));
  INV_X1    g713(.A(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n901), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n675), .A2(new_n896), .ZN(new_n917));
  AOI211_X1 g716(.A(new_n889), .B(new_n900), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n901), .ZN(new_n919));
  INV_X1    g718(.A(new_n903), .ZN(new_n920));
  INV_X1    g719(.A(new_n890), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n891), .B1(new_n844), .B2(KEYINPUT119), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n336), .B1(new_n922), .B2(new_n907), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n923), .B2(new_n909), .ZN(new_n924));
  INV_X1    g723(.A(new_n912), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n920), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n919), .B(new_n917), .C1(new_n926), .C2(new_n914), .ZN(new_n927));
  INV_X1    g726(.A(new_n900), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n888), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n918), .A2(new_n929), .ZN(G1344gat));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n916), .A2(new_n931), .A3(new_n385), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n919), .A2(new_n385), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n855), .A2(new_n264), .B1(new_n675), .B2(new_n386), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n902), .B1(new_n934), .B2(new_n512), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n893), .A2(new_n903), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(G148gat), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n931), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n893), .A2(new_n559), .A3(new_n385), .A4(new_n894), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(KEYINPUT59), .ZN(new_n942));
  AOI22_X1  g741(.A1(new_n938), .A2(new_n940), .B1(new_n939), .B2(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n932), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n385), .A2(new_n931), .ZN(new_n946));
  AOI211_X1 g745(.A(new_n901), .B(new_n946), .C1(new_n913), .C2(new_n915), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n942), .A2(new_n939), .ZN(new_n948));
  INV_X1    g747(.A(new_n940), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n937), .B2(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT123), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n945), .A2(new_n951), .ZN(G1345gat));
  AND3_X1   g751(.A1(new_n893), .A2(new_n559), .A3(new_n894), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n953), .A2(new_n490), .A3(new_n336), .ZN(new_n954));
  AND2_X1   g753(.A1(new_n916), .A2(new_n336), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n954), .B1(new_n955), .B2(new_n490), .ZN(G1346gat));
  AOI21_X1  g755(.A(G162gat), .B1(new_n953), .B2(new_n334), .ZN(new_n957));
  NOR2_X1   g756(.A1(new_n337), .A2(new_n491), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n957), .B1(new_n916), .B2(new_n958), .ZN(G1347gat));
  NOR2_X1   g758(.A1(new_n585), .A2(new_n559), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n706), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n893), .A2(new_n512), .A3(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n675), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n863), .A2(new_n868), .A3(new_n961), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n966), .A2(new_n411), .A3(new_n681), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT124), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n968), .B(new_n969), .ZN(G1348gat));
  OAI21_X1  g769(.A(G176gat), .B1(new_n964), .B2(new_n763), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n966), .A2(new_n412), .A3(new_n385), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1349gat));
  NAND2_X1  g772(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n974));
  XOR2_X1   g773(.A(new_n974), .B(KEYINPUT126), .Z(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n421), .B1(new_n963), .B2(new_n336), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n264), .A2(new_n418), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n966), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n977), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g779(.A1(KEYINPUT125), .A2(KEYINPUT60), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n976), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI221_X1 g781(.A(new_n975), .B1(KEYINPUT125), .B2(KEYINPUT60), .C1(new_n977), .C2(new_n979), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n982), .A2(new_n983), .ZN(G1350gat));
  NAND3_X1  g783(.A1(new_n966), .A2(new_n425), .A3(new_n334), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n963), .A2(new_n334), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(G190gat), .ZN(new_n988));
  AOI211_X1 g787(.A(KEYINPUT61), .B(new_n425), .C1(new_n963), .C2(new_n334), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n985), .B1(new_n988), .B2(new_n989), .ZN(G1351gat));
  NAND2_X1  g789(.A1(new_n935), .A2(new_n936), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n961), .A2(new_n708), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n991), .A2(new_n681), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT127), .ZN(new_n994));
  AOI21_X1  g793(.A(new_n656), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n995), .B1(new_n994), .B2(new_n993), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n863), .A2(new_n961), .ZN(new_n997));
  NOR2_X1   g796(.A1(new_n708), .A2(new_n512), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n999), .A2(new_n656), .A3(new_n681), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n996), .A2(new_n1000), .ZN(G1352gat));
  NOR2_X1   g800(.A1(new_n763), .A2(G204gat), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g802(.A(new_n1003), .B(KEYINPUT62), .Z(new_n1004));
  NAND2_X1  g803(.A1(new_n991), .A2(new_n992), .ZN(new_n1005));
  OAI21_X1  g804(.A(G204gat), .B1(new_n1005), .B2(new_n763), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1004), .A2(new_n1006), .ZN(G1353gat));
  INV_X1    g806(.A(G211gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n999), .A2(new_n1008), .A3(new_n336), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n991), .A2(new_n336), .A3(new_n992), .ZN(new_n1010));
  AND3_X1   g809(.A1(new_n1010), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1011));
  AOI21_X1  g810(.A(KEYINPUT63), .B1(new_n1010), .B2(G211gat), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(G1354gat));
  OAI21_X1  g812(.A(G218gat), .B1(new_n1005), .B2(new_n337), .ZN(new_n1014));
  INV_X1    g813(.A(G218gat), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n999), .A2(new_n1015), .A3(new_n334), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(G1355gat));
endmodule


