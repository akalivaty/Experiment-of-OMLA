//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 1 1 1 1 1 0 1 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983;
  NAND2_X1  g000(.A1(KEYINPUT2), .A2(G113), .ZN(new_n187));
  OAI21_X1  g001(.A(KEYINPUT66), .B1(KEYINPUT2), .B2(G113), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  NOR3_X1   g003(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G116), .ZN(new_n193));
  INV_X1    g007(.A(G116), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G119), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(new_n196), .ZN(new_n197));
  XNOR2_X1  g011(.A(G116), .B(G119), .ZN(new_n198));
  OAI211_X1 g012(.A(new_n198), .B(new_n187), .C1(new_n189), .C2(new_n190), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G143), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G146), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n202), .A2(new_n204), .A3(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(new_n203), .A3(G143), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n205), .B(G146), .C1(new_n201), .C2(KEYINPUT1), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G134), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G137), .ZN(new_n212));
  INV_X1    g026(.A(G137), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(G131), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT11), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n211), .B2(G137), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT65), .B1(new_n213), .B2(G134), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n211), .A3(G137), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(KEYINPUT11), .A3(G134), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n218), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n210), .B(new_n215), .C1(G131), .C2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT0), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(new_n201), .ZN(new_n226));
  NAND2_X1  g040(.A1(KEYINPUT0), .A2(G128), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n204), .A2(new_n206), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n204), .A2(new_n206), .A3(new_n227), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n217), .A2(new_n221), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n218), .A4(new_n220), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n222), .A2(G131), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n230), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n200), .B1(new_n224), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n237));
  XNOR2_X1  g051(.A(G143), .B(G146), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(new_n227), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n226), .A2(new_n227), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n239), .B1(new_n240), .B2(new_n238), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n222), .A2(G131), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n222), .A2(G131), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n241), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n200), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n245), .A3(new_n223), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n236), .A2(new_n237), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(new_n223), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT70), .A3(new_n200), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n247), .A2(KEYINPUT28), .A3(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n251), .B(G101), .ZN(new_n252));
  INV_X1    g066(.A(G953), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT67), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT67), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G953), .ZN(new_n256));
  AOI21_X1  g070(.A(G237), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G210), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n252), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n246), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n250), .A2(KEYINPUT29), .A3(new_n259), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G902), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT29), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n233), .A2(new_n234), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n230), .A2(KEYINPUT64), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT64), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n241), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n223), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n200), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n244), .A2(new_n245), .A3(KEYINPUT28), .A4(new_n223), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n261), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n259), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n264), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n244), .A2(KEYINPUT30), .A3(new_n223), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n234), .A2(new_n233), .B1(new_n230), .B2(KEYINPUT64), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n224), .B1(new_n277), .B2(new_n268), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n200), .B(new_n276), .C1(new_n278), .C2(KEYINPUT30), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n259), .B1(new_n279), .B2(new_n246), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n262), .B(new_n263), .C1(new_n275), .C2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT71), .ZN(new_n282));
  AND3_X1   g096(.A1(new_n281), .A2(new_n282), .A3(G472), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n282), .B1(new_n281), .B2(G472), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n273), .A2(new_n274), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n246), .A2(new_n259), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(KEYINPUT68), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n246), .A2(new_n289), .A3(new_n259), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT31), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n279), .A2(new_n288), .A3(KEYINPUT31), .A4(new_n290), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n286), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NOR2_X1   g109(.A1(G472), .A2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g111(.A(KEYINPUT69), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT32), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n293), .A2(new_n294), .ZN(new_n300));
  INV_X1    g114(.A(new_n286), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n299), .B1(new_n302), .B2(new_n296), .ZN(new_n303));
  NOR3_X1   g117(.A1(new_n295), .A2(KEYINPUT32), .A3(new_n297), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI211_X1 g119(.A(KEYINPUT69), .B(new_n299), .C1(new_n295), .C2(new_n297), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n285), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT72), .B1(new_n192), .B2(G128), .ZN(new_n308));
  OR2_X1    g122(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n309), .B(new_n310), .C1(G119), .C2(new_n201), .ZN(new_n311));
  XNOR2_X1  g125(.A(G119), .B(G128), .ZN(new_n312));
  XOR2_X1   g126(.A(KEYINPUT24), .B(G110), .Z(new_n313));
  OAI22_X1  g127(.A1(new_n311), .A2(G110), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  INV_X1    g130(.A(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G140), .ZN(new_n318));
  NAND4_X1  g132(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT73), .A4(KEYINPUT16), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n316), .A2(new_n318), .A3(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT73), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n316), .B2(KEYINPUT16), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n319), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G146), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n316), .A2(new_n318), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n314), .B(new_n324), .C1(G146), .C2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n203), .B(new_n319), .C1(new_n320), .C2(new_n322), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n324), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  OR3_X1    g143(.A1(new_n323), .A2(new_n327), .A3(G146), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n313), .A2(new_n312), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n311), .A2(G110), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n329), .A2(new_n330), .A3(new_n331), .A4(new_n332), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n326), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n254), .A2(new_n256), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n338), .B(KEYINPUT76), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n339), .A2(KEYINPUT22), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(KEYINPUT22), .ZN(new_n341));
  AND3_X1   g155(.A1(new_n340), .A2(G137), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(G137), .B1(new_n340), .B2(new_n341), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n336), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n333), .B(KEYINPUT75), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n342), .A2(new_n343), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n347), .A3(new_n326), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT25), .B1(new_n349), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(G217), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n351), .B1(G234), .B2(new_n263), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n348), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n354), .A3(new_n263), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n350), .A2(new_n352), .A3(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n349), .A2(KEYINPUT77), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n352), .A2(G902), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT77), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n357), .A2(new_n358), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n356), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(KEYINPUT78), .B1(new_n307), .B2(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n283), .A2(new_n284), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n302), .A2(new_n299), .A3(new_n296), .ZN(new_n365));
  OAI21_X1  g179(.A(KEYINPUT32), .B1(new_n295), .B2(new_n297), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n302), .A2(new_n296), .ZN(new_n367));
  AOI22_X1  g181(.A1(new_n365), .A2(new_n366), .B1(new_n367), .B2(KEYINPUT69), .ZN(new_n368));
  INV_X1    g182(.A(new_n306), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AND2_X1   g184(.A1(new_n356), .A2(new_n361), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT78), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(G475), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  INV_X1    g190(.A(G104), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n376), .B(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G237), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n337), .A2(G214), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n205), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT18), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n381), .B(new_n382), .C1(new_n383), .C2(new_n232), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n325), .B(G146), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n257), .A2(G143), .A3(G214), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n257), .B2(G214), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n384), .B(new_n385), .C1(new_n388), .C2(new_n383), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n329), .A2(new_n330), .ZN(new_n390));
  OAI211_X1 g204(.A(KEYINPUT17), .B(G131), .C1(new_n386), .C2(new_n387), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(KEYINPUT89), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n390), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT17), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n381), .A2(new_n232), .A3(new_n382), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT89), .B1(new_n396), .B2(new_n391), .ZN(new_n397));
  OAI211_X1 g211(.A(new_n378), .B(new_n389), .C1(new_n393), .C2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n388), .A2(new_n395), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n325), .A2(KEYINPUT19), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT19), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n401), .B1(new_n316), .B2(new_n318), .ZN(new_n402));
  NOR3_X1   g216(.A1(new_n400), .A2(G146), .A3(new_n402), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n403), .A2(KEYINPUT87), .ZN(new_n404));
  AOI22_X1  g218(.A1(new_n403), .A2(KEYINPUT87), .B1(G146), .B2(new_n323), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n399), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n389), .ZN(new_n407));
  INV_X1    g221(.A(new_n378), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n407), .A2(KEYINPUT88), .A3(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n398), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT88), .B1(new_n407), .B2(new_n408), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n375), .B(new_n263), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(KEYINPUT20), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT90), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n407), .A2(new_n408), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT88), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n419), .A2(new_n398), .A3(new_n409), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT20), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n420), .A2(new_n421), .A3(new_n375), .A4(new_n263), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n415), .A2(new_n416), .A3(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G952), .ZN(new_n424));
  AOI211_X1 g238(.A(G953), .B(new_n424), .C1(G234), .C2(G237), .ZN(new_n425));
  INV_X1    g239(.A(new_n337), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n263), .B1(G234), .B2(G237), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  XNOR2_X1  g242(.A(new_n428), .B(KEYINPUT94), .ZN(new_n429));
  XOR2_X1   g243(.A(KEYINPUT21), .B(G898), .Z(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n425), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g246(.A(G214), .B1(G237), .B2(G902), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G122), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n437));
  INV_X1    g251(.A(G107), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n437), .A2(G104), .A3(new_n438), .ZN(new_n439));
  AOI22_X1  g253(.A1(new_n377), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n440));
  OAI22_X1  g254(.A1(new_n377), .A2(G107), .B1(KEYINPUT79), .B2(KEYINPUT3), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G101), .ZN(new_n443));
  INV_X1    g257(.A(G101), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n439), .A2(new_n440), .A3(new_n441), .A4(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n443), .A2(KEYINPUT4), .A3(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT4), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n447), .A3(G101), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n446), .A2(new_n200), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT83), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT83), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT5), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n196), .A2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT83), .B(KEYINPUT5), .ZN(new_n456));
  OAI21_X1  g270(.A(G113), .B1(new_n456), .B2(new_n193), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n199), .B1(new_n455), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n438), .A2(G104), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n377), .A2(G107), .ZN(new_n460));
  OAI21_X1  g274(.A(G101), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n445), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT80), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n445), .A2(new_n464), .A3(new_n461), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n458), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n436), .B1(new_n449), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(G113), .ZN(new_n468));
  INV_X1    g282(.A(new_n193), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n468), .B1(new_n454), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n198), .A2(new_n456), .ZN(new_n471));
  OR3_X1    g285(.A1(KEYINPUT66), .A2(KEYINPUT2), .A3(G113), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n472), .A2(new_n188), .B1(KEYINPUT2), .B2(G113), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n470), .A2(new_n471), .B1(new_n473), .B2(new_n198), .ZN(new_n474));
  INV_X1    g288(.A(new_n465), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n464), .B1(new_n445), .B2(new_n461), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n446), .A2(new_n200), .A3(new_n448), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n435), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n467), .A2(KEYINPUT6), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n435), .B1(new_n477), .B2(new_n478), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT6), .ZN(new_n482));
  AOI21_X1  g296(.A(KEYINPUT84), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n467), .A2(KEYINPUT84), .A3(KEYINPUT6), .A4(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  OR3_X1    g300(.A1(new_n210), .A2(KEYINPUT85), .A3(G125), .ZN(new_n487));
  OAI21_X1  g301(.A(KEYINPUT85), .B1(new_n210), .B2(G125), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n487), .B(new_n488), .C1(new_n317), .C2(new_n241), .ZN(new_n489));
  INV_X1    g303(.A(G224), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n490), .A2(G953), .ZN(new_n491));
  XOR2_X1   g305(.A(new_n489), .B(new_n491), .Z(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n486), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT7), .B1(new_n490), .B2(G953), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n489), .B(new_n496), .ZN(new_n497));
  OR2_X1    g311(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n470), .A2(KEYINPUT86), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n498), .B(new_n499), .C1(new_n450), .C2(new_n196), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n462), .B1(new_n500), .B2(new_n199), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n435), .B(KEYINPUT8), .ZN(new_n502));
  AND2_X1   g316(.A1(new_n445), .A2(new_n461), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n502), .B1(new_n458), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n479), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n263), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n495), .A3(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(new_n495), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n492), .B1(new_n484), .B2(new_n485), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n509), .B1(new_n510), .B2(new_n506), .ZN(new_n511));
  AOI211_X1 g325(.A(new_n432), .B(new_n434), .C1(new_n508), .C2(new_n511), .ZN(new_n512));
  XNOR2_X1  g326(.A(G128), .B(G143), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(new_n211), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n194), .A2(KEYINPUT14), .A3(G122), .ZN(new_n515));
  XNOR2_X1  g329(.A(G116), .B(G122), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(G107), .B(new_n515), .C1(new_n517), .C2(KEYINPUT14), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n514), .B(new_n518), .C1(G107), .C2(new_n517), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n211), .B1(new_n513), .B2(KEYINPUT13), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n205), .A2(G128), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(KEYINPUT13), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT91), .Z(new_n523));
  XNOR2_X1  g337(.A(new_n516), .B(new_n438), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n513), .A2(new_n211), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n519), .B1(new_n523), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g341(.A(KEYINPUT9), .B(G234), .Z(new_n528));
  NAND3_X1  g342(.A1(new_n528), .A2(G217), .A3(new_n253), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT92), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n527), .A2(new_n529), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  OR3_X1    g347(.A1(new_n527), .A2(new_n531), .A3(new_n529), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n533), .A2(new_n534), .A3(new_n263), .ZN(new_n535));
  INV_X1    g349(.A(G478), .ZN(new_n536));
  NOR2_X1   g350(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT93), .A2(KEYINPUT15), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n536), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n535), .B(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n389), .B1(new_n393), .B2(new_n397), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n408), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n398), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n375), .B1(new_n545), .B2(new_n263), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n423), .A2(new_n512), .A3(new_n542), .A4(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n222), .B(new_n232), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n503), .A2(new_n210), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n462), .A2(new_n208), .A3(new_n209), .A4(new_n207), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n549), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT12), .B1(new_n265), .B2(KEYINPUT81), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  OAI211_X1 g368(.A(KEYINPUT10), .B(new_n210), .C1(new_n475), .C2(new_n476), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT10), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n446), .A2(new_n241), .A3(new_n448), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n555), .A2(new_n557), .A3(new_n549), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n337), .A2(G227), .ZN(new_n560));
  XNOR2_X1  g374(.A(G110), .B(G140), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n554), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n555), .A2(new_n557), .A3(new_n558), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(new_n265), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n562), .B1(new_n566), .B2(new_n559), .ZN(new_n567));
  OR2_X1    g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT82), .ZN(new_n569));
  INV_X1    g383(.A(G469), .ZN(new_n570));
  NAND4_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .A4(new_n263), .ZN(new_n571));
  OAI211_X1 g385(.A(new_n570), .B(new_n263), .C1(new_n564), .C2(new_n567), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT82), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(new_n559), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n554), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n576), .A2(new_n562), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n563), .B1(new_n265), .B2(new_n565), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g393(.A(G469), .B1(new_n579), .B2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n574), .A2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(G221), .ZN(new_n582));
  AOI21_X1  g396(.A(new_n582), .B1(new_n528), .B2(new_n263), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n548), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n374), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n587), .B(G101), .ZN(G3));
  OAI21_X1  g402(.A(G472), .B1(new_n295), .B2(G902), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n367), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n362), .A2(new_n585), .A3(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n432), .ZN(new_n592));
  AND3_X1   g406(.A1(new_n412), .A2(KEYINPUT90), .A3(KEYINPUT20), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT90), .B1(new_n412), .B2(KEYINPUT20), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n546), .B1(new_n595), .B2(new_n422), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n533), .A2(new_n534), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n530), .A2(KEYINPUT33), .A3(new_n532), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(G478), .A3(new_n263), .A4(new_n599), .ZN(new_n600));
  AND2_X1   g414(.A1(new_n536), .A2(KEYINPUT97), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n536), .A2(KEYINPUT97), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n535), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n600), .A2(new_n603), .ZN(new_n604));
  INV_X1    g418(.A(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n596), .A2(new_n605), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n510), .A2(new_n509), .A3(new_n506), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n434), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n508), .A2(KEYINPUT95), .A3(new_n511), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT96), .ZN(new_n611));
  AOI21_X1  g425(.A(KEYINPUT96), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n591), .A2(new_n592), .A3(new_n606), .A4(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(KEYINPUT98), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n614), .B(new_n616), .ZN(G6));
  XNOR2_X1  g431(.A(new_n422), .B(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n595), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n535), .B(new_n540), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n547), .A3(new_n620), .A4(new_n592), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT100), .ZN(new_n622));
  OR2_X1    g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n622), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n623), .A2(new_n591), .A3(new_n613), .A4(new_n624), .ZN(new_n625));
  XOR2_X1   g439(.A(KEYINPUT35), .B(G107), .Z(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G9));
  AOI21_X1  g441(.A(new_n354), .B1(new_n353), .B2(new_n263), .ZN(new_n628));
  AOI211_X1 g442(.A(KEYINPUT25), .B(G902), .C1(new_n345), .C2(new_n348), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n347), .A2(KEYINPUT36), .ZN(new_n631));
  OAI22_X1  g445(.A1(new_n345), .A2(KEYINPUT36), .B1(new_n631), .B2(new_n336), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n630), .A2(new_n352), .B1(new_n358), .B2(new_n632), .ZN(new_n633));
  NOR4_X1   g447(.A1(new_n548), .A2(new_n633), .A3(new_n585), .A4(new_n590), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(KEYINPUT37), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G110), .ZN(G12));
  INV_X1    g450(.A(new_n585), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n632), .A2(new_n358), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n356), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n613), .A2(new_n370), .A3(new_n637), .A4(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n546), .B1(new_n618), .B2(new_n595), .ZN(new_n641));
  INV_X1    g455(.A(G900), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n425), .B1(new_n429), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n641), .A2(new_n620), .A3(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n640), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(new_n201), .ZN(G30));
  XNOR2_X1  g461(.A(new_n643), .B(KEYINPUT39), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n585), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT40), .Z(new_n650));
  INV_X1    g464(.A(G472), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n247), .A2(new_n274), .A3(new_n249), .ZN(new_n652));
  AOI21_X1  g466(.A(G902), .B1(new_n291), .B2(new_n652), .ZN(new_n653));
  OAI22_X1  g467(.A1(new_n368), .A2(new_n369), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n596), .A2(new_n542), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n508), .A2(new_n511), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(KEYINPUT38), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n655), .A2(new_n657), .A3(new_n433), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n650), .A2(new_n633), .A3(new_n654), .A4(new_n658), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(G143), .ZN(G45));
  NAND2_X1  g474(.A1(new_n606), .A2(new_n644), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n640), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n203), .ZN(G48));
  NOR2_X1   g477(.A1(new_n307), .A2(new_n362), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n568), .A2(new_n263), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G469), .ZN(new_n666));
  AND3_X1   g480(.A1(new_n574), .A2(new_n584), .A3(new_n666), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n664), .A2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n606), .A2(new_n592), .A3(new_n613), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT41), .B(G113), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G15));
  NAND3_X1  g486(.A1(new_n623), .A2(new_n613), .A3(new_n624), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n668), .ZN(new_n674));
  XNOR2_X1  g488(.A(KEYINPUT101), .B(G116), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G18));
  INV_X1    g490(.A(KEYINPUT96), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n508), .A2(KEYINPUT95), .A3(new_n511), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n433), .B1(new_n508), .B2(KEYINPUT95), .ZN(new_n679));
  OAI21_X1  g493(.A(new_n677), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT96), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n667), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n680), .A2(new_n667), .A3(KEYINPUT102), .A4(new_n681), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n423), .A2(new_n547), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n687), .A2(new_n620), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n307), .A2(new_n432), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n686), .A2(new_n688), .A3(new_n639), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT103), .ZN(new_n691));
  INV_X1    g505(.A(new_n688), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n692), .B1(new_n684), .B2(new_n685), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT103), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n639), .A4(new_n689), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n691), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND2_X1  g511(.A1(new_n250), .A2(new_n261), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(new_n274), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n297), .B1(new_n300), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n589), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(KEYINPUT104), .B(G472), .C1(new_n295), .C2(G902), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n700), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n362), .ZN(new_n706));
  INV_X1    g520(.A(new_n682), .ZN(new_n707));
  AND4_X1   g521(.A1(new_n592), .A2(new_n706), .A3(new_n707), .A4(new_n655), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(G122), .Z(G24));
  NAND2_X1  g523(.A1(new_n639), .A2(new_n644), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n687), .A2(new_n604), .A3(new_n704), .ZN(new_n712));
  INV_X1    g526(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n686), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G125), .ZN(G27));
  INV_X1    g529(.A(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n580), .A2(KEYINPUT105), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT105), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n579), .A2(new_n718), .A3(new_n263), .ZN(new_n719));
  OAI21_X1  g533(.A(new_n717), .B1(new_n570), .B2(new_n719), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n583), .B1(new_n720), .B2(new_n574), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n656), .A2(new_n434), .ZN(new_n722));
  AND2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n664), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n716), .B1(new_n724), .B2(new_n661), .ZN(new_n725));
  INV_X1    g539(.A(new_n722), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n661), .A2(new_n726), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n303), .A2(new_n304), .A3(KEYINPUT106), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n285), .ZN(new_n729));
  OAI21_X1  g543(.A(KEYINPUT106), .B1(new_n303), .B2(new_n304), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n362), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n721), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G131), .ZN(G33));
  NOR2_X1   g548(.A1(new_n724), .A2(new_n645), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(new_n211), .ZN(G36));
  NOR2_X1   g550(.A1(new_n687), .A2(new_n605), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(KEYINPUT43), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n590), .A3(new_n639), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT44), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n722), .B1(new_n739), .B2(new_n740), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n579), .A2(KEYINPUT45), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n579), .A2(KEYINPUT45), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(G469), .A3(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(G469), .A2(G902), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT46), .ZN(new_n748));
  AOI22_X1  g562(.A1(new_n747), .A2(new_n748), .B1(new_n571), .B2(new_n573), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(new_n748), .B2(new_n747), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n584), .ZN(new_n751));
  NOR4_X1   g565(.A1(new_n741), .A2(new_n742), .A3(new_n648), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n213), .ZN(G39));
  XNOR2_X1  g567(.A(new_n751), .B(KEYINPUT47), .ZN(new_n754));
  INV_X1    g568(.A(new_n727), .ZN(new_n755));
  NOR4_X1   g569(.A1(new_n754), .A2(new_n371), .A3(new_n370), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(new_n315), .ZN(G42));
  AND2_X1   g571(.A1(new_n574), .A2(new_n666), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n758), .B(KEYINPUT49), .Z(new_n759));
  NOR4_X1   g573(.A1(new_n759), .A2(new_n657), .A3(new_n362), .A4(new_n605), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n654), .A2(new_n583), .A3(new_n687), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n760), .A2(new_n433), .A3(new_n761), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n708), .A2(new_n670), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n596), .A2(KEYINPUT107), .A3(new_n620), .A4(new_n512), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n423), .A2(new_n512), .A3(new_n547), .A4(new_n620), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT107), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n434), .B1(new_n508), .B2(new_n511), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n687), .A2(new_n604), .A3(new_n592), .A4(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n764), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(new_n591), .ZN(new_n771));
  INV_X1    g585(.A(new_n634), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n587), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n634), .B1(new_n374), .B2(new_n586), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n776), .A2(KEYINPUT108), .A3(new_n771), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n763), .B1(new_n775), .B2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n735), .B1(new_n725), .B2(new_n732), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n723), .A2(new_n713), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n641), .A2(new_n542), .ZN(new_n781));
  NOR4_X1   g595(.A1(new_n781), .A2(new_n307), .A3(new_n585), .A4(new_n726), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n711), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n674), .B1(new_n695), .B2(new_n691), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n778), .A2(new_n779), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n710), .B(new_n712), .C1(new_n684), .C2(new_n685), .ZN(new_n786));
  OAI21_X1  g600(.A(KEYINPUT109), .B1(new_n786), .B2(new_n646), .ZN(new_n787));
  OR2_X1    g601(.A1(new_n640), .A2(new_n645), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n714), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n596), .A2(new_n611), .A3(new_n612), .A4(new_n542), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n643), .B(KEYINPUT110), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n639), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n791), .A2(new_n654), .A3(new_n721), .A4(new_n793), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  INV_X1    g609(.A(new_n662), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n787), .A2(new_n790), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n796), .A2(new_n714), .A3(new_n788), .A4(new_n794), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n785), .A2(new_n801), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n708), .A2(new_n670), .ZN(new_n805));
  AND4_X1   g619(.A1(KEYINPUT108), .A2(new_n587), .A3(new_n771), .A4(new_n772), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT108), .B1(new_n776), .B2(new_n771), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n674), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n696), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n798), .B(new_n799), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n811), .A2(new_n779), .A3(new_n783), .A4(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT111), .B1(new_n813), .B2(new_n803), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n778), .A2(new_n783), .A3(new_n784), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n797), .A2(new_n800), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(KEYINPUT53), .A3(new_n779), .A4(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n804), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT112), .B1(new_n818), .B2(KEYINPUT54), .ZN(new_n819));
  XOR2_X1   g633(.A(KEYINPUT113), .B(KEYINPUT51), .Z(new_n820));
  AND2_X1   g634(.A1(new_n738), .A2(new_n425), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n821), .A2(new_n706), .ZN(new_n822));
  INV_X1    g636(.A(new_n667), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n822), .A2(new_n433), .A3(new_n657), .A4(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(KEYINPUT50), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n823), .A2(new_n726), .ZN(new_n826));
  INV_X1    g640(.A(new_n654), .ZN(new_n827));
  AND4_X1   g641(.A1(new_n371), .A2(new_n826), .A3(new_n827), .A4(new_n425), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n828), .A2(new_n596), .A3(new_n605), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n821), .A2(new_n826), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n639), .A2(new_n704), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n825), .B(new_n829), .C1(new_n830), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n758), .A2(new_n583), .ZN(new_n833));
  AOI211_X1 g647(.A(new_n726), .B(new_n822), .C1(new_n754), .C2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT114), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n820), .B1(new_n832), .B2(new_n835), .ZN(new_n836));
  XNOR2_X1  g650(.A(new_n798), .B(KEYINPUT52), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n803), .B1(new_n785), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n817), .A2(new_n802), .A3(new_n838), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n785), .A2(new_n801), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(KEYINPUT111), .A3(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT112), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT54), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  OR2_X1    g659(.A1(new_n813), .A2(new_n803), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n803), .B1(new_n785), .B2(new_n801), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n844), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n819), .A2(new_n836), .A3(new_n845), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT51), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n832), .A2(new_n851), .A3(new_n834), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n821), .A2(new_n731), .A3(new_n826), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT48), .B1(new_n853), .B2(KEYINPUT115), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(new_n686), .ZN(new_n857));
  OAI211_X1 g671(.A(G952), .B(new_n253), .C1(new_n822), .C2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(new_n858), .B1(new_n606), .B2(new_n828), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n854), .A2(new_n855), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n856), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT116), .ZN(new_n862));
  NOR3_X1   g676(.A1(new_n850), .A2(new_n852), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(G952), .A2(G953), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n762), .B1(new_n863), .B2(new_n864), .ZN(G75));
  INV_X1    g679(.A(KEYINPUT56), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n818), .A2(G902), .ZN(new_n867));
  INV_X1    g681(.A(G210), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n486), .B(new_n493), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT55), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n869), .A2(new_n871), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n337), .A2(G952), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n872), .A2(new_n873), .A3(new_n874), .ZN(G51));
  NAND2_X1  g689(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n842), .A2(new_n844), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n746), .A2(KEYINPUT57), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n746), .A2(KEYINPUT57), .ZN(new_n881));
  OAI21_X1  g695(.A(new_n568), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n867), .A2(new_n745), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n874), .B1(new_n882), .B2(new_n883), .ZN(G54));
  NAND4_X1  g698(.A1(new_n818), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n885));
  INV_X1    g699(.A(new_n420), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n874), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT117), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n839), .A2(KEYINPUT58), .A3(G902), .A4(new_n841), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n375), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n890), .B2(new_n420), .ZN(new_n891));
  NOR4_X1   g705(.A1(new_n889), .A2(KEYINPUT117), .A3(new_n375), .A4(new_n886), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT118), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n895), .B(new_n887), .C1(new_n891), .C2(new_n892), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n896), .ZN(G60));
  INV_X1    g711(.A(KEYINPUT119), .ZN(new_n898));
  AND2_X1   g712(.A1(new_n598), .A2(new_n599), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n819), .A2(new_n845), .A3(new_n849), .ZN(new_n900));
  NAND2_X1  g714(.A1(G478), .A2(G902), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT59), .Z(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n899), .B1(new_n900), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n899), .A2(new_n903), .ZN(new_n905));
  INV_X1    g719(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n878), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n874), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n898), .B1(new_n904), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n874), .B1(new_n878), .B2(new_n906), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n848), .B1(new_n877), .B2(KEYINPUT112), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n902), .B1(new_n912), .B2(new_n845), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(KEYINPUT119), .C1(new_n913), .C2(new_n899), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(G63));
  NAND2_X1  g729(.A1(new_n357), .A2(new_n360), .ZN(new_n916));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT60), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n916), .B1(new_n842), .B2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT61), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n918), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n818), .A2(new_n632), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n908), .A3(new_n924), .A4(new_n925), .ZN(new_n926));
  OR2_X1    g740(.A1(new_n924), .A2(KEYINPUT120), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n924), .A2(KEYINPUT120), .ZN(new_n928));
  AND4_X1   g742(.A1(new_n908), .A2(new_n927), .A3(new_n919), .A4(new_n928), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n926), .B1(new_n929), .B2(KEYINPUT61), .ZN(G66));
  AOI21_X1  g744(.A(new_n253), .B1(new_n430), .B2(G224), .ZN(new_n931));
  INV_X1    g745(.A(new_n811), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n337), .ZN(new_n933));
  OAI211_X1 g747(.A(new_n484), .B(new_n485), .C1(G898), .C2(new_n337), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT122), .Z(new_n935));
  XNOR2_X1  g749(.A(new_n933), .B(new_n935), .ZN(G69));
  MUX2_X1   g750(.A(new_n278), .B(new_n248), .S(KEYINPUT30), .Z(new_n937));
  NOR2_X1   g751(.A1(new_n400), .A2(new_n402), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n937), .B(new_n938), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n752), .A2(new_n756), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n649), .B1(new_n363), .B2(new_n373), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n687), .A2(new_n542), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n941), .B(new_n722), .C1(new_n606), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n787), .A2(new_n796), .A3(new_n790), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT123), .Z(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n659), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n946), .A2(KEYINPUT62), .A3(new_n659), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n944), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n939), .B1(new_n951), .B2(new_n426), .ZN(new_n952));
  INV_X1    g766(.A(new_n939), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n426), .A2(G900), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n751), .A2(new_n648), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n955), .A2(new_n731), .A3(new_n791), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT126), .Z(new_n957));
  NAND4_X1  g771(.A1(new_n940), .A2(new_n946), .A3(new_n779), .A4(new_n957), .ZN(new_n958));
  OAI211_X1 g772(.A(new_n953), .B(new_n954), .C1(new_n958), .C2(new_n426), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n952), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n337), .B1(G227), .B2(G900), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n952), .A2(KEYINPUT124), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n952), .A2(KEYINPUT124), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n959), .A3(new_n964), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n961), .B(KEYINPUT125), .Z(new_n966));
  OAI21_X1  g780(.A(new_n962), .B1(new_n965), .B2(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(new_n846), .A2(new_n847), .ZN(new_n968));
  NAND2_X1  g782(.A1(G472), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT63), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n279), .A2(new_n246), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n291), .B1(new_n972), .B2(new_n259), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n968), .A2(new_n970), .A3(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n951), .A2(new_n811), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n975), .A2(new_n970), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n976), .A2(new_n259), .A3(new_n971), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n970), .B1(new_n958), .B2(new_n932), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n978), .A2(new_n274), .A3(new_n972), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n908), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(KEYINPUT127), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n974), .B(new_n977), .C1(new_n981), .C2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(G57));
endmodule


