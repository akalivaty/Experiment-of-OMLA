//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:28 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n770, new_n771,
    new_n772, new_n773, new_n775, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n853, new_n854, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n967,
    new_n968;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(G22gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT2), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n207), .B1(new_n209), .B2(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT72), .B1(new_n209), .B2(new_n211), .ZN(new_n213));
  AND2_X1   g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n212), .A2(new_n213), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n210), .A2(G141gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n208), .A2(G148gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n207), .B(new_n221), .C1(new_n216), .C2(KEYINPUT72), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n218), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(G197gat), .B(G204gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT22), .ZN(new_n226));
  INV_X1    g025(.A(G211gat), .ZN(new_n227));
  INV_X1    g026(.A(G218gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n226), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G211gat), .B(G218gat), .ZN(new_n231));
  INV_X1    g030(.A(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n225), .A3(new_n229), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT29), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n224), .B1(new_n235), .B2(KEYINPUT3), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n218), .B2(new_n222), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n238), .B1(new_n239), .B2(KEYINPUT29), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n204), .B1(new_n236), .B2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n236), .A2(new_n240), .A3(new_n204), .ZN(new_n243));
  XOR2_X1   g042(.A(G78gat), .B(G106gat), .Z(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n243), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n244), .B1(new_n247), .B2(new_n241), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n203), .B1(new_n246), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(G228gat), .A2(G233gat), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n251), .B1(new_n240), .B2(KEYINPUT79), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n248), .A3(new_n203), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(new_n253), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n255), .B1(new_n256), .B2(new_n249), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n254), .A2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  AND3_X1   g058(.A1(new_n218), .A2(KEYINPUT3), .A3(new_n222), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n260), .A2(new_n239), .ZN(new_n261));
  INV_X1    g060(.A(G120gat), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G113gat), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(G120gat), .ZN(new_n265));
  AOI21_X1  g064(.A(KEYINPUT1), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AND2_X1   g065(.A1(G127gat), .A2(G134gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(G127gat), .A2(G134gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n269));
  NOR3_X1   g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OR2_X1    g069(.A1(G127gat), .A2(G134gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(G127gat), .A2(G134gat), .ZN(new_n272));
  AOI21_X1  g071(.A(KEYINPUT66), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n266), .B1(new_n270), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n271), .A2(new_n272), .ZN(new_n275));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(new_n266), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n271), .A2(KEYINPUT66), .A3(new_n272), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n269), .B1(new_n267), .B2(new_n268), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n266), .ZN(new_n282));
  AND3_X1   g081(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n278), .B1(new_n277), .B2(new_n282), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n261), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n261), .B(KEYINPUT74), .C1(new_n283), .C2(new_n284), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G113gat), .B(G120gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n271), .B(new_n272), .C1(new_n290), .C2(KEYINPUT1), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n291), .A2(KEYINPUT67), .B1(new_n281), .B2(new_n266), .ZN(new_n292));
  AND3_X1   g091(.A1(new_n281), .A2(KEYINPUT67), .A3(new_n266), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n223), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT76), .B1(new_n295), .B2(KEYINPUT4), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT75), .B(KEYINPUT4), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT76), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT4), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n294), .A2(new_n299), .A3(new_n300), .A4(new_n223), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n296), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(G225gat), .A2(G233gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n289), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT5), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n283), .A2(new_n284), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n295), .B1(new_n306), .B2(new_n223), .ZN(new_n307));
  INV_X1    g106(.A(new_n303), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n305), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n294), .A2(new_n223), .A3(new_n297), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n277), .A2(new_n282), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n300), .B1(new_n312), .B2(new_n224), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n308), .A2(KEYINPUT5), .ZN(new_n316));
  INV_X1    g115(.A(new_n288), .ZN(new_n317));
  OAI21_X1  g116(.A(KEYINPUT73), .B1(new_n292), .B2(new_n293), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n277), .A2(new_n278), .A3(new_n282), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT74), .B1(new_n320), .B2(new_n261), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n315), .B(new_n316), .C1(new_n317), .C2(new_n321), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT77), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n314), .B1(new_n287), .B2(new_n288), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n324), .B1(new_n325), .B2(new_n316), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n310), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G1gat), .B(G29gat), .ZN(new_n328));
  INV_X1    g127(.A(G85gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT0), .B(G57gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  XNOR2_X1  g132(.A(KEYINPUT78), .B(KEYINPUT6), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n327), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT83), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n327), .A2(KEYINPUT83), .A3(new_n333), .A4(new_n334), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n332), .B(new_n310), .C1(new_n323), .C2(new_n326), .ZN(new_n339));
  INV_X1    g138(.A(new_n334), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n322), .A2(KEYINPUT77), .ZN(new_n341));
  NAND4_X1  g140(.A1(new_n289), .A2(new_n324), .A3(new_n315), .A4(new_n316), .ZN(new_n342));
  AOI22_X1  g141(.A1(new_n341), .A2(new_n342), .B1(new_n304), .B2(new_n309), .ZN(new_n343));
  XNOR2_X1  g142(.A(new_n332), .B(KEYINPUT80), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI211_X1 g144(.A(new_n339), .B(new_n340), .C1(new_n343), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G169gat), .A2(G176gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(G183gat), .A2(G190gat), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n347), .B1(new_n348), .B2(KEYINPUT24), .ZN(new_n349));
  NOR2_X1   g148(.A1(G183gat), .A2(G190gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT24), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n352), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n349), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g153(.A1(G169gat), .A2(G176gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT23), .B1(new_n355), .B2(KEYINPUT64), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT64), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  OAI211_X1 g157(.A(new_n357), .B(new_n358), .C1(G169gat), .C2(G176gat), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n356), .A4(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT25), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n356), .A2(new_n359), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n352), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT24), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n363), .B(new_n347), .C1(new_n364), .C2(new_n350), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n361), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT28), .ZN(new_n368));
  XNOR2_X1  g167(.A(KEYINPUT27), .B(G183gat), .ZN(new_n369));
  INV_X1    g168(.A(G190gat), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT26), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n355), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n374), .A2(KEYINPUT65), .ZN(new_n375));
  INV_X1    g174(.A(new_n348), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n374), .A2(KEYINPUT65), .A3(new_n347), .A4(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n369), .A2(new_n368), .A3(new_n370), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n372), .A2(new_n377), .A3(new_n379), .A4(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G226gat), .ZN(new_n382));
  INV_X1    g181(.A(G233gat), .ZN(new_n383));
  NOR2_X1   g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND3_X1   g183(.A1(new_n367), .A2(new_n381), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n386), .B1(new_n382), .B2(new_n383), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n387), .B1(new_n367), .B2(new_n381), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n237), .B1(new_n385), .B2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n367), .A2(new_n381), .A3(new_n384), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n377), .A2(new_n379), .ZN(new_n391));
  INV_X1    g190(.A(new_n380), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n371), .ZN(new_n393));
  AOI22_X1  g192(.A1(new_n391), .A2(new_n393), .B1(new_n360), .B2(new_n366), .ZN(new_n394));
  OAI211_X1 g193(.A(new_n390), .B(new_n238), .C1(new_n394), .C2(new_n387), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n389), .A2(KEYINPUT69), .A3(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n385), .A2(new_n388), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT69), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n397), .A2(new_n398), .A3(new_n238), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT37), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G8gat), .B(G36gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(G64gat), .B(G92gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(new_n403), .B(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n395), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT38), .B1(new_n406), .B2(KEYINPUT37), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n405), .B1(new_n396), .B2(new_n399), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT38), .ZN(new_n412));
  INV_X1    g211(.A(new_n405), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n400), .B2(new_n401), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n396), .A2(KEYINPUT37), .A3(new_n399), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n337), .A2(new_n338), .A3(new_n346), .A4(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n341), .A2(new_n342), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n345), .B1(new_n419), .B2(new_n310), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n396), .A2(new_n399), .A3(new_n405), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT70), .ZN(new_n422));
  AOI22_X1  g221(.A1(KEYINPUT30), .A2(new_n409), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  AND4_X1   g222(.A1(new_n422), .A2(new_n400), .A3(KEYINPUT30), .A4(new_n413), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT30), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n420), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT81), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n325), .A2(KEYINPUT39), .A3(new_n303), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n429), .B1(new_n430), .B2(new_n344), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n315), .B1(new_n317), .B2(new_n321), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT39), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(new_n308), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(KEYINPUT81), .A3(new_n345), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n295), .B(new_n303), .C1(new_n306), .C2(new_n223), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n436), .B2(KEYINPUT82), .ZN(new_n437));
  OAI221_X1 g236(.A(new_n437), .B1(KEYINPUT82), .B2(new_n436), .C1(new_n303), .C2(new_n325), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n431), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n431), .A2(KEYINPUT40), .A3(new_n438), .A4(new_n435), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n428), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n259), .B1(new_n418), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT71), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n409), .A2(new_n422), .A3(KEYINPUT30), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n410), .A2(new_n426), .ZN(new_n447));
  AND2_X1   g246(.A1(new_n421), .A2(new_n422), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n445), .B(new_n446), .C1(new_n447), .C2(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(KEYINPUT71), .B1(new_n423), .B2(new_n424), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n449), .A2(new_n450), .A3(new_n427), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n339), .A2(new_n340), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n343), .A2(new_n332), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n335), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n451), .A2(new_n454), .A3(new_n259), .ZN(new_n455));
  INV_X1    g254(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n394), .A2(new_n312), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n367), .A2(new_n381), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(new_n294), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n457), .A2(new_n459), .A3(G227gat), .A4(G233gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT32), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(KEYINPUT34), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT33), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n457), .A2(new_n459), .ZN(new_n465));
  NAND2_X1  g264(.A1(G227gat), .A2(G233gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(G71gat), .B(G99gat), .ZN(new_n469));
  XOR2_X1   g268(.A(new_n468), .B(new_n469), .Z(new_n470));
  NAND3_X1  g269(.A1(new_n464), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT34), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n460), .A2(KEYINPUT32), .A3(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n470), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n465), .B(new_n466), .C1(new_n463), .C2(new_n474), .ZN(new_n475));
  AND4_X1   g274(.A1(new_n462), .A2(new_n471), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  AOI22_X1  g275(.A1(new_n471), .A2(new_n475), .B1(new_n462), .B2(new_n473), .ZN(new_n477));
  AND2_X1   g276(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n478));
  NOR2_X1   g277(.A1(KEYINPUT68), .A2(KEYINPUT36), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NOR3_X1   g279(.A1(new_n476), .A2(new_n477), .A3(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n476), .A2(new_n477), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n482), .A2(new_n478), .ZN(new_n483));
  OAI22_X1  g282(.A1(new_n444), .A2(new_n456), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n334), .B1(new_n343), .B2(new_n332), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n327), .A2(new_n344), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n336), .A2(new_n335), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n487), .A2(new_n338), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n258), .A2(new_n482), .A3(new_n427), .A4(new_n425), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT35), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n258), .A2(new_n482), .A3(KEYINPUT84), .ZN(new_n493));
  AOI21_X1  g292(.A(KEYINPUT84), .B1(new_n258), .B2(new_n482), .ZN(new_n494));
  NOR3_X1   g293(.A1(new_n493), .A2(new_n494), .A3(new_n492), .ZN(new_n495));
  AND2_X1   g294(.A1(new_n451), .A2(new_n454), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n491), .A2(new_n492), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n484), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NOR3_X1   g299(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n501));
  INV_X1    g300(.A(G29gat), .ZN(new_n502));
  INV_X1    g301(.A(G36gat), .ZN(new_n503));
  OAI22_X1  g302(.A1(new_n500), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G43gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(G50gat), .ZN(new_n506));
  INV_X1    g305(.A(G50gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(G43gat), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT15), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n509), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT85), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n508), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT86), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n506), .B(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT15), .ZN(new_n517));
  AOI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n510), .B1(new_n518), .B2(new_n504), .ZN(new_n519));
  OAI21_X1  g318(.A(KEYINPUT87), .B1(new_n519), .B2(KEYINPUT17), .ZN(new_n520));
  XNOR2_X1  g319(.A(G15gat), .B(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT16), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n521), .B1(new_n522), .B2(G1gat), .ZN(new_n523));
  OAI21_X1  g322(.A(new_n523), .B1(G1gat), .B2(new_n521), .ZN(new_n524));
  INV_X1    g323(.A(G8gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n520), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT17), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT87), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n528), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n530), .A2(new_n519), .ZN(new_n531));
  OR2_X1    g330(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(G229gat), .A2(G233gat), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n533), .B(KEYINPUT88), .Z(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(KEYINPUT18), .A3(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n527), .B2(new_n531), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT18), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n519), .B(new_n526), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT89), .B(KEYINPUT13), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n534), .B(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n535), .A2(new_n538), .A3(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G113gat), .B(G141gat), .ZN(new_n544));
  INV_X1    g343(.A(G197gat), .ZN(new_n545));
  XNOR2_X1  g344(.A(new_n544), .B(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT11), .B(G169gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT12), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n543), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n535), .A2(new_n538), .A3(new_n542), .A4(new_n549), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT9), .ZN(new_n555));
  XOR2_X1   g354(.A(G57gat), .B(G64gat), .Z(new_n556));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n557), .B2(new_n556), .ZN(new_n559));
  XOR2_X1   g358(.A(G71gat), .B(G78gat), .Z(new_n560));
  NAND2_X1  g359(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n564), .B1(new_n562), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n565), .A2(new_n556), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(KEYINPUT91), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT91), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n556), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT92), .B(KEYINPUT21), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  XOR2_X1   g372(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n574));
  XNOR2_X1  g373(.A(new_n573), .B(new_n574), .ZN(new_n575));
  AOI22_X1  g374(.A1(new_n559), .A2(new_n560), .B1(new_n569), .B2(new_n567), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(KEYINPUT21), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n526), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n579));
  INV_X1    g378(.A(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n575), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n574), .ZN(new_n583));
  XNOR2_X1  g382(.A(new_n573), .B(new_n583), .ZN(new_n584));
  OR2_X1    g383(.A1(new_n578), .A2(KEYINPUT95), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n584), .A2(new_n585), .A3(new_n579), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(G127gat), .B(G155gat), .Z(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(new_n588), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n582), .A2(new_n586), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(G183gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(G211gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT93), .B(KEYINPUT94), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n592), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n589), .A2(new_n591), .A3(new_n597), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G92gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n329), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT7), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n605), .B1(new_n329), .B2(new_n603), .ZN(new_n606));
  NAND3_X1  g405(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n604), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(G99gat), .B(G106gat), .Z(new_n609));
  OAI21_X1  g408(.A(KEYINPUT99), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n561), .A2(new_n610), .A3(new_n570), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n608), .B(new_n609), .ZN(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G230gat), .A2(G233gat), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n576), .A2(new_n612), .A3(new_n610), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G120gat), .B(G148gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G176gat), .B(G204gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT10), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n571), .A2(new_n623), .A3(new_n612), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n576), .A2(new_n612), .A3(new_n610), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n612), .B1(new_n576), .B2(new_n610), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n617), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n630), .A2(KEYINPUT100), .A3(new_n623), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n624), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n615), .B1(new_n632), .B2(KEYINPUT101), .ZN(new_n633));
  INV_X1    g432(.A(new_n624), .ZN(new_n634));
  AOI21_X1  g433(.A(KEYINPUT100), .B1(new_n630), .B2(new_n623), .ZN(new_n635));
  AOI211_X1 g434(.A(new_n628), .B(KEYINPUT10), .C1(new_n614), .C2(new_n617), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT101), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  OAI211_X1 g438(.A(new_n618), .B(new_n622), .C1(new_n633), .C2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n637), .A2(new_n615), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n641), .A2(new_n618), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n621), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(G190gat), .B(G218gat), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT41), .ZN(new_n647));
  NAND2_X1  g446(.A1(G232gat), .A2(G233gat), .ZN(new_n648));
  OAI22_X1  g447(.A1(new_n519), .A2(new_n612), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT97), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT97), .ZN(new_n651));
  OAI221_X1 g450(.A(new_n651), .B1(new_n647), .B2(new_n648), .C1(new_n519), .C2(new_n612), .ZN(new_n652));
  AND2_X1   g451(.A1(new_n650), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n519), .ZN(new_n654));
  AOI21_X1  g453(.A(new_n613), .B1(new_n654), .B2(new_n528), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n519), .A2(KEYINPUT17), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n646), .B1(new_n653), .B2(new_n657), .ZN(new_n658));
  AOI22_X1  g457(.A1(new_n650), .A2(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n645), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n648), .A2(new_n647), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT96), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  AND4_X1   g463(.A1(KEYINPUT98), .A2(new_n658), .A3(new_n660), .A4(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT98), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n659), .B2(new_n645), .ZN(new_n667));
  AOI22_X1  g466(.A1(new_n667), .A2(new_n664), .B1(new_n658), .B2(new_n660), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NOR4_X1   g468(.A1(new_n554), .A2(new_n601), .A3(new_n644), .A4(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n498), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n454), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(G1gat), .ZN(G1324gat));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n425), .A2(new_n427), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n671), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n671), .ZN(new_n680));
  INV_X1    g479(.A(new_n676), .ZN(new_n681));
  OAI21_X1  g480(.A(G8gat), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n675), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(KEYINPUT42), .B1(new_n677), .B2(new_n678), .ZN(new_n684));
  OR3_X1    g483(.A1(new_n683), .A2(KEYINPUT102), .A3(new_n684), .ZN(new_n685));
  OAI21_X1  g484(.A(KEYINPUT102), .B1(new_n683), .B2(new_n684), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(G1325gat));
  AOI21_X1  g486(.A(G15gat), .B1(new_n671), .B2(new_n482), .ZN(new_n688));
  INV_X1    g487(.A(new_n481), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT103), .ZN(new_n690));
  OAI211_X1 g489(.A(new_n689), .B(new_n690), .C1(new_n482), .C2(new_n478), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT103), .B1(new_n483), .B2(new_n481), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT104), .Z(new_n695));
  AOI21_X1  g494(.A(new_n688), .B1(new_n671), .B2(new_n695), .ZN(G1326gat));
  NAND2_X1  g495(.A1(new_n671), .A2(new_n259), .ZN(new_n697));
  XNOR2_X1  g496(.A(KEYINPUT43), .B(G22gat), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n697), .B(new_n698), .ZN(G1327gat));
  INV_X1    g498(.A(new_n669), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n484), .B2(new_n497), .ZN(new_n701));
  INV_X1    g500(.A(new_n601), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n702), .A2(new_n554), .A3(new_n644), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n704), .A2(new_n502), .A3(new_n672), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n418), .A2(new_n443), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n258), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n693), .B1(new_n710), .B2(new_n455), .ZN(new_n711));
  INV_X1    g510(.A(new_n494), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n258), .A2(new_n482), .A3(KEYINPUT84), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n712), .A2(KEYINPUT35), .A3(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n451), .A2(new_n454), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n489), .B1(new_n487), .B2(new_n338), .ZN(new_n716));
  OAI22_X1  g515(.A1(new_n714), .A2(new_n715), .B1(new_n716), .B2(KEYINPUT35), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT106), .B1(new_n711), .B2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n693), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n719), .B1(new_n444), .B2(new_n456), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT106), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n497), .A2(new_n720), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n708), .B1(new_n718), .B2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT44), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n701), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n723), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n703), .B(KEYINPUT105), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n728), .A2(KEYINPUT107), .A3(new_n672), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G29gat), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT107), .B1(new_n728), .B2(new_n672), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n706), .B1(new_n730), .B2(new_n731), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n704), .A2(new_n503), .A3(new_n676), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(KEYINPUT46), .Z(new_n734));
  NOR3_X1   g533(.A1(new_n726), .A2(new_n681), .A3(new_n727), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n503), .B2(new_n735), .ZN(G1329gat));
  NAND4_X1  g535(.A1(new_n701), .A2(new_n505), .A3(new_n482), .A4(new_n703), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT109), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g539(.A(new_n727), .ZN(new_n741));
  OAI211_X1 g540(.A(new_n693), .B(new_n741), .C1(new_n723), .C2(new_n725), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(KEYINPUT110), .ZN(new_n743));
  OAI21_X1  g542(.A(G43gat), .B1(new_n742), .B2(KEYINPUT110), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT108), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n742), .A2(new_n746), .A3(G43gat), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n742), .B2(G43gat), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(new_n748), .A3(new_n738), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND3_X1  g549(.A1(new_n704), .A2(new_n507), .A3(new_n259), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n726), .A2(new_n258), .A3(new_n727), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n751), .B1(new_n752), .B2(new_n507), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT48), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OAI211_X1 g554(.A(KEYINPUT48), .B(new_n751), .C1(new_n752), .C2(new_n507), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(G1331gat));
  NAND2_X1  g556(.A1(new_n718), .A2(new_n722), .ZN(new_n758));
  INV_X1    g557(.A(new_n644), .ZN(new_n759));
  NOR4_X1   g558(.A1(new_n759), .A2(new_n601), .A3(new_n553), .A4(new_n669), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(new_n761));
  NOR2_X1   g560(.A1(new_n761), .A2(new_n454), .ZN(new_n762));
  XNOR2_X1  g561(.A(KEYINPUT111), .B(G57gat), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(G1332gat));
  NOR2_X1   g563(.A1(new_n761), .A2(new_n681), .ZN(new_n765));
  NOR2_X1   g564(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n766));
  AND2_X1   g565(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n768), .B1(new_n765), .B2(new_n766), .ZN(G1333gat));
  OAI21_X1  g568(.A(G71gat), .B1(new_n761), .B2(new_n719), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n482), .A2(new_n562), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n770), .B1(new_n761), .B2(new_n771), .ZN(new_n772));
  XNOR2_X1  g571(.A(KEYINPUT112), .B(KEYINPUT50), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1334gat));
  NOR2_X1   g573(.A1(new_n761), .A2(new_n258), .ZN(new_n775));
  XOR2_X1   g574(.A(KEYINPUT113), .B(G78gat), .Z(new_n776));
  XNOR2_X1  g575(.A(new_n775), .B(new_n776), .ZN(G1335gat));
  NAND2_X1  g576(.A1(new_n497), .A2(new_n720), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n702), .A2(new_n553), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT114), .ZN(new_n780));
  INV_X1    g579(.A(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n778), .A2(new_n669), .A3(new_n781), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(KEYINPUT51), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n783), .A2(new_n759), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g584(.A(G85gat), .B1(new_n785), .B2(new_n672), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n726), .A2(new_n759), .A3(new_n780), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n672), .A2(G85gat), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(G1336gat));
  NOR2_X1   g589(.A1(new_n681), .A2(G92gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n785), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n780), .A2(new_n759), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n676), .B(new_n794), .C1(new_n723), .C2(new_n725), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT115), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g600(.A(KEYINPUT51), .B1(new_n782), .B2(new_n798), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n759), .A3(new_n802), .ZN(new_n803));
  AOI22_X1  g602(.A1(new_n803), .A2(new_n791), .B1(G92gat), .B2(new_n795), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n797), .B1(new_n804), .B2(new_n793), .ZN(G1337gat));
  AOI21_X1  g604(.A(G99gat), .B1(new_n785), .B2(new_n482), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n693), .A2(G99gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n787), .B2(new_n807), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n258), .A2(G106gat), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT53), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n259), .B(new_n794), .C1(new_n723), .C2(new_n725), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G106gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n810), .A2(new_n811), .A3(new_n813), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n803), .A2(new_n809), .B1(G106gat), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n815), .B2(new_n811), .ZN(G1339gat));
  NOR4_X1   g615(.A1(new_n601), .A2(new_n644), .A3(new_n553), .A4(new_n669), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT55), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n616), .B(new_n634), .C1(new_n635), .C2(new_n636), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT54), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n616), .B1(new_n637), .B2(new_n638), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n632), .A2(KEYINPUT101), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n621), .B1(new_n641), .B2(KEYINPUT54), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n818), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT54), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n632), .B2(new_n616), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n633), .B2(new_n639), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n632), .A2(new_n616), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n622), .B1(new_n829), .B2(new_n826), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n828), .A2(KEYINPUT55), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n532), .A2(new_n534), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n539), .A2(new_n541), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n548), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  AND2_X1   g633(.A1(new_n552), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n825), .A2(new_n831), .A3(new_n640), .A4(new_n835), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n702), .B1(new_n836), .B2(new_n669), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n669), .B1(new_n644), .B2(new_n835), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n825), .A2(new_n831), .A3(new_n640), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n838), .B1(new_n839), .B2(new_n554), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n817), .B1(new_n837), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n672), .A2(new_n681), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n493), .A2(new_n494), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n264), .A3(new_n553), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n258), .A2(new_n482), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n841), .A2(new_n848), .A3(new_n842), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  OAI21_X1  g649(.A(G113gat), .B1(new_n850), .B2(new_n554), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n847), .A2(new_n851), .ZN(G1340gat));
  NAND3_X1  g651(.A1(new_n846), .A2(new_n262), .A3(new_n644), .ZN(new_n853));
  OAI21_X1  g652(.A(G120gat), .B1(new_n850), .B2(new_n759), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(G1341gat));
  NAND3_X1  g654(.A1(new_n849), .A2(G127gat), .A3(new_n702), .ZN(new_n856));
  OAI21_X1  g655(.A(KEYINPUT116), .B1(new_n845), .B2(new_n601), .ZN(new_n857));
  INV_X1    g656(.A(G127gat), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n845), .A2(KEYINPUT116), .A3(new_n601), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n861), .B(KEYINPUT117), .ZN(G1342gat));
  NOR3_X1   g661(.A1(new_n845), .A2(G134gat), .A3(new_n700), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT56), .ZN(new_n864));
  OAI21_X1  g663(.A(G134gat), .B1(new_n850), .B2(new_n700), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  NAND2_X1  g668(.A1(new_n837), .A2(new_n840), .ZN(new_n870));
  INV_X1    g669(.A(new_n817), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n872), .A2(KEYINPUT57), .A3(new_n259), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT57), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n841), .B2(new_n258), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n693), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n842), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(G141gat), .B1(new_n878), .B2(new_n554), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n693), .A2(new_n258), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n843), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n553), .A2(new_n208), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g683(.A(new_n881), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n210), .A3(new_n644), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n873), .A2(new_n875), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n887), .A2(new_n644), .A3(new_n719), .A4(new_n877), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  AND3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(G148gat), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n889), .B1(new_n888), .B2(G148gat), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n886), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT119), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g693(.A(KEYINPUT119), .B(new_n886), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(G1345gat));
  AOI21_X1  g695(.A(G155gat), .B1(new_n885), .B2(new_n702), .ZN(new_n897));
  INV_X1    g696(.A(new_n878), .ZN(new_n898));
  NOR2_X1   g697(.A1(new_n601), .A2(new_n205), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n897), .B1(new_n898), .B2(new_n899), .ZN(G1346gat));
  NAND3_X1  g699(.A1(new_n885), .A2(new_n206), .A3(new_n669), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT120), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n669), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(G162gat), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n902), .B1(new_n898), .B2(new_n669), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n672), .A2(new_n681), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n872), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n908), .A2(new_n494), .A3(new_n493), .ZN(new_n909));
  INV_X1    g708(.A(G169gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n909), .A2(new_n910), .A3(new_n553), .ZN(new_n911));
  NOR3_X1   g710(.A1(new_n841), .A2(new_n672), .A3(new_n681), .ZN(new_n912));
  INV_X1    g711(.A(new_n848), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n554), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n911), .A2(new_n915), .ZN(G1348gat));
  AOI21_X1  g715(.A(G176gat), .B1(new_n909), .B2(new_n644), .ZN(new_n917));
  INV_X1    g716(.A(G176gat), .ZN(new_n918));
  NOR3_X1   g717(.A1(new_n914), .A2(new_n918), .A3(new_n759), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n917), .A2(new_n919), .ZN(G1349gat));
  OAI21_X1  g719(.A(G183gat), .B1(new_n914), .B2(new_n601), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n702), .A2(new_n369), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n912), .A2(new_n844), .A3(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT121), .ZN(new_n924));
  AND2_X1   g723(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n923), .A2(new_n924), .ZN(new_n926));
  OAI211_X1 g725(.A(KEYINPUT123), .B(new_n921), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT60), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT60), .ZN(new_n932));
  OAI211_X1 g731(.A(KEYINPUT122), .B(new_n921), .C1(new_n925), .C2(new_n926), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n931), .A2(new_n932), .A3(new_n933), .ZN(G1350gat));
  NAND3_X1  g733(.A1(new_n909), .A2(new_n370), .A3(new_n669), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT124), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n908), .A2(new_n848), .A3(new_n700), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n936), .B(KEYINPUT61), .C1(new_n937), .C2(new_n370), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  OAI211_X1 g738(.A(new_n939), .B(G190gat), .C1(new_n914), .C2(new_n700), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g740(.A(G190gat), .B1(new_n914), .B2(new_n700), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n936), .B1(new_n942), .B2(KEYINPUT61), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(KEYINPUT125), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT125), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n946), .B(new_n935), .C1(new_n941), .C2(new_n943), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1351gat));
  NAND2_X1  g747(.A1(new_n876), .A2(new_n907), .ZN(new_n949));
  OAI21_X1  g748(.A(G197gat), .B1(new_n949), .B2(new_n554), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n908), .A2(new_n258), .A3(new_n693), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT126), .Z(new_n952));
  NAND2_X1  g751(.A1(new_n553), .A2(new_n545), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1352gat));
  XNOR2_X1  g753(.A(KEYINPUT127), .B(G204gat), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n759), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n951), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g756(.A(new_n957), .B(KEYINPUT62), .Z(new_n958));
  OAI21_X1  g757(.A(new_n955), .B1(new_n949), .B2(new_n759), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1353gat));
  OAI21_X1  g759(.A(G211gat), .B1(new_n949), .B2(new_n601), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT63), .ZN(new_n962));
  AND2_X1   g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(new_n962), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n702), .A2(new_n227), .ZN(new_n965));
  OAI22_X1  g764(.A1(new_n963), .A2(new_n964), .B1(new_n952), .B2(new_n965), .ZN(G1354gat));
  NOR3_X1   g765(.A1(new_n949), .A2(new_n228), .A3(new_n700), .ZN(new_n967));
  OR2_X1    g766(.A1(new_n952), .A2(new_n700), .ZN(new_n968));
  AOI21_X1  g767(.A(new_n967), .B1(new_n968), .B2(new_n228), .ZN(G1355gat));
endmodule


