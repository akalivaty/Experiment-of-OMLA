//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  XOR2_X1   g000(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n187));
  NOR2_X1   g001(.A1(G237), .A2(G953), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G210), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT26), .B(G101), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT65), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(KEYINPUT11), .A2(G134), .ZN(new_n196));
  NAND2_X1  g010(.A1(KEYINPUT65), .A2(G137), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n195), .A2(new_n196), .A3(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT11), .A2(G134), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT11), .A2(G134), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n199), .B1(new_n200), .B2(G137), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n198), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n197), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT65), .A2(G137), .ZN(new_n206));
  NOR3_X1   g020(.A1(new_n205), .A2(new_n206), .A3(G134), .ZN(new_n207));
  INV_X1    g021(.A(G134), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(new_n194), .ZN(new_n209));
  OAI21_X1  g023(.A(G131), .B1(new_n207), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n204), .A2(new_n210), .A3(KEYINPUT70), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n195), .A2(new_n208), .A3(new_n197), .ZN(new_n213));
  INV_X1    g027(.A(new_n209), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n203), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(G131), .B1(new_n198), .B2(new_n201), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G146), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G143), .ZN(new_n219));
  INV_X1    g033(.A(G143), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G146), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT1), .B1(new_n220), .B2(G146), .ZN(new_n223));
  OAI21_X1  g037(.A(G128), .B1(new_n223), .B2(KEYINPUT67), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT67), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n225), .B1(new_n219), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n222), .B1(new_n224), .B2(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(G143), .B(G146), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT1), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n228), .A2(new_n229), .A3(G128), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n211), .A2(new_n217), .A3(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G119), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT68), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G119), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n236), .A3(G116), .ZN(new_n237));
  INV_X1    g051(.A(G116), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n238), .A2(G119), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT2), .B(G113), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(new_n241), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(new_n237), .A3(new_n239), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n242), .A2(new_n244), .A3(KEYINPUT69), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT69), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n240), .A2(new_n246), .A3(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT0), .ZN(new_n249));
  INV_X1    g063(.A(G128), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n228), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n249), .A2(new_n250), .A3(KEYINPUT64), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT64), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n253), .B1(KEYINPUT0), .B2(G128), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n252), .A2(new_n254), .B1(KEYINPUT0), .B2(G128), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n251), .B1(new_n255), .B2(new_n228), .ZN(new_n256));
  OR2_X1    g070(.A1(new_n203), .A2(KEYINPUT66), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n257), .B1(new_n198), .B2(new_n201), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n198), .A2(new_n257), .A3(new_n201), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n256), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n232), .A2(new_n248), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(KEYINPUT28), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT28), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n232), .A2(new_n263), .A3(new_n248), .A4(new_n260), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n248), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n229), .B1(G143), .B2(new_n218), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n250), .B1(new_n267), .B2(new_n225), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n223), .A2(KEYINPUT67), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n228), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND4_X1   g084(.A1(new_n229), .A2(new_n219), .A3(new_n221), .A4(G128), .ZN(new_n271));
  OAI22_X1  g085(.A1(new_n270), .A2(new_n271), .B1(new_n215), .B2(new_n216), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n260), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n266), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n192), .B1(new_n265), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT30), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n276), .B1(new_n232), .B2(new_n260), .ZN(new_n277));
  AND3_X1   g091(.A1(new_n272), .A2(new_n276), .A3(new_n260), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n266), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n261), .A2(new_n192), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT31), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT31), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n275), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NOR2_X1   g099(.A1(G472), .A2(G902), .ZN(new_n286));
  INV_X1    g100(.A(new_n286), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n285), .A2(KEYINPUT32), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  AND3_X1   g103(.A1(new_n279), .A2(new_n280), .A3(KEYINPUT31), .ZN(new_n290));
  AOI21_X1  g104(.A(KEYINPUT31), .B1(new_n279), .B2(new_n280), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n262), .A2(new_n264), .B1(new_n266), .B2(new_n273), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n290), .A2(new_n291), .B1(new_n192), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n289), .B1(new_n293), .B2(new_n286), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n288), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G472), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n279), .A2(new_n261), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT72), .B1(new_n298), .B2(new_n192), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT72), .ZN(new_n300));
  INV_X1    g114(.A(new_n192), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT29), .B1(new_n292), .B2(new_n192), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n299), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n248), .B1(new_n232), .B2(new_n260), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(new_n262), .B2(new_n264), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n192), .A2(KEYINPUT29), .ZN(new_n307));
  AOI21_X1  g121(.A(G902), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n296), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g123(.A(KEYINPUT73), .B1(new_n295), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n308), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT32), .B1(new_n285), .B2(new_n287), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n293), .A2(new_n289), .A3(new_n286), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n312), .A2(new_n313), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n310), .A2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT74), .B(G217), .ZN(new_n319));
  INV_X1    g133(.A(G902), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(G234), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G140), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n322), .A2(new_n323), .A3(G125), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n325), .A2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(G146), .B(new_n324), .C1(new_n328), .C2(new_n322), .ZN(new_n329));
  XNOR2_X1  g143(.A(G125), .B(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(new_n218), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n234), .A2(new_n236), .A3(G128), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  OAI21_X1  g148(.A(KEYINPUT75), .B1(new_n233), .B2(G128), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT68), .B(G119), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n335), .B1(new_n336), .B2(G128), .ZN(new_n337));
  XOR2_X1   g151(.A(KEYINPUT24), .B(G110), .Z(new_n338));
  NOR3_X1   g152(.A1(new_n334), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n234), .A2(new_n236), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT23), .B1(new_n340), .B2(new_n250), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n250), .A2(KEYINPUT23), .A3(G119), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n333), .A2(new_n342), .ZN(new_n343));
  NOR3_X1   g157(.A1(new_n341), .A2(new_n343), .A3(G110), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n332), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n324), .B1(new_n328), .B2(new_n322), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n218), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n329), .ZN(new_n348));
  OAI21_X1  g162(.A(G110), .B1(new_n341), .B2(new_n343), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n338), .B1(new_n334), .B2(new_n337), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT76), .B1(new_n345), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n345), .A2(KEYINPUT76), .A3(new_n351), .ZN(new_n354));
  XOR2_X1   g168(.A(KEYINPUT22), .B(G137), .Z(new_n355));
  INV_X1    g169(.A(G953), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n356), .A2(G221), .A3(G234), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n355), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n353), .A2(new_n354), .A3(new_n359), .ZN(new_n360));
  AOI211_X1 g174(.A(KEYINPUT76), .B(new_n359), .C1(new_n345), .C2(new_n351), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(KEYINPUT25), .B1(new_n363), .B2(new_n320), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  AOI211_X1 g179(.A(new_n365), .B(G902), .C1(new_n360), .C2(new_n362), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n321), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n321), .A2(G902), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n363), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT81), .B(G469), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n219), .A2(new_n225), .A3(KEYINPUT1), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n269), .A2(G128), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n271), .B1(new_n374), .B2(new_n222), .ZN(new_n375));
  XNOR2_X1  g189(.A(G104), .B(G107), .ZN(new_n376));
  INV_X1    g190(.A(G101), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT77), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G104), .ZN(new_n379));
  OAI21_X1  g193(.A(KEYINPUT3), .B1(new_n379), .B2(G107), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT3), .ZN(new_n381));
  INV_X1    g195(.A(G107), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n381), .A2(new_n382), .A3(G104), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n379), .A2(G107), .ZN(new_n384));
  NAND4_X1  g198(.A1(new_n380), .A2(new_n383), .A3(new_n377), .A4(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT77), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n379), .A2(G107), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n382), .A2(G104), .ZN(new_n388));
  OAI211_X1 g202(.A(new_n386), .B(G101), .C1(new_n387), .C2(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n378), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n375), .A2(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n222), .B1(new_n267), .B2(new_n250), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n230), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n393), .A2(new_n385), .A3(new_n389), .A4(new_n378), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n259), .A2(new_n258), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NOR2_X1   g211(.A1(KEYINPUT79), .A2(KEYINPUT12), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n395), .A2(new_n397), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n396), .B1(new_n391), .B2(new_n394), .ZN(new_n401));
  XOR2_X1   g215(.A(KEYINPUT79), .B(KEYINPUT12), .Z(new_n402));
  OAI21_X1  g216(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n390), .A2(KEYINPUT78), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT78), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n378), .A2(new_n405), .A3(new_n389), .A4(new_n385), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n404), .A2(KEYINPUT10), .A3(new_n231), .A4(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  AOI22_X1  g222(.A1(new_n223), .A2(G128), .B1(new_n219), .B2(new_n221), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n271), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n408), .B1(new_n390), .B2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n380), .A2(new_n383), .A3(new_n384), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(G101), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(KEYINPUT4), .A3(new_n385), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n415), .A3(G101), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n256), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n407), .A2(new_n396), .A3(new_n411), .A4(new_n417), .ZN(new_n418));
  XNOR2_X1  g232(.A(G110), .B(G140), .ZN(new_n419));
  INV_X1    g233(.A(G227), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(G953), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n419), .B(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n403), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n407), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n411), .A2(new_n417), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n397), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n423), .B1(new_n427), .B2(new_n418), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n320), .B(new_n372), .C1(new_n424), .C2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n423), .B1(new_n403), .B2(new_n418), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n418), .A2(new_n423), .ZN(new_n431));
  INV_X1    g245(.A(new_n426), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n396), .B1(new_n432), .B2(new_n407), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT80), .B1(new_n430), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n401), .A2(new_n402), .ZN(new_n436));
  AOI211_X1 g250(.A(new_n396), .B(new_n398), .C1(new_n391), .C2(new_n394), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n418), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n422), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT80), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n427), .A2(new_n418), .A3(new_n423), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n435), .B2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G469), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n429), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n234), .A2(new_n236), .A3(new_n446), .A4(G116), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n447), .A2(G113), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n237), .A2(KEYINPUT5), .A3(new_n239), .ZN(new_n449));
  INV_X1    g263(.A(new_n240), .ZN(new_n450));
  AOI22_X1  g264(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n243), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n404), .A3(new_n406), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n245), .A2(new_n414), .A3(new_n247), .A4(new_n416), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT6), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(KEYINPUT6), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n452), .B2(new_n453), .ZN(new_n461));
  OAI211_X1 g275(.A(KEYINPUT82), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n461), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT82), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n463), .A2(new_n464), .A3(KEYINPUT6), .A4(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n256), .A2(G125), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(G125), .B2(new_n375), .ZN(new_n468));
  INV_X1    g282(.A(G224), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n468), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n466), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G210), .B1(G237), .B2(G902), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n474), .A2(KEYINPUT84), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT7), .B1(new_n469), .B2(G953), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n468), .A2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n477), .ZN(new_n479));
  OAI211_X1 g293(.A(new_n467), .B(new_n479), .C1(G125), .C2(new_n375), .ZN(new_n480));
  XOR2_X1   g294(.A(new_n456), .B(KEYINPUT8), .Z(new_n481));
  NAND2_X1  g295(.A1(new_n448), .A2(new_n449), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n244), .ZN(new_n483));
  INV_X1    g297(.A(new_n390), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n481), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n451), .A2(new_n390), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n478), .A2(new_n480), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT83), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n459), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n490), .B1(new_n487), .B2(new_n488), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n473), .A2(new_n476), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n471), .B1(new_n462), .B2(new_n465), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n478), .A2(new_n480), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n485), .A2(new_n486), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n488), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n459), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n487), .A2(new_n488), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n320), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n475), .B1(new_n494), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n493), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT9), .B(G234), .ZN(new_n503));
  OAI21_X1  g317(.A(G221), .B1(new_n503), .B2(G902), .ZN(new_n504));
  OAI21_X1  g318(.A(G214), .B1(G237), .B2(G902), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n445), .A2(new_n502), .A3(new_n504), .A4(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n379), .ZN(new_n508));
  INV_X1    g322(.A(G237), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n509), .A2(new_n356), .A3(G214), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT85), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n510), .A2(new_n511), .A3(new_n220), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n188), .B(G214), .C1(KEYINPUT85), .C2(G143), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT18), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(new_n203), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n514), .A2(KEYINPUT18), .A3(G131), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n328), .A2(G146), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(new_n331), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT86), .B1(new_n514), .B2(G131), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT86), .ZN(new_n523));
  AOI211_X1 g337(.A(new_n523), .B(new_n203), .C1(new_n512), .C2(new_n513), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT17), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n348), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(KEYINPUT88), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n522), .ZN(new_n528));
  INV_X1    g342(.A(new_n524), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n515), .A2(new_n203), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n528), .A2(new_n529), .A3(new_n530), .A4(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT88), .B1(new_n525), .B2(new_n526), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n508), .B(new_n521), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT19), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n330), .B(new_n536), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n329), .B1(new_n537), .B2(G146), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT87), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g354(.A(KEYINPUT87), .B(new_n329), .C1(new_n537), .C2(G146), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AND3_X1   g356(.A1(new_n528), .A2(new_n529), .A3(new_n531), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n521), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(new_n508), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n535), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(G475), .A2(G902), .ZN(new_n548));
  XOR2_X1   g362(.A(new_n548), .B(KEYINPUT90), .Z(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n535), .A2(new_n546), .A3(KEYINPUT89), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT89), .B1(new_n535), .B2(new_n546), .ZN(new_n553));
  NOR3_X1   g367(.A1(new_n552), .A2(new_n553), .A3(new_n549), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT20), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n521), .B1(new_n533), .B2(new_n534), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(new_n545), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n535), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(new_n320), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  NAND2_X1  g375(.A1(G234), .A2(G237), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(G952), .A3(new_n356), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n563), .B(KEYINPUT93), .ZN(new_n564));
  AND3_X1   g378(.A1(new_n562), .A2(G902), .A3(G953), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT21), .B(G898), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n564), .A2(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT92), .ZN(new_n569));
  XNOR2_X1  g383(.A(G116), .B(G122), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n571), .A2(G107), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  XNOR2_X1  g387(.A(G128), .B(G143), .ZN(new_n574));
  XNOR2_X1  g388(.A(new_n574), .B(new_n208), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n238), .A2(KEYINPUT14), .A3(G122), .ZN(new_n576));
  OAI211_X1 g390(.A(G107), .B(new_n576), .C1(new_n571), .C2(KEYINPUT14), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n575), .A3(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n319), .A2(new_n503), .A3(G953), .ZN(new_n579));
  OAI21_X1  g393(.A(KEYINPUT13), .B1(new_n220), .B2(G128), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n250), .B2(G143), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n250), .A2(G143), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n581), .A2(KEYINPUT91), .B1(KEYINPUT13), .B2(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n583), .B1(KEYINPUT91), .B2(new_n581), .ZN(new_n584));
  AND2_X1   g398(.A1(new_n584), .A2(G134), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n574), .A2(new_n208), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n570), .A2(new_n382), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n586), .B1(new_n572), .B2(new_n587), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n578), .B(new_n579), .C1(new_n585), .C2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n579), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n588), .B1(new_n584), .B2(G134), .ZN(new_n591));
  INV_X1    g405(.A(new_n578), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n590), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n589), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n594), .A2(new_n320), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n597), .B1(new_n594), .B2(new_n320), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n569), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g415(.A(new_n600), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(KEYINPUT92), .A3(new_n598), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n568), .B1(new_n601), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n556), .A2(new_n561), .A3(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n506), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n318), .A2(new_n371), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  NAND2_X1  g422(.A1(new_n445), .A2(new_n504), .ZN(new_n609));
  OAI21_X1  g423(.A(G472), .B1(new_n285), .B2(G902), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n293), .A2(new_n286), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n610), .A2(new_n367), .A3(new_n611), .A4(new_n369), .ZN(new_n612));
  OR2_X1    g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  XOR2_X1   g427(.A(new_n594), .B(KEYINPUT33), .Z(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(G478), .ZN(new_n615));
  AOI211_X1 g429(.A(G478), .B(G902), .C1(new_n589), .C2(new_n593), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n595), .A2(new_n320), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT89), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n547), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n549), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n535), .A2(new_n546), .A3(KEYINPUT89), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  AOI22_X1  g438(.A1(new_n624), .A2(KEYINPUT20), .B1(new_n547), .B2(new_n550), .ZN(new_n625));
  INV_X1    g439(.A(new_n561), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n619), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n474), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n473), .A2(new_n628), .A3(new_n492), .ZN(new_n629));
  OAI21_X1  g443(.A(new_n474), .B1(new_n494), .B2(new_n500), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n629), .A2(new_n630), .A3(new_n505), .ZN(new_n631));
  NOR4_X1   g445(.A1(new_n613), .A2(new_n568), .A3(new_n627), .A4(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT34), .B(G104), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND3_X1  g448(.A1(new_n621), .A2(new_n623), .A3(new_n550), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n635), .B1(new_n554), .B2(new_n555), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n601), .A2(new_n603), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n636), .A2(new_n561), .A3(new_n638), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n568), .A3(new_n631), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n613), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n345), .A2(new_n351), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n359), .A2(KEYINPUT36), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n368), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n367), .A2(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n649), .A2(new_n611), .A3(new_n610), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n606), .A2(new_n650), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT37), .B(G110), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G12));
  INV_X1    g467(.A(new_n609), .ZN(new_n654));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n565), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n564), .A2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n639), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n630), .A2(new_n505), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n659), .A2(new_n649), .A3(new_n629), .ZN(new_n660));
  INV_X1    g474(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n318), .A2(new_n654), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G128), .ZN(G30));
  XNOR2_X1  g477(.A(KEYINPUT96), .B(KEYINPUT39), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n657), .B(new_n664), .Z(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n654), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(KEYINPUT40), .Z(new_n668));
  AND2_X1   g482(.A1(new_n493), .A2(new_n501), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT94), .B(KEYINPUT38), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n625), .A2(new_n626), .ZN(new_n673));
  INV_X1    g487(.A(new_n261), .ZN(new_n674));
  OAI21_X1  g488(.A(new_n301), .B1(new_n674), .B2(new_n305), .ZN(new_n675));
  OR2_X1    g489(.A1(new_n675), .A2(KEYINPUT95), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(KEYINPUT95), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n676), .A2(new_n281), .A3(new_n677), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n316), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n354), .A2(new_n359), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n681), .A2(new_n352), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n320), .B1(new_n682), .B2(new_n361), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n365), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n320), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n686), .A2(new_n321), .B1(new_n368), .B2(new_n647), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n505), .A3(new_n687), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n672), .A2(new_n673), .A3(new_n637), .A4(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n668), .A2(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(KEYINPUT97), .B(G143), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n690), .B(new_n691), .ZN(G45));
  INV_X1    g506(.A(new_n657), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n619), .B(new_n693), .C1(new_n625), .C2(new_n626), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n318), .A2(new_n654), .A3(new_n661), .A4(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT98), .B(G146), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G48));
  NOR3_X1   g512(.A1(new_n627), .A2(new_n568), .A3(new_n631), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n427), .A2(new_n418), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n422), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n403), .A2(new_n418), .A3(new_n423), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n429), .B(new_n504), .C1(new_n703), .C2(new_n444), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n318), .A2(new_n699), .A3(new_n371), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT99), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n706), .B(new_n708), .ZN(G15));
  NAND4_X1  g523(.A1(new_n318), .A2(new_n640), .A3(new_n371), .A4(new_n705), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND4_X1  g525(.A1(new_n659), .A2(new_n649), .A3(new_n705), .A4(new_n629), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n605), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n318), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  NOR3_X1   g529(.A1(new_n673), .A2(new_n637), .A3(new_n631), .ZN(new_n716));
  OAI22_X1  g530(.A1(new_n290), .A2(new_n291), .B1(new_n192), .B2(new_n306), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n286), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n610), .A2(new_n718), .ZN(new_n719));
  NOR4_X1   g533(.A1(new_n719), .A2(new_n370), .A3(new_n568), .A4(new_n704), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n716), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR2_X1   g536(.A1(new_n719), .A2(new_n687), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n631), .A2(new_n704), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n695), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(new_n326), .ZN(G27));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n727), .B1(new_n288), .B2(new_n294), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT101), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(new_n312), .A3(new_n729), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n439), .A2(G469), .A3(new_n441), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n439), .A2(KEYINPUT100), .A3(G469), .A4(new_n441), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n444), .A2(new_n320), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n736), .B1(new_n703), .B2(new_n372), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n504), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n493), .A2(new_n501), .A3(new_n505), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n695), .A2(new_n730), .A3(new_n741), .A4(new_n371), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT42), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n694), .A2(KEYINPUT42), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n318), .A2(new_n744), .A3(new_n371), .A4(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n203), .ZN(G33));
  AND3_X1   g561(.A1(new_n318), .A2(new_n371), .A3(new_n741), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n658), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  NAND2_X1  g564(.A1(new_n615), .A2(new_n618), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n625), .A2(new_n751), .A3(new_n626), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT102), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n754));
  OR2_X1    g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n687), .B1(new_n611), .B2(new_n610), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n755), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT104), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n504), .ZN(new_n764));
  INV_X1    g578(.A(new_n429), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n439), .A2(KEYINPUT45), .A3(new_n441), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n435), .A2(new_n442), .ZN(new_n767));
  OAI211_X1 g581(.A(G469), .B(new_n766), .C1(new_n767), .C2(KEYINPUT45), .ZN(new_n768));
  INV_X1    g582(.A(new_n736), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT46), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n765), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n769), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n764), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n666), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n740), .B(KEYINPUT103), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n759), .A2(KEYINPUT104), .A3(new_n760), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n759), .A2(new_n760), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n763), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G137), .ZN(G39));
  XNOR2_X1  g595(.A(new_n774), .B(KEYINPUT47), .ZN(new_n782));
  OR4_X1    g596(.A1(new_n318), .A2(new_n371), .A3(new_n694), .A4(new_n740), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT105), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NOR3_X1   g599(.A1(new_n318), .A2(new_n371), .A3(new_n740), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n786), .A2(KEYINPUT105), .A3(new_n695), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G140), .ZN(G42));
  OAI21_X1  g603(.A(new_n429), .B1(new_n703), .B2(new_n444), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n791), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(KEYINPUT106), .B2(KEYINPUT49), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n796));
  AND4_X1   g610(.A1(new_n504), .A2(new_n795), .A3(new_n505), .A4(new_n796), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n680), .A2(new_n370), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n797), .A2(new_n672), .A3(new_n752), .A4(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n564), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n755), .A2(new_n800), .A3(new_n757), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT111), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n755), .A2(KEYINPUT111), .A3(new_n800), .A4(new_n757), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n719), .A2(new_n370), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n671), .A2(new_n505), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n805), .A2(new_n705), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT114), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT115), .A3(KEYINPUT50), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT115), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n808), .B2(KEYINPUT114), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT50), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n808), .B2(new_n811), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n810), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n740), .A2(new_n704), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n798), .A2(new_n800), .A3(new_n816), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n817), .A2(new_n673), .A3(new_n751), .ZN(new_n818));
  INV_X1    g632(.A(new_n816), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n803), .B2(new_n804), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT116), .ZN(new_n821));
  AND3_X1   g635(.A1(new_n820), .A2(new_n821), .A3(new_n723), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n821), .B1(new_n820), .B2(new_n723), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n806), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n803), .B2(new_n804), .ZN(new_n826));
  INV_X1    g640(.A(new_n776), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n790), .A2(KEYINPUT112), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(new_n764), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n826), .B(new_n827), .C1(new_n782), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT51), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n824), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n815), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n356), .A2(G952), .ZN(new_n836));
  INV_X1    g650(.A(new_n627), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n817), .B2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT48), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n730), .A2(new_n371), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n820), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n820), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n826), .A2(new_n629), .A3(new_n659), .A4(new_n705), .ZN(new_n844));
  OR2_X1    g658(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(KEYINPUT117), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g661(.A(new_n830), .B(KEYINPUT113), .ZN(new_n848));
  OAI211_X1 g662(.A(new_n826), .B(new_n827), .C1(new_n782), .C2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n849), .B(new_n818), .C1(new_n822), .C2(new_n823), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n809), .A2(KEYINPUT115), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n808), .A2(new_n811), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT50), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n850), .B1(new_n854), .B2(new_n810), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n835), .B(new_n847), .C1(new_n855), .C2(KEYINPUT51), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n857));
  AOI22_X1  g671(.A1(new_n318), .A2(new_n713), .B1(new_n716), .B2(new_n720), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n706), .A3(new_n710), .ZN(new_n859));
  INV_X1    g673(.A(new_n568), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n502), .A2(new_n860), .A3(new_n505), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n861), .A2(new_n609), .A3(new_n612), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n556), .A2(new_n561), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT107), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n599), .B2(new_n600), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n602), .A2(KEYINPUT107), .A3(new_n598), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n627), .B1(new_n863), .B2(new_n867), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n862), .A2(new_n868), .B1(new_n606), .B2(new_n650), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT108), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n657), .B1(new_n865), .B2(new_n866), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n636), .A2(new_n870), .A3(new_n561), .A4(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n740), .A2(new_n687), .ZN(new_n873));
  AND2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n636), .A2(new_n561), .A3(new_n871), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT108), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n318), .A2(new_n874), .A3(new_n654), .A4(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n869), .A2(new_n877), .A3(new_n607), .ZN(new_n878));
  NOR3_X1   g692(.A1(new_n694), .A2(new_n687), .A3(new_n719), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n741), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n295), .A2(new_n309), .A3(KEYINPUT73), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n313), .B1(new_n312), .B2(new_n316), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n371), .B(new_n741), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n658), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n880), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NOR4_X1   g699(.A1(new_n859), .A2(new_n878), .A3(new_n746), .A4(new_n885), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n879), .A2(new_n724), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n649), .A2(new_n764), .A3(new_n657), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n716), .A2(new_n738), .A3(new_n680), .A4(new_n888), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n662), .A2(new_n696), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT52), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n890), .B(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(new_n892), .A3(KEYINPUT53), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n609), .B(new_n660), .C1(new_n310), .C2(new_n317), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n725), .B1(new_n895), .B2(new_n658), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n896), .A2(new_n891), .A3(new_n696), .A4(new_n889), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n890), .A2(KEYINPUT52), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n878), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n858), .A2(new_n706), .A3(new_n710), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n743), .A2(new_n745), .ZN(new_n902));
  INV_X1    g716(.A(new_n885), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n900), .A2(new_n901), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n894), .B1(new_n899), .B2(new_n904), .ZN(new_n905));
  AOI211_X1 g719(.A(KEYINPUT109), .B(new_n857), .C1(new_n893), .C2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT109), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n893), .A2(new_n905), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n907), .B1(new_n908), .B2(KEYINPUT54), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n901), .A2(new_n902), .A3(KEYINPUT110), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT110), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n859), .B2(new_n746), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n878), .A2(new_n885), .A3(new_n894), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n892), .A2(new_n910), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n857), .A3(new_n905), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n906), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n856), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(G952), .A2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n799), .B1(new_n917), .B2(new_n918), .ZN(G75));
  NOR2_X1   g733(.A1(new_n356), .A2(G952), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT118), .Z(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n914), .A2(new_n905), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(G902), .ZN(new_n925));
  INV_X1    g739(.A(G210), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n466), .B(new_n472), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT55), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  OR2_X1    g744(.A1(new_n927), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n927), .A2(new_n930), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n922), .B1(new_n931), .B2(new_n932), .ZN(G51));
  XNOR2_X1  g747(.A(new_n736), .B(KEYINPUT57), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n914), .A2(new_n857), .A3(new_n905), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n857), .B1(new_n914), .B2(new_n905), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n701), .A2(new_n702), .ZN(new_n940));
  OAI211_X1 g754(.A(KEYINPUT119), .B(new_n934), .C1(new_n935), .C2(new_n936), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n925), .A2(new_n768), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n920), .B1(new_n942), .B2(new_n943), .ZN(G54));
  INV_X1    g758(.A(new_n925), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n552), .A2(new_n553), .ZN(new_n946));
  NAND2_X1  g760(.A1(KEYINPUT58), .A2(G475), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT120), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n945), .A2(new_n946), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n946), .B1(new_n945), .B2(new_n948), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n920), .ZN(G60));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n614), .B(KEYINPUT121), .Z(new_n953));
  XOR2_X1   g767(.A(new_n617), .B(KEYINPUT59), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT53), .B1(new_n886), .B2(new_n892), .ZN(new_n956));
  NAND3_X1  g770(.A1(new_n910), .A2(new_n913), .A3(new_n912), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n957), .A2(new_n899), .ZN(new_n958));
  OAI21_X1  g772(.A(KEYINPUT54), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n959), .B2(new_n915), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n952), .B1(new_n960), .B2(new_n922), .ZN(new_n961));
  INV_X1    g775(.A(new_n955), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n935), .B2(new_n936), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(KEYINPUT122), .A3(new_n921), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n961), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n953), .B1(new_n916), .B2(new_n954), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT60), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n969), .B1(new_n914), .B2(new_n905), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n647), .ZN(new_n971));
  NOR2_X1   g785(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n922), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n971), .B(new_n973), .C1(new_n363), .C2(new_n970), .ZN(new_n974));
  NAND2_X1  g788(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n974), .B(new_n975), .ZN(G66));
  OAI21_X1  g790(.A(G953), .B1(new_n566), .B2(new_n469), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n869), .A2(new_n607), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n859), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n977), .B1(new_n979), .B2(G953), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n462), .B(new_n465), .C1(G898), .C2(new_n356), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(G69));
  OR2_X1    g796(.A1(new_n277), .A2(new_n278), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n983), .B(new_n537), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT125), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n840), .A2(new_n716), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n902), .B(new_n749), .C1(new_n775), .C2(new_n987), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n662), .A2(new_n696), .A3(new_n887), .ZN(new_n989));
  OR2_X1    g803(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n989), .A2(KEYINPUT124), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n780), .A2(new_n788), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n356), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n356), .A2(G900), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n986), .B1(new_n995), .B2(new_n997), .ZN(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n992), .B2(new_n993), .ZN(new_n999));
  NOR3_X1   g813(.A1(new_n999), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n985), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n990), .A2(new_n991), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n1002), .A2(new_n690), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT62), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1002), .A2(new_n1005), .A3(new_n690), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n667), .A2(new_n740), .ZN(new_n1007));
  NAND4_X1  g821(.A1(new_n1007), .A2(new_n318), .A3(new_n371), .A4(new_n868), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .A4(new_n993), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n356), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n984), .ZN(new_n1011));
  OAI221_X1 g825(.A(G953), .B1(new_n420), .B2(new_n655), .C1(new_n984), .C2(KEYINPUT126), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1001), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g827(.A(new_n1012), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n995), .A2(new_n986), .A3(new_n997), .ZN(new_n1015));
  OAI21_X1  g829(.A(KEYINPUT125), .B1(new_n999), .B2(new_n996), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n984), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n985), .B1(new_n1009), .B2(new_n356), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1013), .A2(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  INV_X1    g836(.A(new_n979), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1022), .B1(new_n994), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n297), .A2(new_n192), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n920), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n908), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n299), .A2(new_n302), .A3(new_n281), .ZN(new_n1028));
  NAND2_X1  g842(.A1(new_n1028), .A2(new_n1022), .ZN(new_n1029));
  XNOR2_X1  g843(.A(new_n1029), .B(KEYINPUT127), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1026), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1022), .B1(new_n1009), .B2(new_n1023), .ZN(new_n1032));
  NOR2_X1   g846(.A1(new_n298), .A2(new_n301), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(G57));
endmodule


