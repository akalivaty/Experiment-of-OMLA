//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:48 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n790, new_n791, new_n792, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  INV_X1    g004(.A(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT76), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n193), .A2(KEYINPUT76), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  XOR2_X1   g012(.A(KEYINPUT24), .B(G110), .Z(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT77), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n193), .B1(new_n201), .B2(KEYINPUT23), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n195), .A2(KEYINPUT23), .ZN(new_n203));
  OAI21_X1  g017(.A(KEYINPUT77), .B1(new_n192), .B2(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n202), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G110), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n200), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G140), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G125), .ZN(new_n209));
  INV_X1    g023(.A(G125), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G140), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n211), .A3(KEYINPUT16), .ZN(new_n212));
  OR3_X1    g026(.A1(new_n210), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n212), .A2(new_n213), .A3(KEYINPUT78), .A4(G146), .ZN(new_n214));
  AOI21_X1  g028(.A(G146), .B1(new_n212), .B2(new_n213), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT78), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n213), .A3(G146), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n215), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n207), .B1(new_n214), .B2(new_n218), .ZN(new_n219));
  OAI22_X1  g033(.A1(new_n198), .A2(new_n199), .B1(new_n205), .B2(G110), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT64), .A2(G146), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(KEYINPUT64), .A2(G146), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(new_n209), .A3(new_n211), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n220), .A2(new_n217), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n191), .B1(new_n219), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n214), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n228), .A2(new_n200), .A3(new_n206), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n220), .A2(new_n217), .A3(new_n225), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n229), .A2(new_n230), .A3(new_n190), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT75), .B(G902), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT25), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n227), .A2(new_n231), .A3(KEYINPUT25), .A4(new_n232), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(G217), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n232), .B2(G234), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n239), .A2(G902), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n227), .A2(new_n231), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  XOR2_X1   g058(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XOR2_X1   g061(.A(new_n247), .B(KEYINPUT27), .Z(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT26), .B(G101), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g064(.A(KEYINPUT28), .ZN(new_n251));
  INV_X1    g065(.A(G137), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n252), .A2(KEYINPUT11), .A3(G134), .ZN(new_n253));
  INV_X1    g067(.A(G134), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G137), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT66), .B(G131), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT11), .ZN(new_n258));
  OAI211_X1 g072(.A(KEYINPUT65), .B(new_n258), .C1(new_n254), .C2(G137), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n252), .A2(G134), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT65), .B1(new_n261), .B2(new_n258), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n256), .B(new_n257), .C1(new_n260), .C2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n253), .A2(new_n255), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n258), .B1(new_n254), .B2(G137), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n266), .B1(new_n269), .B2(new_n259), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(KEYINPUT67), .A3(new_n257), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT64), .ZN(new_n273));
  INV_X1    g087(.A(G146), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n275), .A2(G143), .A3(new_n221), .ZN(new_n276));
  INV_X1    g090(.A(G143), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G146), .ZN(new_n278));
  INV_X1    g092(.A(G128), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(KEYINPUT1), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n279), .B1(new_n276), .B2(KEYINPUT1), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n274), .A2(G143), .ZN(new_n283));
  INV_X1    g097(.A(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n275), .A2(new_n221), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n284), .B1(new_n285), .B2(new_n277), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n281), .B1(new_n282), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n261), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n290));
  OAI21_X1  g104(.A(G131), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n272), .A2(new_n287), .A3(new_n291), .ZN(new_n292));
  OR2_X1    g106(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n293));
  INV_X1    g107(.A(G131), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n270), .B2(KEYINPUT68), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n293), .A2(new_n295), .B1(new_n265), .B2(new_n271), .ZN(new_n296));
  AND2_X1   g110(.A1(KEYINPUT0), .A2(G128), .ZN(new_n297));
  NOR2_X1   g111(.A1(KEYINPUT0), .A2(G128), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G143), .B1(new_n275), .B2(new_n221), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n284), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n276), .A2(new_n278), .A3(new_n297), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n292), .B1(new_n296), .B2(new_n303), .ZN(new_n304));
  XNOR2_X1  g118(.A(KEYINPUT70), .B(G116), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G119), .ZN(new_n306));
  INV_X1    g120(.A(G116), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n306), .B1(new_n307), .B2(G119), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT2), .B(G113), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n309), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n306), .B(new_n311), .C1(new_n307), .C2(G119), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n251), .B1(new_n304), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n304), .A2(new_n313), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  AND3_X1   g130(.A1(new_n272), .A2(new_n287), .A3(new_n291), .ZN(new_n317));
  OAI21_X1  g131(.A(KEYINPUT71), .B1(new_n296), .B2(new_n303), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n263), .A2(new_n264), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT67), .B1(new_n270), .B2(new_n257), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n256), .B(KEYINPUT68), .C1(new_n260), .C2(new_n262), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(G131), .ZN(new_n322));
  NOR2_X1   g136(.A1(new_n270), .A2(KEYINPUT68), .ZN(new_n323));
  OAI22_X1  g137(.A1(new_n319), .A2(new_n320), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT71), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n301), .A2(new_n302), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n317), .B1(new_n318), .B2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n313), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT28), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n250), .B1(new_n316), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n318), .A2(new_n327), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n329), .A3(new_n292), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT30), .ZN(new_n334));
  AOI211_X1 g148(.A(new_n334), .B(new_n317), .C1(new_n318), .C2(new_n327), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n304), .A2(new_n334), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n313), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n250), .B(new_n333), .C1(new_n335), .C2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT31), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NOR3_X1   g154(.A1(new_n296), .A2(KEYINPUT71), .A3(new_n303), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n325), .B1(new_n324), .B2(new_n326), .ZN(new_n342));
  OAI211_X1 g156(.A(KEYINPUT30), .B(new_n292), .C1(new_n341), .C2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n329), .B1(new_n304), .B2(new_n334), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n343), .A2(new_n344), .B1(new_n328), .B2(new_n329), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(KEYINPUT31), .A3(new_n250), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n331), .B1(new_n340), .B2(new_n346), .ZN(new_n347));
  NOR2_X1   g161(.A1(G472), .A2(G902), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n245), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(new_n331), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n343), .A2(new_n344), .ZN(new_n352));
  AND4_X1   g166(.A1(KEYINPUT31), .A2(new_n352), .A3(new_n250), .A4(new_n333), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT31), .B1(new_n345), .B2(new_n250), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n351), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT32), .A3(new_n348), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n350), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G472), .ZN(new_n358));
  INV_X1    g172(.A(new_n232), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT74), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n329), .B1(new_n332), .B2(new_n292), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n313), .B(new_n317), .C1(new_n318), .C2(new_n327), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n360), .B(KEYINPUT28), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n292), .B1(new_n341), .B2(new_n342), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n313), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n251), .B1(new_n365), .B2(new_n333), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n314), .A2(KEYINPUT74), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n250), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT29), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n359), .B1(new_n368), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n345), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT73), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n369), .ZN(new_n375));
  OAI21_X1  g189(.A(KEYINPUT73), .B1(new_n345), .B2(new_n250), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n316), .A2(new_n250), .A3(new_n330), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n375), .A2(new_n376), .A3(new_n370), .A4(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n358), .B1(new_n372), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n244), .B1(new_n357), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G221), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT9), .B(G234), .ZN(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G902), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n381), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT3), .B1(new_n386), .B2(G107), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT3), .ZN(new_n388));
  INV_X1    g202(.A(G107), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G104), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n386), .A2(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n387), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AND2_X1   g206(.A1(new_n392), .A2(G101), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n387), .A2(new_n390), .A3(new_n394), .A4(new_n391), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT79), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT4), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n393), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n392), .A2(G101), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT79), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT4), .A4(new_n395), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n397), .A2(new_n326), .A3(new_n399), .A4(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT80), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n395), .ZN(new_n405));
  AOI22_X1  g219(.A1(new_n405), .A2(KEYINPUT79), .B1(new_n398), .B2(new_n393), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT80), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n326), .A4(new_n402), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n391), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n386), .A2(G107), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n395), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT81), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT81), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n395), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n287), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(KEYINPUT10), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n276), .A2(new_n278), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n279), .B1(new_n283), .B2(KEYINPUT1), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n281), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  INV_X1    g236(.A(new_n413), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n421), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n409), .A2(new_n296), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n276), .A2(KEYINPUT1), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G128), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n283), .B1(new_n224), .B2(G143), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n430), .A2(new_n281), .A3(new_n413), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n421), .A2(new_n423), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n324), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT12), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n324), .A3(KEYINPUT12), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n426), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G110), .B(G140), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n188), .A2(G227), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n440), .B(new_n441), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n404), .A2(new_n408), .B1(new_n418), .B2(new_n424), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n442), .B1(new_n443), .B2(new_n296), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n409), .A2(new_n425), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n324), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n439), .A2(new_n442), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(G469), .B1(new_n447), .B2(G902), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT82), .ZN(new_n449));
  INV_X1    g263(.A(G469), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n443), .A2(new_n296), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n409), .A2(new_n296), .A3(new_n425), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n442), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n444), .A2(new_n438), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n359), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n439), .A2(new_n442), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n444), .A2(new_n446), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n450), .B1(new_n459), .B2(new_n384), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT82), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n385), .B1(new_n456), .B2(new_n461), .ZN(new_n462));
  OAI21_X1  g276(.A(G214), .B1(G237), .B2(G902), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n303), .B2(G125), .ZN(new_n466));
  AOI211_X1 g280(.A(KEYINPUT84), .B(new_n210), .C1(new_n301), .C2(new_n302), .ZN(new_n467));
  OR2_X1    g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  OAI211_X1 g282(.A(new_n210), .B(new_n281), .C1(new_n282), .C2(new_n286), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT85), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n469), .B(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT7), .ZN(new_n472));
  INV_X1    g286(.A(G224), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G953), .ZN(new_n474));
  OAI22_X1  g288(.A1(new_n468), .A2(new_n471), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT86), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI221_X1 g291(.A(KEYINPUT86), .B1(new_n472), .B2(new_n474), .C1(new_n468), .C2(new_n471), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n466), .A2(new_n467), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n430), .A2(new_n470), .A3(new_n210), .A4(new_n281), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n469), .A2(KEYINPUT85), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n474), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n480), .A2(new_n483), .A3(KEYINPUT7), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n192), .A3(G116), .ZN(new_n487));
  OAI211_X1 g301(.A(G113), .B(new_n487), .C1(new_n308), .C2(new_n486), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(new_n312), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n423), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n312), .A3(new_n413), .ZN(new_n491));
  XNOR2_X1  g305(.A(G110), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT8), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n406), .A2(new_n313), .A3(new_n402), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n488), .A2(new_n312), .A3(new_n414), .A4(new_n416), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(new_n496), .A3(new_n492), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n485), .A2(new_n494), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n479), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n495), .A2(new_n496), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n492), .B(KEYINPUT83), .Z(new_n501));
  AOI22_X1  g315(.A1(new_n497), .A2(KEYINPUT6), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n500), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n468), .A2(new_n471), .A3(new_n474), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n484), .B1(new_n480), .B2(new_n483), .ZN(new_n505));
  OAI22_X1  g319(.A1(new_n502), .A2(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(new_n384), .A3(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(G210), .B1(G237), .B2(G902), .ZN(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(G902), .B1(new_n479), .B2(new_n498), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n508), .A3(new_n506), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n464), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT20), .ZN(new_n514));
  NOR2_X1   g328(.A1(G475), .A2(G902), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n515), .B(KEYINPUT88), .Z(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n257), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(G143), .B1(new_n246), .B2(G214), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n518), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n523));
  INV_X1    g337(.A(G237), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n188), .A3(G214), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n277), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n257), .A3(new_n519), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n519), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n529), .A2(KEYINPUT17), .A3(new_n518), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n218), .A2(new_n528), .A3(new_n214), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G113), .B(G122), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n532), .B(new_n386), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n209), .A2(new_n211), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n534), .A2(G146), .ZN(new_n535));
  NAND2_X1  g349(.A1(KEYINPUT18), .A2(G131), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  AOI22_X1  g351(.A1(new_n225), .A2(new_n535), .B1(new_n529), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n520), .A2(new_n521), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT87), .B1(new_n539), .B2(new_n536), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT87), .ZN(new_n541));
  NOR3_X1   g355(.A1(new_n529), .A2(new_n541), .A3(new_n537), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n538), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n531), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n522), .A2(new_n527), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n534), .B(KEYINPUT19), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(new_n217), .C1(new_n285), .C2(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n533), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n514), .B(new_n517), .C1(new_n544), .C2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT89), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n544), .A2(new_n548), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT20), .B1(new_n552), .B2(new_n516), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n531), .A2(new_n533), .A3(new_n543), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n543), .A2(new_n547), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n554), .B1(new_n555), .B2(new_n533), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(KEYINPUT89), .A3(new_n514), .A4(new_n517), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n551), .A2(new_n553), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n533), .B1(new_n531), .B2(new_n543), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n384), .B1(new_n544), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G475), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n558), .A2(KEYINPUT90), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT90), .B1(new_n558), .B2(new_n561), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(G478), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT15), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n565), .B1(KEYINPUT94), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n567), .B1(KEYINPUT94), .B2(new_n566), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n307), .A2(KEYINPUT70), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT70), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G116), .ZN(new_n571));
  AND3_X1   g385(.A1(new_n569), .A2(new_n571), .A3(G122), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT91), .ZN(new_n573));
  INV_X1    g387(.A(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(KEYINPUT91), .A2(G122), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n307), .B1(new_n575), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g391(.A(G107), .B1(new_n572), .B2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n576), .ZN(new_n579));
  NOR2_X1   g393(.A1(KEYINPUT91), .A2(G122), .ZN(new_n580));
  OAI21_X1  g394(.A(G116), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n569), .A2(new_n571), .A3(G122), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n389), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n578), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n277), .A2(G128), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n279), .A2(G143), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n585), .A2(new_n586), .A3(new_n254), .ZN(new_n587));
  XNOR2_X1  g401(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n586), .B1(new_n588), .B2(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n585), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n588), .A2(KEYINPUT93), .A3(new_n585), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n589), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n584), .B(new_n587), .C1(new_n594), .C2(new_n254), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n582), .A2(KEYINPUT14), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT14), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n305), .A2(new_n597), .A3(G122), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n598), .A3(new_n581), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G107), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n585), .A2(new_n586), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(G134), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n587), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n583), .A3(new_n603), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n382), .A2(new_n238), .A3(G953), .ZN(new_n605));
  AND3_X1   g419(.A1(new_n595), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n605), .B1(new_n595), .B2(new_n604), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n232), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT95), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n592), .A2(new_n593), .ZN(new_n611));
  INV_X1    g425(.A(new_n589), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n254), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n583), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n389), .B1(new_n581), .B2(new_n582), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n587), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n577), .B1(KEYINPUT14), .B2(new_n582), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n389), .B1(new_n617), .B2(new_n598), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n603), .A2(new_n583), .ZN(new_n619));
  OAI22_X1  g433(.A1(new_n613), .A2(new_n616), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n605), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n595), .A2(new_n604), .A3(new_n605), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n624), .A2(KEYINPUT95), .A3(new_n232), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n568), .B1(new_n610), .B2(new_n625), .ZN(new_n626));
  AOI21_X1  g440(.A(KEYINPUT95), .B1(new_n624), .B2(new_n232), .ZN(new_n627));
  INV_X1    g441(.A(new_n568), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(KEYINPUT96), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  AOI211_X1 g444(.A(new_n609), .B(new_n359), .C1(new_n622), .C2(new_n623), .ZN(new_n631));
  OAI21_X1  g445(.A(new_n628), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n610), .A2(new_n568), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n188), .A2(G952), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n637), .B1(G234), .B2(G237), .ZN(new_n638));
  AOI211_X1 g452(.A(new_n188), .B(new_n232), .C1(G234), .C2(G237), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT21), .B(G898), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n638), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n564), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n462), .A2(new_n513), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n380), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(new_n394), .ZN(G3));
  NAND2_X1  g460(.A1(new_n355), .A2(new_n232), .ZN(new_n647));
  AOI22_X1  g461(.A1(new_n647), .A2(G472), .B1(new_n348), .B2(new_n355), .ZN(new_n648));
  AND3_X1   g462(.A1(new_n648), .A2(new_n244), .A3(new_n462), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n608), .A2(new_n565), .ZN(new_n650));
  INV_X1    g464(.A(new_n620), .ZN(new_n651));
  OAI21_X1  g465(.A(KEYINPUT33), .B1(new_n651), .B2(KEYINPUT97), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(new_n624), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n232), .A2(G478), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n650), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n655), .B1(new_n562), .B2(new_n563), .ZN(new_n656));
  INV_X1    g470(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n649), .A2(new_n513), .A3(new_n642), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT34), .B(G104), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G6));
  AND4_X1   g474(.A1(new_n384), .A2(new_n499), .A3(new_n508), .A4(new_n506), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n508), .B1(new_n511), .B2(new_n506), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n463), .B(new_n642), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n553), .A2(new_n549), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n630), .A2(new_n635), .A3(new_n561), .A4(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n649), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT98), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT35), .B(G107), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G9));
  NAND2_X1  g484(.A1(new_n229), .A2(new_n230), .ZN(new_n671));
  OR2_X1    g485(.A1(new_n191), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n241), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n675), .B1(new_n237), .B2(new_n239), .ZN(new_n676));
  AOI211_X1 g490(.A(new_n464), .B(new_n676), .C1(new_n510), .C2(new_n512), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n648), .A2(new_n462), .A3(new_n643), .A4(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(G900), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n638), .B1(new_n639), .B2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n514), .B1(new_n556), .B2(new_n517), .ZN(new_n684));
  INV_X1    g498(.A(new_n549), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n561), .B(new_n683), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n630), .A2(new_n635), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT99), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n357), .B2(new_n379), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n462), .A2(new_n677), .ZN(new_n691));
  OAI21_X1  g505(.A(KEYINPUT100), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n350), .A2(new_n356), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n372), .A2(new_n378), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(G472), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n448), .A2(new_n449), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n453), .A2(new_n454), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n450), .A3(new_n232), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n461), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n385), .ZN(new_n701));
  AND3_X1   g515(.A1(new_n677), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT100), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n696), .A2(new_n702), .A3(new_n703), .A4(new_n689), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n692), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G128), .ZN(G30));
  XOR2_X1   g520(.A(new_n682), .B(KEYINPUT39), .Z(new_n707));
  NAND2_X1  g521(.A1(new_n462), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g522(.A(new_n708), .B(KEYINPUT40), .Z(new_n709));
  NAND3_X1  g523(.A1(new_n365), .A2(new_n369), .A3(new_n333), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(new_n384), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n345), .A2(new_n369), .ZN(new_n712));
  OAI21_X1  g526(.A(G472), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n350), .A2(new_n356), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT101), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n630), .A2(new_n635), .A3(new_n463), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n564), .A2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  INV_X1    g533(.A(new_n676), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n510), .A2(new_n512), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(KEYINPUT38), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(KEYINPUT102), .B1(new_n717), .B2(new_n676), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n721), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n709), .A2(new_n715), .A3(new_n726), .ZN(new_n727));
  XOR2_X1   g541(.A(KEYINPUT103), .B(G143), .Z(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G45));
  OAI211_X1 g543(.A(new_n655), .B(new_n683), .C1(new_n562), .C2(new_n563), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n731), .B1(new_n357), .B2(new_n379), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n691), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(new_n274), .ZN(G48));
  INV_X1    g548(.A(new_n442), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n735), .B1(new_n446), .B2(new_n426), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n426), .A2(new_n438), .A3(new_n735), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n232), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(G469), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n699), .A3(new_n701), .ZN(new_n740));
  NOR3_X1   g554(.A1(new_n663), .A2(new_n740), .A3(new_n656), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n741), .B(new_n244), .C1(new_n357), .C2(new_n379), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  NOR3_X1   g558(.A1(new_n663), .A2(new_n740), .A3(new_n665), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n745), .B(new_n244), .C1(new_n357), .C2(new_n379), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  OAI211_X1 g561(.A(new_n463), .B(new_n720), .C1(new_n661), .C2(new_n662), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(new_n740), .ZN(new_n749));
  OAI211_X1 g563(.A(new_n749), .B(new_n643), .C1(new_n357), .C2(new_n379), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  INV_X1    g565(.A(new_n740), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n717), .A2(new_n752), .A3(new_n722), .A4(new_n642), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n340), .A2(new_n346), .ZN(new_n754));
  OAI211_X1 g568(.A(new_n363), .B(new_n369), .C1(new_n366), .C2(new_n367), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n348), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n647), .A2(G472), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT104), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(new_n760), .A3(new_n348), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n758), .A2(new_n244), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI22_X1  g578(.A1(new_n757), .A2(KEYINPUT104), .B1(new_n647), .B2(G472), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n765), .A2(KEYINPUT105), .A3(new_n244), .A4(new_n761), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n753), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n574), .ZN(G24));
  NAND3_X1  g582(.A1(new_n758), .A2(new_n759), .A3(new_n761), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n749), .A2(new_n731), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT106), .B(G125), .Z(new_n772));
  XNOR2_X1  g586(.A(new_n771), .B(new_n772), .ZN(G27));
  INV_X1    g587(.A(KEYINPUT32), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n347), .B2(new_n349), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n695), .A2(new_n356), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n738), .A2(G469), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n701), .B1(new_n777), .B2(new_n460), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n510), .A2(new_n463), .A3(new_n512), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n778), .A2(new_n730), .A3(new_n779), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n776), .A2(KEYINPUT42), .A3(new_n244), .A4(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(KEYINPUT108), .B(KEYINPUT42), .ZN(new_n782));
  OAI211_X1 g596(.A(new_n780), .B(new_n244), .C1(new_n357), .C2(new_n379), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT107), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n782), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n243), .B1(new_n693), .B2(new_n695), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT107), .B1(new_n786), .B2(new_n780), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n781), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G131), .ZN(G33));
  AOI21_X1  g603(.A(new_n385), .B1(new_n699), .B2(new_n448), .ZN(new_n790));
  INV_X1    g604(.A(new_n779), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n689), .A2(new_n790), .A3(new_n791), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n792), .A2(new_n380), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(new_n254), .ZN(G36));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  INV_X1    g609(.A(new_n648), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n720), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n564), .A2(new_n655), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(KEYINPUT43), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n795), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT43), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n798), .B(new_n801), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n802), .A2(KEYINPUT44), .A3(new_n796), .A4(new_n720), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(new_n791), .A3(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n450), .A2(new_n384), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT45), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n450), .B1(new_n459), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n447), .A2(KEYINPUT45), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n805), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n777), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(KEYINPUT109), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT110), .ZN(new_n813));
  OAI21_X1  g627(.A(new_n813), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n809), .A2(new_n813), .A3(KEYINPUT46), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n811), .A2(new_n812), .A3(new_n814), .A4(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n816), .A2(new_n701), .A3(new_n707), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n804), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(new_n252), .ZN(G39));
  NOR4_X1   g633(.A1(new_n696), .A2(new_n244), .A3(new_n730), .A4(new_n779), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n816), .A2(KEYINPUT47), .A3(new_n701), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT47), .B1(new_n816), .B2(new_n701), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n820), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT111), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI211_X1 g639(.A(KEYINPUT111), .B(new_n820), .C1(new_n821), .C2(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  XOR2_X1   g641(.A(KEYINPUT112), .B(G140), .Z(new_n828));
  XNOR2_X1  g642(.A(new_n827), .B(new_n828), .ZN(G42));
  NAND2_X1  g643(.A1(new_n739), .A2(new_n699), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT113), .Z(new_n832));
  NAND2_X1  g646(.A1(new_n830), .A2(KEYINPUT49), .ZN(new_n833));
  NOR4_X1   g647(.A1(new_n798), .A2(new_n243), .A3(new_n464), .A4(new_n385), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n724), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  OR3_X1    g649(.A1(new_n715), .A2(new_n832), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n752), .A2(new_n791), .A3(new_n638), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n715), .A2(new_n243), .A3(new_n837), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n562), .A2(new_n563), .A3(new_n655), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n799), .A2(new_n837), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n841), .A2(new_n720), .A3(new_n761), .A4(new_n765), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n821), .A2(new_n822), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n739), .A2(new_n699), .A3(new_n385), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n764), .A2(new_n766), .ZN(new_n847));
  AND2_X1   g661(.A1(new_n802), .A2(new_n638), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n791), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n723), .A2(new_n463), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n847), .A2(new_n752), .A3(new_n848), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT50), .Z(new_n854));
  AOI21_X1  g668(.A(KEYINPUT51), .B1(new_n851), .B2(new_n854), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n637), .B(KEYINPUT118), .Z(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n776), .A2(new_n244), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n841), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT48), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT48), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n841), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n857), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n849), .A2(new_n513), .A3(new_n752), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n838), .A2(new_n657), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT119), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n855), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n851), .A2(KEYINPUT51), .A3(new_n854), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT117), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n869), .A2(new_n870), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n868), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT54), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT53), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n732), .A2(new_n691), .B1(new_n769), .B2(new_n770), .ZN(new_n876));
  INV_X1    g690(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n682), .B1(new_n510), .B2(new_n512), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n717), .A2(new_n676), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n350), .A2(new_n356), .A3(new_n713), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n879), .A2(KEYINPUT115), .A3(new_n880), .A4(new_n790), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT115), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n717), .A2(new_n676), .A3(new_n790), .A4(new_n878), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n882), .B1(new_n714), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n705), .A2(new_n877), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n886), .A2(KEYINPUT116), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n876), .B1(new_n704), .B2(new_n692), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n889), .B1(new_n890), .B2(new_n885), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n891), .B2(new_n887), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n632), .A2(new_n634), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n564), .A2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n663), .B1(new_n894), .B2(new_n656), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n244), .A3(new_n648), .A4(new_n462), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n742), .A2(new_n746), .A3(new_n896), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n750), .B(new_n678), .C1(new_n380), .C2(new_n644), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n767), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NOR3_X1   g713(.A1(new_n779), .A2(new_n893), .A3(new_n686), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n696), .A2(new_n462), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n765), .A2(new_n780), .A3(new_n761), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n793), .B1(new_n903), .B2(new_n720), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n899), .A2(new_n788), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT114), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n892), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n905), .A2(new_n906), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n875), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND3_X1   g724(.A1(new_n899), .A2(new_n788), .A3(new_n904), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n886), .A2(new_n887), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n890), .A2(KEYINPUT52), .A3(new_n885), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n911), .A2(new_n914), .A3(KEYINPUT53), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n874), .B1(new_n910), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT52), .B1(new_n890), .B2(new_n885), .ZN(new_n917));
  AND4_X1   g731(.A1(KEYINPUT52), .A2(new_n705), .A3(new_n877), .A4(new_n885), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n875), .B1(new_n919), .B2(new_n905), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n892), .A2(KEYINPUT53), .A3(new_n911), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n873), .A2(new_n916), .A3(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(G952), .A2(G953), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n836), .B1(new_n924), .B2(new_n925), .ZN(G75));
  INV_X1    g740(.A(KEYINPUT120), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n188), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n232), .B1(new_n920), .B2(new_n921), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT56), .B1(new_n930), .B2(new_n509), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n502), .A2(new_n503), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n504), .A2(new_n505), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n506), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(KEYINPUT55), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n929), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  AOI211_X1 g752(.A(KEYINPUT56), .B(new_n936), .C1(new_n930), .C2(new_n509), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n927), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT53), .B1(new_n911), .B2(new_n914), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n899), .A2(KEYINPUT53), .A3(new_n788), .A4(new_n904), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n886), .A2(KEYINPUT116), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(KEYINPUT52), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n942), .B1(new_n944), .B2(new_n888), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n941), .A2(new_n945), .ZN(new_n946));
  NOR3_X1   g760(.A1(new_n946), .A2(new_n232), .A3(new_n508), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n936), .B1(new_n947), .B2(KEYINPUT56), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n931), .A2(new_n937), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n948), .A2(new_n949), .A3(KEYINPUT120), .A4(new_n929), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n940), .A2(new_n950), .ZN(G51));
  XNOR2_X1  g765(.A(new_n946), .B(new_n874), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n805), .B(KEYINPUT57), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n698), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n930), .A2(new_n808), .A3(new_n807), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n928), .B1(new_n955), .B2(new_n956), .ZN(G54));
  NAND3_X1  g771(.A1(new_n930), .A2(KEYINPUT58), .A3(G475), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n958), .A2(new_n552), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n552), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n959), .A2(new_n960), .A3(new_n928), .ZN(G60));
  NOR2_X1   g775(.A1(new_n916), .A2(new_n923), .ZN(new_n962));
  NAND2_X1  g776(.A1(G478), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT59), .Z(new_n964));
  OAI21_X1  g778(.A(new_n653), .B1(new_n962), .B2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n653), .A2(new_n964), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n928), .B1(new_n952), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n965), .A2(new_n967), .ZN(G63));
  NAND2_X1  g782(.A1(G217), .A2(G902), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT60), .Z(new_n970));
  OAI21_X1  g784(.A(new_n970), .B1(new_n941), .B2(new_n945), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n227), .A2(new_n231), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n928), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT122), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n673), .B(KEYINPUT121), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n922), .A2(new_n974), .A3(new_n970), .A4(new_n975), .ZN(new_n976));
  OAI211_X1 g790(.A(new_n970), .B(new_n975), .C1(new_n941), .C2(new_n945), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n977), .A2(KEYINPUT122), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n973), .A2(new_n976), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n980));
  NOR2_X1   g794(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT124), .ZN(new_n982));
  AND3_X1   g796(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n982), .B1(new_n979), .B2(new_n980), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  OAI21_X1  g799(.A(G953), .B1(new_n640), .B2(new_n473), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n899), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n932), .B1(G898), .B2(new_n188), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  AND2_X1   g803(.A1(new_n825), .A2(new_n826), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n727), .A2(new_n890), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(KEYINPUT62), .ZN(new_n992));
  OR2_X1    g806(.A1(new_n804), .A2(new_n817), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT62), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n727), .A2(new_n994), .A3(new_n890), .ZN(new_n995));
  AOI21_X1  g809(.A(new_n779), .B1(new_n894), .B2(new_n656), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n786), .A2(new_n462), .A3(new_n707), .A4(new_n996), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n992), .A2(new_n993), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n188), .B1(new_n990), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n343), .A2(new_n336), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(new_n546), .Z(new_n1001));
  NAND2_X1  g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n993), .A2(KEYINPUT126), .A3(new_n890), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT126), .ZN(new_n1004));
  INV_X1    g818(.A(new_n890), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1004), .B1(new_n818), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1003), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(new_n788), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n858), .A2(new_n722), .A3(new_n717), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n817), .A2(new_n1009), .ZN(new_n1010));
  NOR3_X1   g824(.A1(new_n1008), .A2(new_n1010), .A3(new_n793), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n1007), .A2(new_n827), .A3(new_n188), .A4(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1001), .B1(G900), .B2(G953), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1002), .A2(KEYINPUT125), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT127), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND3_X1  g833(.A1(new_n1002), .A2(KEYINPUT127), .A3(new_n1014), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1020), .A2(new_n1017), .ZN(new_n1021));
  AOI22_X1  g835(.A1(new_n999), .A2(new_n1001), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1022));
  AOI21_X1  g836(.A(KEYINPUT127), .B1(new_n1022), .B2(KEYINPUT125), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n1024), .ZN(G72));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  OR2_X1    g841(.A1(new_n990), .A2(new_n998), .ZN(new_n1028));
  INV_X1    g842(.A(new_n899), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n928), .B1(new_n1030), .B2(new_n712), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1007), .A2(new_n827), .A3(new_n1011), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1027), .B1(new_n1032), .B2(new_n1029), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1033), .A2(new_n369), .A3(new_n345), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n910), .A2(new_n915), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n375), .A2(new_n376), .A3(new_n338), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1035), .A2(new_n1027), .A3(new_n1036), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1031), .A2(new_n1034), .A3(new_n1037), .ZN(G57));
endmodule


