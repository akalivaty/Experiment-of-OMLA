//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 0 0 0 1 1 1 1 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:45 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n964, new_n965, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020;
  INV_X1    g000(.A(KEYINPUT23), .ZN(new_n202));
  OAI21_X1  g001(.A(new_n202), .B1(G169gat), .B2(G176gat), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT25), .ZN(new_n204));
  NAND2_X1  g003(.A1(G169gat), .A2(G176gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  AND4_X1   g007(.A1(KEYINPUT66), .A2(new_n207), .A3(new_n208), .A4(KEYINPUT23), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT66), .B1(new_n210), .B2(KEYINPUT23), .ZN(new_n211));
  NOR3_X1   g010(.A1(new_n206), .A2(new_n209), .A3(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n213));
  INV_X1    g012(.A(G183gat), .ZN(new_n214));
  INV_X1    g013(.A(G190gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G183gat), .A2(G190gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n216), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n227), .A2(KEYINPUT65), .A3(new_n221), .A4(new_n216), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n224), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n214), .A2(new_n215), .A3(KEYINPUT67), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT67), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(G183gat), .B2(G190gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n219), .A2(new_n230), .A3(new_n232), .A4(new_n220), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n207), .A2(new_n208), .A3(KEYINPUT23), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n234), .A2(new_n203), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n233), .A2(new_n235), .A3(new_n205), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(KEYINPUT25), .ZN(new_n237));
  AND2_X1   g036(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n238));
  NOR2_X1   g037(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n239));
  OAI21_X1  g038(.A(new_n215), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT68), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT28), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n240), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT27), .B(G183gat), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n246), .A2(new_n241), .A3(new_n242), .A4(new_n215), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT26), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n210), .A2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n249), .A2(new_n205), .A3(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n245), .A2(new_n247), .A3(new_n217), .A4(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n229), .A2(new_n237), .A3(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(G127gat), .B(G134gat), .Z(new_n254));
  INV_X1    g053(.A(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(G120gat), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(G120gat), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n257), .B1(new_n261), .B2(new_n263), .ZN(new_n264));
  OAI211_X1 g063(.A(new_n255), .B(new_n256), .C1(new_n259), .C2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n260), .A2(G113gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n258), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(new_n256), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n258), .B2(new_n266), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n254), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n265), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G227gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n265), .A2(new_n271), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n277), .A2(new_n237), .A3(new_n229), .A4(new_n252), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(KEYINPUT32), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT71), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g081(.A(G15gat), .B(G43gat), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(G71gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(G99gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT33), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n285), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n279), .A2(KEYINPUT71), .A3(KEYINPUT32), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n282), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n278), .ZN(new_n290));
  INV_X1    g089(.A(new_n276), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  OAI211_X1 g091(.A(new_n279), .B(KEYINPUT32), .C1(new_n286), .C2(new_n285), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n289), .B2(new_n293), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT72), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n289), .A2(new_n293), .ZN(new_n297));
  INV_X1    g096(.A(new_n292), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n289), .A2(new_n292), .A3(new_n293), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AND3_X1   g101(.A1(new_n296), .A2(new_n302), .A3(KEYINPUT34), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT34), .B1(new_n296), .B2(new_n302), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT36), .ZN(new_n305));
  NOR3_X1   g104(.A1(new_n303), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT34), .ZN(new_n307));
  NOR3_X1   g106(.A1(new_n294), .A2(new_n295), .A3(KEYINPUT72), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n300), .B1(new_n299), .B2(new_n301), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n296), .A2(new_n302), .A3(KEYINPUT34), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT36), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n306), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  INV_X1    g113(.A(G218gat), .ZN(new_n315));
  INV_X1    g114(.A(G211gat), .ZN(new_n316));
  XNOR2_X1  g115(.A(G197gat), .B(G204gat), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT73), .B(G218gat), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT22), .B1(new_n318), .B2(G211gat), .ZN(new_n319));
  AND2_X1   g118(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(KEYINPUT74), .ZN(new_n321));
  OAI211_X1 g120(.A(new_n316), .B(new_n317), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(new_n322), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n319), .B(KEYINPUT74), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n316), .B1(new_n324), .B2(new_n317), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n315), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  OAI21_X1  g125(.A(new_n317), .B1(new_n320), .B2(new_n321), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(G211gat), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n328), .A2(G218gat), .A3(new_n322), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(KEYINPUT75), .A3(new_n329), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT29), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n253), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(G226gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(new_n336), .B2(new_n275), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n253), .A2(G226gat), .A3(G233gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n332), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT76), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n338), .B(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n342), .A2(new_n330), .A3(new_n337), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n340), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g143(.A(G8gat), .B(G36gat), .ZN(new_n345));
  INV_X1    g144(.A(G64gat), .ZN(new_n346));
  XNOR2_X1  g145(.A(new_n345), .B(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(G92gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(new_n314), .B1(new_n344), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT30), .ZN(new_n351));
  INV_X1    g150(.A(new_n349), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n340), .A2(KEYINPUT78), .A3(new_n343), .A4(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n340), .A2(KEYINPUT30), .A3(new_n343), .A4(new_n352), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT77), .B1(new_n344), .B2(new_n349), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n344), .A2(KEYINPUT77), .A3(new_n349), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n354), .B(new_n355), .C1(new_n356), .C2(new_n357), .ZN(new_n358));
  XNOR2_X1  g157(.A(G155gat), .B(G162gat), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT79), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  XNOR2_X1  g160(.A(G141gat), .B(G148gat), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT2), .ZN(new_n364));
  AND2_X1   g163(.A1(G155gat), .A2(G162gat), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT80), .B(G162gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G155gat), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n362), .B1(new_n369), .B2(KEYINPUT2), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(new_n359), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n367), .A2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT84), .B1(new_n372), .B2(new_n277), .ZN(new_n373));
  AOI22_X1  g172(.A1(new_n366), .A2(new_n361), .B1(new_n370), .B2(new_n359), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT84), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(new_n272), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n373), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n377), .B1(new_n374), .B2(new_n272), .ZN(new_n378));
  NAND2_X1  g177(.A1(G225gat), .A2(G233gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OR2_X1    g179(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n377), .A2(KEYINPUT4), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n372), .A2(KEYINPUT83), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n374), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT4), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(new_n272), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT87), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n382), .A2(new_n388), .A3(KEYINPUT87), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT3), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n374), .A2(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT81), .B(KEYINPUT3), .Z(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n367), .A2(new_n371), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n374), .A2(KEYINPUT82), .A3(new_n396), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n394), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n391), .A2(new_n392), .B1(new_n277), .B2(new_n401), .ZN(new_n402));
  OAI211_X1 g201(.A(KEYINPUT39), .B(new_n381), .C1(new_n402), .C2(new_n379), .ZN(new_n403));
  XOR2_X1   g202(.A(G1gat), .B(G29gat), .Z(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G57gat), .B(G85gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n394), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT82), .B1(new_n374), .B2(new_n396), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n397), .A2(new_n398), .ZN(new_n412));
  OAI211_X1 g211(.A(new_n410), .B(new_n277), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n392), .ZN(new_n414));
  AOI21_X1  g213(.A(KEYINPUT87), .B1(new_n382), .B2(new_n388), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n413), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT39), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n380), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n403), .A2(new_n409), .A3(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT40), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n378), .A2(new_n380), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT4), .B1(new_n373), .B2(new_n376), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n386), .A2(KEYINPUT4), .A3(new_n272), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n424), .A2(new_n413), .A3(new_n425), .A4(new_n379), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n426), .A2(KEYINPUT85), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT85), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n387), .B(new_n277), .C1(new_n383), .C2(new_n385), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n429), .A2(new_n423), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n380), .B1(new_n401), .B2(new_n277), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g231(.A(KEYINPUT5), .B(new_n422), .C1(new_n427), .C2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  OAI211_X1 g233(.A(new_n434), .B(new_n431), .C1(new_n414), .C2(new_n415), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n408), .ZN(new_n437));
  NAND4_X1  g236(.A1(new_n403), .A2(KEYINPUT40), .A3(new_n409), .A4(new_n418), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n358), .A2(new_n421), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n409), .B1(new_n433), .B2(new_n435), .ZN(new_n440));
  XOR2_X1   g239(.A(KEYINPUT88), .B(KEYINPUT6), .Z(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n433), .A2(new_n409), .A3(new_n435), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n442), .B1(new_n444), .B2(new_n441), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n344), .A2(KEYINPUT37), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n340), .A2(new_n447), .A3(new_n343), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n446), .A2(KEYINPUT38), .A3(new_n349), .A4(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n349), .ZN(new_n450));
  INV_X1    g249(.A(new_n339), .ZN(new_n451));
  INV_X1    g250(.A(new_n333), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT75), .B1(new_n326), .B2(new_n329), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT90), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n342), .A2(new_n337), .ZN(new_n457));
  INV_X1    g256(.A(new_n330), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT90), .B(new_n451), .C1(new_n452), .C2(new_n453), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n456), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n450), .B1(new_n461), .B2(KEYINPUT37), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n449), .B1(new_n462), .B2(KEYINPUT38), .ZN(new_n463));
  AND2_X1   g262(.A1(new_n350), .A2(new_n353), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n439), .B1(new_n445), .B2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(G22gat), .B(G50gat), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AND2_X1   g267(.A1(G228gat), .A2(G233gat), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n334), .B1(new_n412), .B2(new_n411), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n332), .A2(new_n470), .A3(new_n333), .ZN(new_n471));
  AOI21_X1  g270(.A(KEYINPUT29), .B1(new_n326), .B2(new_n329), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n374), .B1(new_n473), .B2(new_n393), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n469), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n386), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n472), .B2(new_n395), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT89), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n469), .B1(new_n458), .B2(new_n470), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT89), .B(new_n476), .C1(new_n472), .C2(new_n395), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G78gat), .B(G106gat), .ZN(new_n483));
  XOR2_X1   g282(.A(new_n483), .B(KEYINPUT31), .Z(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n475), .A2(new_n482), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n475), .B2(new_n482), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n468), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n475), .A2(new_n482), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n484), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n475), .A2(new_n482), .A3(new_n485), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(new_n467), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n488), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n466), .A2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n441), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n437), .B2(new_n443), .ZN(new_n496));
  NOR3_X1   g295(.A1(new_n496), .A2(new_n358), .A3(new_n442), .ZN(new_n497));
  INV_X1    g296(.A(new_n493), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n313), .B1(new_n494), .B2(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT35), .ZN(new_n501));
  NOR2_X1   g300(.A1(new_n303), .A2(new_n304), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n354), .A2(new_n355), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n357), .A2(new_n356), .ZN(new_n505));
  NOR2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n443), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n441), .B1(new_n507), .B2(new_n440), .ZN(new_n508));
  INV_X1    g307(.A(new_n442), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n501), .B1(new_n503), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n497), .A2(KEYINPUT35), .A3(new_n502), .A4(new_n493), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  OR2_X1    g312(.A1(new_n500), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT97), .ZN(new_n515));
  INV_X1    g314(.A(G8gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517));
  XNOR2_X1  g316(.A(G15gat), .B(G22gat), .ZN(new_n518));
  INV_X1    g317(.A(G1gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT16), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OR2_X1    g320(.A1(G15gat), .A2(G22gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(G15gat), .A2(G22gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(new_n519), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n516), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(G15gat), .A2(G22gat), .ZN(new_n526));
  NOR2_X1   g325(.A1(G15gat), .A2(G22gat), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n520), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AND4_X1   g327(.A1(KEYINPUT96), .A2(new_n524), .A3(new_n528), .A4(new_n516), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n515), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n524), .A2(new_n528), .A3(KEYINPUT96), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(G8gat), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n521), .A2(new_n516), .A3(new_n524), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT97), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n530), .A2(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT102), .ZN(new_n536));
  INV_X1    g335(.A(G57gat), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n537), .A2(G64gat), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n346), .A2(G57gat), .ZN(new_n539));
  OAI21_X1  g338(.A(KEYINPUT99), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(G71gat), .A2(G78gat), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT9), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n346), .A2(G57gat), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n537), .A2(G64gat), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT99), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n540), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G71gat), .ZN(new_n549));
  INV_X1    g348(.A(G78gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g350(.A1(new_n551), .A2(new_n541), .ZN(new_n552));
  XNOR2_X1  g351(.A(KEYINPUT100), .B(G57gat), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n544), .B1(new_n553), .B2(new_n346), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n541), .B1(new_n551), .B2(new_n542), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n548), .A2(new_n552), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT21), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n535), .A2(new_n536), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n536), .B1(new_n535), .B2(new_n557), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n548), .A2(new_n552), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n554), .A2(new_n555), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(KEYINPUT101), .B(KEYINPUT21), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NOR3_X1   g364(.A1(new_n559), .A2(new_n560), .A3(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n565), .B1(new_n559), .B2(new_n560), .ZN(new_n568));
  XNOR2_X1  g367(.A(G127gat), .B(G155gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(G231gat), .A2(G233gat), .ZN(new_n570));
  XOR2_X1   g369(.A(new_n569), .B(new_n570), .Z(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n567), .A2(new_n568), .A3(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n574));
  XNOR2_X1  g373(.A(G183gat), .B(G211gat), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n565), .ZN(new_n577));
  INV_X1    g376(.A(new_n560), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n577), .B1(new_n578), .B2(new_n558), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n571), .B1(new_n579), .B2(new_n566), .ZN(new_n580));
  AND3_X1   g379(.A1(new_n573), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n576), .B1(new_n573), .B2(new_n580), .ZN(new_n582));
  OR2_X1    g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(G190gat), .B(G218gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT104), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT8), .ZN(new_n588));
  NAND2_X1  g387(.A1(G85gat), .A2(G92gat), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(G85gat), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(new_n348), .ZN(new_n593));
  NAND3_X1  g392(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n588), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(G99gat), .B(G106gat), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT103), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n587), .B1(new_n592), .B2(new_n348), .ZN(new_n600));
  NAND4_X1  g399(.A1(new_n600), .A2(new_n596), .A3(new_n591), .A4(new_n594), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(new_n602));
  AND2_X1   g401(.A1(new_n591), .A2(new_n594), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n603), .A2(KEYINPUT103), .A3(new_n596), .A4(new_n600), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OR3_X1    g405(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n608));
  AOI22_X1  g407(.A1(new_n607), .A2(new_n608), .B1(G29gat), .B2(G36gat), .ZN(new_n609));
  INV_X1    g408(.A(G50gat), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n610), .A2(G43gat), .ZN(new_n611));
  INV_X1    g410(.A(G43gat), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(G50gat), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT15), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n611), .A2(new_n613), .A3(KEYINPUT93), .A4(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT93), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n610), .B2(G43gat), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n618), .A2(new_n614), .B1(new_n611), .B2(new_n613), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n609), .B1(new_n616), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT94), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n609), .B(KEYINPUT94), .C1(new_n616), .C2(new_n619), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n612), .A2(G50gat), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n610), .A2(G43gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT92), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n608), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g427(.A(KEYINPUT92), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n607), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(G29gat), .A2(G36gat), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n614), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n622), .A2(new_n623), .B1(new_n626), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT17), .ZN(new_n635));
  NOR2_X1   g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(KEYINPUT95), .A2(KEYINPUT17), .ZN(new_n637));
  NOR3_X1   g436(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n611), .A3(new_n613), .ZN(new_n640));
  INV_X1    g439(.A(new_n623), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT93), .B1(new_n612), .B2(G50gat), .ZN(new_n642));
  OAI22_X1  g441(.A1(KEYINPUT15), .A2(new_n642), .B1(new_n624), .B2(new_n625), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n615), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT94), .B1(new_n644), .B2(new_n609), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n640), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n636), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n639), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n606), .B1(new_n638), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT41), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n633), .A2(new_n606), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n649), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n646), .A2(new_n647), .A3(new_n639), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n633), .A2(new_n634), .A3(new_n635), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n605), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(new_n651), .B(new_n650), .C1(new_n659), .C2(new_n654), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n586), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(G134gat), .B(G162gat), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n656), .A2(new_n660), .A3(new_n586), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n663), .ZN(new_n666));
  INV_X1    g465(.A(new_n664), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n666), .B1(new_n667), .B2(new_n661), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n665), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n583), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n525), .A2(new_n529), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n638), .B2(new_n648), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT98), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n535), .B2(new_n633), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n530), .A2(new_n534), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n646), .A2(new_n675), .A3(KEYINPUT98), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G229gat), .A2(G233gat), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n672), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT18), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n677), .B1(new_n675), .B2(new_n646), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n678), .B(KEYINPUT13), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n672), .A2(new_n677), .A3(KEYINPUT18), .A4(new_n678), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n681), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(G113gat), .B(G141gat), .ZN(new_n687));
  XNOR2_X1  g486(.A(G169gat), .B(G197gat), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g488(.A(KEYINPUT91), .B(KEYINPUT11), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT12), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g493(.A1(new_n681), .A2(new_n684), .A3(new_n685), .A4(new_n692), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(G230gat), .A2(G233gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n605), .A2(new_n563), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n598), .A2(new_n601), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n556), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(KEYINPUT10), .B1(new_n698), .B2(new_n700), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n556), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT105), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n697), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n698), .A2(new_n706), .A3(new_n700), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT10), .ZN(new_n708));
  AOI22_X1  g507(.A1(new_n604), .A2(new_n602), .B1(new_n561), .B2(new_n562), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n561), .A2(new_n562), .A3(new_n699), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n708), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n605), .A2(KEYINPUT10), .A3(new_n556), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n713), .A2(KEYINPUT105), .A3(new_n697), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n705), .A2(new_n707), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(G120gat), .B(G148gat), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(new_n208), .ZN(new_n717));
  INV_X1    g516(.A(G204gat), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n717), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n715), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n719), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n707), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n696), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n670), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n514), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n445), .ZN(new_n728));
  XOR2_X1   g527(.A(KEYINPUT106), .B(G1gat), .Z(new_n729));
  XNOR2_X1  g528(.A(new_n728), .B(new_n729), .ZN(G1324gat));
  INV_X1    g529(.A(new_n727), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n358), .ZN(new_n732));
  XNOR2_X1  g531(.A(KEYINPUT16), .B(G8gat), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT107), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(KEYINPUT42), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(G8gat), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT42), .ZN(new_n737));
  OAI211_X1 g536(.A(KEYINPUT107), .B(new_n737), .C1(new_n732), .C2(new_n733), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(G1325gat));
  OAI21_X1  g538(.A(KEYINPUT108), .B1(new_n306), .B2(new_n312), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n305), .B1(new_n303), .B2(new_n304), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n310), .A2(KEYINPUT36), .A3(new_n311), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n740), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n731), .A2(G15gat), .A3(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(new_n502), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n727), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n747), .B1(G15gat), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT109), .ZN(G1326gat));
  NOR2_X1   g550(.A1(new_n727), .A2(new_n493), .ZN(new_n752));
  XOR2_X1   g551(.A(KEYINPUT43), .B(G22gat), .Z(new_n753));
  XNOR2_X1  g552(.A(new_n752), .B(new_n753), .ZN(G1327gat));
  AND2_X1   g553(.A1(new_n665), .A2(new_n668), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n583), .A2(new_n725), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n514), .A2(new_n755), .A3(new_n756), .ZN(new_n757));
  OR3_X1    g556(.A1(new_n757), .A2(G29gat), .A3(new_n445), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n758), .B(KEYINPUT45), .ZN(new_n759));
  OAI211_X1 g558(.A(KEYINPUT44), .B(new_n755), .C1(new_n500), .C2(new_n513), .ZN(new_n760));
  INV_X1    g559(.A(new_n513), .ZN(new_n761));
  OAI211_X1 g560(.A(new_n464), .B(new_n463), .C1(new_n496), .C2(new_n442), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n498), .B1(new_n762), .B2(new_n439), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n510), .A2(new_n493), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n745), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n669), .B1(new_n761), .B2(new_n765), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n760), .B(new_n756), .C1(new_n766), .C2(KEYINPUT44), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n767), .B2(new_n445), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n759), .A2(new_n768), .ZN(G1328gat));
  INV_X1    g568(.A(G36gat), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n514), .A2(new_n770), .A3(new_n755), .A4(new_n756), .ZN(new_n771));
  OR3_X1    g570(.A1(new_n771), .A2(KEYINPUT110), .A3(new_n506), .ZN(new_n772));
  OAI21_X1  g571(.A(KEYINPUT110), .B1(new_n771), .B2(new_n506), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT46), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g575(.A(G36gat), .B1(new_n767), .B2(new_n506), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(KEYINPUT46), .A3(new_n773), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n776), .A2(new_n777), .A3(new_n778), .ZN(G1329gat));
  OR3_X1    g578(.A1(new_n767), .A2(new_n612), .A3(new_n745), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(KEYINPUT111), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n612), .B1(new_n757), .B2(new_n748), .ZN(new_n784));
  NAND4_X1  g583(.A1(new_n780), .A2(new_n782), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n767), .A2(new_n612), .A3(new_n745), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n514), .A2(new_n755), .A3(new_n756), .ZN(new_n787));
  AOI21_X1  g586(.A(G43gat), .B1(new_n787), .B2(new_n502), .ZN(new_n788));
  OAI211_X1 g587(.A(KEYINPUT111), .B(new_n781), .C1(new_n786), .C2(new_n788), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n785), .A2(new_n789), .ZN(G1330gat));
  OAI21_X1  g589(.A(G50gat), .B1(new_n767), .B2(new_n493), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT48), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n787), .A2(new_n610), .A3(new_n498), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n791), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n791), .B(new_n794), .C1(new_n792), .C2(KEYINPUT48), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(G1331gat));
  NAND2_X1  g597(.A1(new_n494), .A2(new_n499), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n513), .B1(new_n799), .B2(new_n745), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n800), .A2(new_n724), .ZN(new_n801));
  NOR2_X1   g600(.A1(new_n670), .A2(new_n696), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n445), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(new_n553), .ZN(G1332gat));
  INV_X1    g605(.A(KEYINPUT49), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n803), .B(new_n358), .C1(new_n807), .C2(new_n346), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n346), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n808), .B(new_n809), .ZN(G1333gat));
  NAND3_X1  g609(.A1(new_n803), .A2(G71gat), .A3(new_n746), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n801), .A2(new_n802), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n549), .B1(new_n812), .B2(new_n748), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n814), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g614(.A1(new_n812), .A2(new_n493), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(new_n550), .ZN(G1335gat));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n583), .A2(new_n696), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  NOR4_X1   g619(.A1(new_n800), .A2(KEYINPUT51), .A3(new_n669), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT51), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n822), .B1(new_n766), .B2(new_n819), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n824), .A2(new_n592), .A3(new_n804), .A4(new_n723), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n820), .A2(new_n724), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n760), .B(new_n826), .C1(new_n766), .C2(KEYINPUT44), .ZN(new_n827));
  OAI21_X1  g626(.A(G85gat), .B1(new_n827), .B2(new_n445), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n818), .B1(new_n825), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n761), .A2(new_n765), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n830), .A2(new_n755), .A3(new_n819), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(KEYINPUT51), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n766), .A2(new_n822), .A3(new_n819), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n832), .A2(new_n804), .A3(new_n723), .A4(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n828), .B(new_n818), .C1(new_n834), .C2(G85gat), .ZN(new_n835));
  INV_X1    g634(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n829), .A2(new_n836), .ZN(G1336gat));
  OAI21_X1  g636(.A(G92gat), .B1(new_n827), .B2(new_n506), .ZN(new_n838));
  NOR2_X1   g637(.A1(new_n506), .A2(G92gat), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n832), .A2(new_n723), .A3(new_n833), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n841), .A2(new_n842), .A3(KEYINPUT52), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n838), .B(new_n840), .C1(KEYINPUT114), .C2(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(G1337gat));
  XOR2_X1   g645(.A(KEYINPUT115), .B(G99gat), .Z(new_n847));
  NAND3_X1  g646(.A1(new_n824), .A2(new_n723), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n827), .A2(new_n745), .ZN(new_n849));
  OAI22_X1  g648(.A1(new_n848), .A2(new_n748), .B1(new_n849), .B2(new_n847), .ZN(G1338gat));
  OAI21_X1  g649(.A(G106gat), .B1(new_n827), .B2(new_n493), .ZN(new_n851));
  INV_X1    g650(.A(G106gat), .ZN(new_n852));
  NAND4_X1  g651(.A1(new_n832), .A2(new_n852), .A3(new_n723), .A4(new_n833), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n851), .B1(new_n853), .B2(new_n493), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT53), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n851), .B(new_n856), .C1(new_n853), .C2(new_n493), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n855), .A2(new_n857), .ZN(G1339gat));
  NOR3_X1   g657(.A1(new_n670), .A2(new_n723), .A3(new_n696), .ZN(new_n859));
  INV_X1    g658(.A(new_n722), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT54), .ZN(new_n861));
  AOI21_X1  g660(.A(KEYINPUT105), .B1(new_n713), .B2(new_n697), .ZN(new_n862));
  AOI211_X1 g661(.A(new_n704), .B(new_n706), .C1(new_n711), .C2(new_n712), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n698), .A2(new_n700), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n702), .B1(new_n865), .B2(new_n708), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n861), .B1(new_n866), .B2(new_n706), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n721), .B1(new_n867), .B2(new_n703), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT55), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n864), .A2(new_n868), .A3(KEYINPUT55), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n872), .A2(KEYINPUT116), .ZN(new_n873));
  INV_X1    g672(.A(KEYINPUT116), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n864), .A2(new_n868), .A3(new_n874), .A4(KEYINPUT55), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n871), .A2(new_n873), .A3(new_n875), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n678), .B1(new_n672), .B2(new_n677), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n646), .A2(new_n675), .ZN(new_n878));
  AOI211_X1 g677(.A(new_n683), .B(new_n878), .C1(new_n674), .C2(new_n676), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n691), .B1(new_n877), .B2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(KEYINPUT117), .B(new_n691), .C1(new_n877), .C2(new_n879), .ZN(new_n883));
  AND3_X1   g682(.A1(new_n882), .A2(new_n695), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n755), .A2(new_n876), .A3(new_n884), .ZN(new_n885));
  AND4_X1   g684(.A1(new_n723), .A2(new_n882), .A3(new_n695), .A4(new_n883), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n886), .B1(new_n876), .B2(new_n696), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n755), .ZN(new_n888));
  INV_X1    g687(.A(new_n583), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n859), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n445), .A2(new_n358), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(new_n503), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n696), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n897), .B(new_n257), .ZN(G1340gat));
  NOR2_X1   g697(.A1(new_n895), .A2(new_n724), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n261), .A2(new_n263), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n901), .B1(new_n260), .B2(new_n899), .ZN(G1341gat));
  INV_X1    g701(.A(new_n895), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n903), .A2(new_n583), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(G127gat), .ZN(G1342gat));
  INV_X1    g704(.A(G134gat), .ZN(new_n906));
  NAND2_X1  g705(.A1(KEYINPUT118), .A2(KEYINPUT56), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n903), .A2(new_n906), .A3(new_n755), .A4(new_n907), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n908), .A2(KEYINPUT118), .A3(KEYINPUT56), .ZN(new_n909));
  OAI21_X1  g708(.A(G134gat), .B1(new_n895), .B2(new_n669), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(KEYINPUT118), .B2(KEYINPUT56), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n909), .A2(new_n910), .A3(new_n911), .ZN(G1343gat));
  INV_X1    g711(.A(KEYINPUT121), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n913), .B1(new_n746), .B2(new_n493), .ZN(new_n914));
  INV_X1    g713(.A(G141gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n745), .A2(KEYINPUT121), .A3(new_n498), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n914), .A2(new_n893), .A3(new_n915), .A4(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n917), .A2(new_n896), .ZN(new_n918));
  XNOR2_X1  g717(.A(new_n918), .B(KEYINPUT122), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n890), .A2(KEYINPUT57), .A3(new_n493), .ZN(new_n920));
  INV_X1    g719(.A(new_n859), .ZN(new_n921));
  INV_X1    g720(.A(new_n885), .ZN(new_n922));
  NAND4_X1  g721(.A1(new_n882), .A2(new_n695), .A3(new_n723), .A4(new_n883), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n876), .A2(KEYINPUT119), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n871), .A2(new_n873), .A3(new_n875), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n696), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g727(.A(new_n922), .B1(new_n928), .B2(new_n669), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n921), .B1(new_n929), .B2(new_n583), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(new_n498), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n920), .B1(new_n931), .B2(KEYINPUT57), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n746), .A2(new_n892), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(KEYINPUT123), .B1(new_n934), .B2(new_n896), .ZN(new_n935));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n936));
  NAND4_X1  g735(.A1(new_n932), .A2(new_n936), .A3(new_n696), .A4(new_n933), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n935), .A2(G141gat), .A3(new_n937), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT58), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n919), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT120), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n932), .A2(new_n941), .A3(new_n933), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n932), .B2(new_n933), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n696), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n918), .B1(new_n945), .B2(G141gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n940), .B1(new_n946), .B2(new_n939), .ZN(G1344gat));
  INV_X1    g746(.A(KEYINPUT57), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n930), .A2(new_n948), .A3(new_n498), .ZN(new_n949));
  OAI21_X1  g748(.A(KEYINPUT57), .B1(new_n890), .B2(new_n493), .ZN(new_n950));
  AND2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(new_n723), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(KEYINPUT59), .A3(new_n933), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n934), .A2(KEYINPUT120), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n724), .B1(new_n954), .B2(new_n942), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n953), .B1(new_n955), .B2(KEYINPUT59), .ZN(new_n956));
  AND3_X1   g755(.A1(new_n914), .A2(new_n893), .A3(new_n916), .ZN(new_n957));
  AOI21_X1  g756(.A(G148gat), .B1(new_n957), .B2(new_n723), .ZN(new_n958));
  AOI22_X1  g757(.A1(new_n956), .A2(G148gat), .B1(KEYINPUT59), .B2(new_n958), .ZN(G1345gat));
  AOI21_X1  g758(.A(G155gat), .B1(new_n957), .B2(new_n583), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n943), .A2(new_n944), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n961), .A2(new_n889), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n960), .B1(new_n962), .B2(G155gat), .ZN(G1346gat));
  AOI21_X1  g762(.A(new_n368), .B1(new_n957), .B2(new_n755), .ZN(new_n964));
  NOR2_X1   g763(.A1(new_n961), .A2(new_n669), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n964), .B1(new_n965), .B2(new_n368), .ZN(G1347gat));
  NOR2_X1   g765(.A1(new_n890), .A2(new_n804), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n503), .A2(new_n506), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G169gat), .B1(new_n970), .B2(new_n896), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT124), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n972), .B1(new_n890), .B2(new_n804), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n923), .B1(new_n896), .B2(new_n925), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n669), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n583), .B1(new_n975), .B2(new_n885), .ZN(new_n976));
  OAI211_X1 g775(.A(KEYINPUT124), .B(new_n445), .C1(new_n976), .C2(new_n859), .ZN(new_n977));
  AND3_X1   g776(.A1(new_n973), .A2(new_n968), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n978), .A2(new_n207), .A3(new_n696), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n971), .A2(new_n979), .ZN(G1348gat));
  NOR3_X1   g779(.A1(new_n970), .A2(new_n208), .A3(new_n724), .ZN(new_n981));
  AOI21_X1  g780(.A(G176gat), .B1(new_n978), .B2(new_n723), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n981), .A2(new_n982), .ZN(G1349gat));
  OAI21_X1  g782(.A(G183gat), .B1(new_n970), .B2(new_n889), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n978), .A2(new_n246), .A3(new_n583), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n986), .B(KEYINPUT60), .ZN(G1350gat));
  AOI21_X1  g786(.A(new_n215), .B1(new_n969), .B2(new_n755), .ZN(new_n988));
  XOR2_X1   g787(.A(new_n988), .B(KEYINPUT61), .Z(new_n989));
  NAND3_X1  g788(.A1(new_n978), .A2(new_n215), .A3(new_n755), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n989), .A2(new_n990), .ZN(G1351gat));
  NOR3_X1   g790(.A1(new_n746), .A2(new_n804), .A3(new_n506), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n951), .A2(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(G197gat), .B1(new_n993), .B2(new_n896), .ZN(new_n994));
  AOI211_X1 g793(.A(new_n493), .B(new_n506), .C1(new_n740), .C2(new_n744), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n973), .A2(new_n995), .A3(new_n977), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n997));
  INV_X1    g796(.A(G197gat), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT125), .ZN(new_n999));
  NAND4_X1  g798(.A1(new_n973), .A2(new_n995), .A3(new_n999), .A4(new_n977), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n997), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n994), .B1(new_n896), .B2(new_n1001), .ZN(G1352gat));
  OR3_X1    g801(.A1(new_n996), .A2(G204gat), .A3(new_n724), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  OR2_X1    g803(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1005));
  AND2_X1   g804(.A1(new_n952), .A2(new_n992), .ZN(new_n1006));
  OAI211_X1 g805(.A(new_n1004), .B(new_n1005), .C1(new_n1006), .C2(new_n718), .ZN(G1353gat));
  NAND4_X1  g806(.A1(new_n997), .A2(new_n316), .A3(new_n583), .A4(new_n1000), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n951), .A2(new_n583), .A3(new_n992), .ZN(new_n1009));
  AND3_X1   g808(.A1(new_n1009), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(KEYINPUT63), .B1(new_n1009), .B2(G211gat), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1008), .B1(new_n1010), .B2(new_n1011), .ZN(G1354gat));
  NAND4_X1  g811(.A1(new_n951), .A2(new_n318), .A3(new_n755), .A4(new_n992), .ZN(new_n1013));
  NAND3_X1  g812(.A1(new_n997), .A2(new_n755), .A3(new_n1000), .ZN(new_n1014));
  AND3_X1   g813(.A1(new_n1014), .A2(KEYINPUT126), .A3(new_n315), .ZN(new_n1015));
  AOI21_X1  g814(.A(KEYINPUT126), .B1(new_n1014), .B2(new_n315), .ZN(new_n1016));
  OAI21_X1  g815(.A(new_n1013), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1017), .A2(KEYINPUT127), .ZN(new_n1018));
  INV_X1    g817(.A(KEYINPUT127), .ZN(new_n1019));
  OAI211_X1 g818(.A(new_n1019), .B(new_n1013), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1020));
  NAND2_X1  g819(.A1(new_n1018), .A2(new_n1020), .ZN(G1355gat));
endmodule


