//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 1 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 0 0 1 1 1 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n766, new_n767, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT83), .Z(new_n189));
  INV_X1    g003(.A(KEYINPUT12), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT11), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G137), .ZN(new_n193));
  AOI21_X1  g007(.A(G131), .B1(new_n192), .B2(G137), .ZN(new_n194));
  INV_X1    g008(.A(G137), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n195), .A2(KEYINPUT11), .A3(G134), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n193), .A2(new_n194), .A3(KEYINPUT65), .A4(new_n196), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(new_n196), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n195), .A2(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(G131), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT69), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n201), .A2(KEYINPUT69), .A3(new_n204), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G128), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n211), .B(new_n213), .C1(KEYINPUT1), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G104), .ZN(new_n220));
  OAI21_X1  g034(.A(KEYINPUT3), .B1(new_n220), .B2(G107), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n222));
  INV_X1    g036(.A(G107), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n222), .A2(new_n223), .A3(G104), .ZN(new_n224));
  INV_X1    g038(.A(G101), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n220), .A2(G107), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n221), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n220), .A2(G107), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n223), .A2(G104), .ZN(new_n229));
  OAI21_X1  g043(.A(G101), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n216), .A2(new_n218), .A3(new_n227), .A4(new_n230), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n190), .B1(new_n209), .B2(new_n234), .ZN(new_n235));
  AND2_X1   g049(.A1(new_n201), .A2(new_n204), .ZN(new_n236));
  OR3_X1    g050(.A1(new_n234), .A2(new_n190), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G110), .B(G140), .ZN(new_n239));
  INV_X1    g053(.A(G953), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G227), .ZN(new_n241));
  XOR2_X1   g055(.A(new_n239), .B(new_n241), .Z(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n221), .A2(new_n224), .A3(new_n226), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n246));
  OAI21_X1  g060(.A(KEYINPUT84), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n244), .A2(G101), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT84), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n249), .A3(KEYINPUT4), .A4(new_n227), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  OAI21_X1  g066(.A(KEYINPUT64), .B1(new_n214), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n252), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT64), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n254), .A2(new_n211), .A3(new_n213), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  OR2_X1    g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n214), .A2(new_n252), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n244), .A2(new_n260), .A3(G101), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n257), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n233), .A2(KEYINPUT10), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n216), .A2(new_n218), .ZN(new_n264));
  INV_X1    g078(.A(new_n231), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT10), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n264), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI22_X1  g081(.A1(new_n251), .A2(new_n262), .B1(new_n263), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT85), .ZN(new_n269));
  AND3_X1   g083(.A1(new_n268), .A2(new_n269), .A3(new_n209), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n269), .B1(new_n268), .B2(new_n209), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n238), .B(new_n243), .C1(new_n270), .C2(new_n271), .ZN(new_n272));
  NOR2_X1   g086(.A1(new_n268), .A2(new_n209), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n251), .A2(new_n262), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n267), .A2(new_n263), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n209), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT85), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n269), .A3(new_n209), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n273), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n272), .B1(new_n279), .B2(new_n243), .ZN(new_n280));
  INV_X1    g094(.A(G469), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT87), .ZN(new_n284));
  INV_X1    g098(.A(new_n273), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n270), .B2(new_n271), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n242), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n287), .B2(new_n272), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT87), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n288), .A2(new_n289), .A3(new_n281), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n277), .A2(new_n278), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(new_n238), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n242), .ZN(new_n294));
  OAI211_X1 g108(.A(KEYINPUT86), .B(new_n243), .C1(new_n270), .C2(new_n271), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n285), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT86), .B1(new_n292), .B2(new_n243), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n294), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(new_n282), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G469), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n189), .B1(new_n291), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(G210), .B1(G237), .B2(G902), .ZN(new_n303));
  XNOR2_X1  g117(.A(G110), .B(G122), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT2), .ZN(new_n306));
  INV_X1    g120(.A(G113), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT66), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(KEYINPUT2), .A3(G113), .ZN(new_n310));
  AOI22_X1  g124(.A1(new_n308), .A2(new_n310), .B1(new_n306), .B2(new_n307), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G116), .ZN(new_n313));
  OAI21_X1  g127(.A(KEYINPUT67), .B1(new_n313), .B2(G119), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT67), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G116), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(G119), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(KEYINPUT68), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT68), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n314), .A2(new_n317), .A3(new_n321), .A4(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n312), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n311), .A2(new_n314), .A3(new_n317), .A4(new_n318), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n323), .A2(new_n324), .B1(new_n260), .B2(new_n245), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n325), .A2(new_n251), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n316), .A2(G116), .ZN(new_n327));
  OAI21_X1  g141(.A(G113), .B1(new_n327), .B2(KEYINPUT5), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n320), .A2(new_n322), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(KEYINPUT5), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n312), .A2(new_n319), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n330), .A2(new_n331), .A3(new_n231), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n305), .B1(new_n326), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n329), .A2(KEYINPUT5), .ZN(new_n334));
  INV_X1    g148(.A(new_n328), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n331), .A2(new_n231), .ZN(new_n337));
  AOI22_X1  g151(.A1(new_n251), .A2(new_n325), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n304), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n333), .A2(new_n339), .A3(KEYINPUT6), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n338), .A2(KEYINPUT6), .A3(new_n304), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n264), .A2(G125), .ZN(new_n342));
  INV_X1    g156(.A(G125), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n343), .B1(new_n257), .B2(new_n259), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n342), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G224), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(G953), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n345), .B(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n340), .A2(new_n341), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n231), .B1(new_n330), .B2(new_n331), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n314), .A2(new_n317), .A3(KEYINPUT5), .A4(new_n318), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n328), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n354), .B1(new_n353), .B2(new_n352), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n337), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n304), .B(KEYINPUT8), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n304), .A2(new_n338), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT7), .ZN(new_n360));
  OAI22_X1  g174(.A1(new_n342), .A2(new_n344), .B1(new_n360), .B2(new_n347), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT89), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n348), .ZN(new_n364));
  OAI221_X1 g178(.A(KEYINPUT89), .B1(new_n360), .B2(new_n347), .C1(new_n342), .C2(new_n344), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n350), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT90), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n303), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n350), .A2(new_n367), .A3(KEYINPUT90), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n350), .A2(new_n367), .A3(new_n303), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT91), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G214), .B1(G237), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT91), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n370), .A2(new_n378), .A3(new_n371), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(G140), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G125), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n343), .A2(G140), .ZN(new_n383));
  AND2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(new_n210), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT79), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n387), .B1(new_n386), .B2(new_n382), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n385), .B1(new_n388), .B2(new_n210), .ZN(new_n389));
  OR2_X1    g203(.A1(KEYINPUT71), .A2(G237), .ZN(new_n390));
  NAND2_X1  g204(.A1(KEYINPUT71), .A2(G237), .ZN(new_n391));
  AOI21_X1  g205(.A(G953), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G143), .A3(G214), .ZN(new_n393));
  AND2_X1   g207(.A1(KEYINPUT71), .A2(G237), .ZN(new_n394));
  NOR2_X1   g208(.A1(KEYINPUT71), .A2(G237), .ZN(new_n395));
  OAI211_X1 g209(.A(G214), .B(new_n240), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n212), .ZN(new_n397));
  NAND2_X1  g211(.A1(KEYINPUT18), .A2(G131), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n393), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n389), .A2(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n398), .B1(new_n393), .B2(new_n397), .ZN(new_n401));
  OAI21_X1  g215(.A(KEYINPUT92), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT92), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n403), .A2(new_n404), .A3(new_n389), .A4(new_n399), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n393), .A2(new_n397), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(G131), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT17), .ZN(new_n409));
  INV_X1    g223(.A(G131), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n393), .A2(new_n397), .A3(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n408), .A2(KEYINPUT93), .A3(new_n409), .A4(new_n411), .ZN(new_n412));
  OAI211_X1 g226(.A(new_n387), .B(KEYINPUT16), .C1(new_n386), .C2(new_n382), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT16), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n382), .A2(new_n414), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n413), .A2(new_n210), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n210), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n410), .B1(new_n393), .B2(new_n397), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(KEYINPUT17), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n412), .A2(new_n418), .A3(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n393), .A2(new_n410), .A3(new_n397), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(new_n419), .ZN(new_n423));
  AOI21_X1  g237(.A(KEYINPUT93), .B1(new_n423), .B2(new_n409), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n406), .B1(new_n421), .B2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(G113), .B(G122), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n426), .B(new_n220), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n425), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n406), .B(new_n427), .C1(new_n421), .C2(new_n424), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(G475), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n413), .A2(new_n415), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G146), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n384), .A2(KEYINPUT19), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n388), .B2(KEYINPUT19), .ZN(new_n437));
  OAI221_X1 g251(.A(new_n435), .B1(new_n437), .B2(G146), .C1(new_n419), .C2(new_n422), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n406), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(new_n428), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(new_n430), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT94), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n444), .B1(new_n440), .B2(new_n430), .ZN(new_n445));
  OAI21_X1  g259(.A(new_n443), .B1(KEYINPUT20), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT20), .ZN(new_n447));
  NAND4_X1  g261(.A1(new_n441), .A2(new_n444), .A3(new_n447), .A4(new_n442), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n433), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(G234), .A2(G237), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n450), .A2(G952), .A3(new_n240), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n450), .A2(G902), .A3(G953), .ZN(new_n452));
  XNOR2_X1  g266(.A(KEYINPUT21), .B(G898), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n313), .A2(KEYINPUT14), .A3(G122), .ZN(new_n456));
  XOR2_X1   g270(.A(G116), .B(G122), .Z(new_n457));
  OAI211_X1 g271(.A(G107), .B(new_n456), .C1(new_n457), .C2(KEYINPUT14), .ZN(new_n458));
  XNOR2_X1  g272(.A(G116), .B(G122), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n223), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n212), .A2(G128), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n217), .A2(G143), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n192), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n192), .B1(new_n461), .B2(new_n462), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n458), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT96), .ZN(new_n467));
  XOR2_X1   g281(.A(KEYINPUT95), .B(KEYINPUT13), .Z(new_n468));
  INV_X1    g282(.A(new_n461), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n467), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT95), .B(KEYINPUT13), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(KEYINPUT96), .A3(new_n461), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n462), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n474), .B1(new_n468), .B2(new_n469), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n192), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n457), .A2(G107), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n477), .A2(new_n460), .B1(KEYINPUT97), .B2(new_n463), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n478), .B1(KEYINPUT97), .B2(new_n463), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n466), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(G217), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n187), .A2(new_n481), .A3(G953), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  OAI211_X1 g298(.A(new_n466), .B(new_n482), .C1(new_n476), .C2(new_n479), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n282), .ZN(new_n487));
  INV_X1    g301(.A(G478), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n488), .A2(KEYINPUT15), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G902), .B1(new_n484), .B2(new_n485), .ZN(new_n491));
  INV_X1    g305(.A(new_n489), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n490), .A2(KEYINPUT98), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT98), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n491), .A2(new_n492), .ZN(new_n496));
  AOI211_X1 g310(.A(G902), .B(new_n489), .C1(new_n484), .C2(new_n485), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n449), .A2(new_n455), .A3(new_n499), .ZN(new_n500));
  NOR3_X1   g314(.A1(new_n302), .A2(new_n380), .A3(new_n500), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT22), .B(G137), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n240), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n502), .B(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT76), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n505), .B1(new_n217), .B2(G119), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n316), .A2(KEYINPUT76), .A3(G128), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n507), .C1(new_n316), .C2(G128), .ZN(new_n508));
  XNOR2_X1  g322(.A(KEYINPUT24), .B(G110), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n508), .A2(KEYINPUT80), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n316), .A2(G128), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n217), .A2(KEYINPUT23), .A3(G119), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n316), .A2(G128), .ZN(new_n513));
  OAI211_X1 g327(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(KEYINPUT23), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n510), .B1(G110), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT80), .B1(new_n508), .B2(new_n509), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n435), .B(new_n385), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n514), .A2(G110), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT78), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT78), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n514), .A2(new_n520), .A3(G110), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n507), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n523), .A2(new_n513), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT77), .ZN(new_n525));
  INV_X1    g339(.A(new_n509), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n524), .A2(new_n525), .A3(new_n526), .A4(new_n506), .ZN(new_n527));
  OAI21_X1  g341(.A(KEYINPUT77), .B1(new_n508), .B2(new_n509), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n522), .B(new_n529), .C1(new_n416), .C2(new_n417), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT81), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n517), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n531), .B1(new_n517), .B2(new_n530), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n504), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n504), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n517), .A2(new_n530), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n535), .B1(new_n536), .B2(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n282), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT25), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n534), .A2(KEYINPUT25), .A3(new_n282), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n481), .B1(G234), .B2(new_n282), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n543), .A2(G902), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n537), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n257), .A2(new_n259), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n207), .A2(new_n208), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(KEYINPUT70), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT70), .ZN(new_n552));
  NAND4_X1  g366(.A1(new_n207), .A2(new_n552), .A3(new_n208), .A4(new_n549), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n192), .A2(G137), .ZN(new_n554));
  OAI21_X1  g368(.A(G131), .B1(new_n554), .B2(new_n203), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n264), .A2(new_n201), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n551), .A2(KEYINPUT30), .A3(new_n553), .A4(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n236), .B2(new_n548), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT30), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n323), .A2(new_n324), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n557), .A2(new_n562), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n556), .A2(new_n323), .A3(new_n324), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n551), .A2(new_n553), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n392), .A2(G210), .ZN(new_n566));
  XNOR2_X1  g380(.A(new_n566), .B(KEYINPUT27), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT26), .B(G101), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n567), .B(new_n568), .ZN(new_n569));
  AND3_X1   g383(.A1(new_n565), .A2(KEYINPUT72), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(KEYINPUT72), .B1(new_n565), .B2(new_n569), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n563), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT73), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT73), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n574), .B(new_n563), .C1(new_n570), .C2(new_n571), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n573), .A2(KEYINPUT31), .A3(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT31), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n577), .B(new_n563), .C1(new_n570), .C2(new_n571), .ZN(new_n578));
  INV_X1    g392(.A(new_n569), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n550), .A2(new_n556), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n561), .B1(new_n580), .B2(KEYINPUT74), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT74), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n550), .A2(new_n582), .A3(new_n556), .ZN(new_n583));
  AOI21_X1  g397(.A(KEYINPUT28), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT28), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n558), .A2(new_n561), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n585), .B1(new_n565), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n579), .B1(new_n584), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g402(.A1(new_n578), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n576), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(G472), .A2(G902), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT32), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(new_n591), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(new_n593), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n581), .A2(new_n583), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n585), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n569), .A2(KEYINPUT29), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n551), .A2(new_n553), .A3(new_n556), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n561), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(new_n565), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT75), .B1(new_n602), .B2(KEYINPUT28), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT75), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n604), .B(new_n585), .C1(new_n601), .C2(new_n565), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n598), .B(new_n599), .C1(new_n603), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n563), .A2(new_n565), .ZN(new_n607));
  AOI21_X1  g421(.A(KEYINPUT29), .B1(new_n607), .B2(new_n579), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n565), .A2(new_n586), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT28), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n598), .A2(new_n569), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(G902), .B1(new_n608), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n590), .A2(new_n596), .B1(new_n613), .B2(G472), .ZN(new_n614));
  AOI211_X1 g428(.A(KEYINPUT82), .B(new_n547), .C1(new_n594), .C2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT82), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n590), .A2(new_n596), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n613), .A2(G472), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n595), .B1(new_n576), .B2(new_n589), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n617), .B(new_n618), .C1(KEYINPUT32), .C2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(new_n547), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n501), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(KEYINPUT99), .B(G101), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT100), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n623), .B(new_n625), .ZN(G3));
  NAND2_X1  g440(.A1(new_n590), .A2(new_n282), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(KEYINPUT101), .A3(G472), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n628), .A2(new_n592), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(G472), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n633), .A2(new_n547), .A3(new_n302), .ZN(new_n634));
  INV_X1    g448(.A(new_n377), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n303), .B1(new_n350), .B2(new_n367), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n635), .B1(new_n637), .B2(new_n373), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n455), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT33), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n486), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(G478), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n488), .A2(new_n282), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n643), .B1(new_n491), .B2(new_n488), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n639), .A2(new_n449), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n634), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT102), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT34), .B(G104), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G6));
  AOI21_X1  g464(.A(new_n447), .B1(new_n441), .B2(new_n442), .ZN(new_n651));
  INV_X1    g465(.A(new_n442), .ZN(new_n652));
  AOI211_X1 g466(.A(KEYINPUT20), .B(new_n652), .C1(new_n440), .C2(new_n430), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR4_X1   g468(.A1(new_n639), .A2(new_n433), .A3(new_n499), .A4(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n634), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G107), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G9));
  INV_X1    g473(.A(new_n545), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT104), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n536), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n536), .B(KEYINPUT104), .ZN(new_n665));
  INV_X1    g479(.A(new_n663), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n660), .B1(new_n664), .B2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n668), .B1(new_n542), .B2(new_n543), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n500), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n670), .A2(new_n380), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n629), .A2(new_n301), .A3(new_n632), .A4(new_n671), .ZN(new_n672));
  XOR2_X1   g486(.A(KEYINPUT37), .B(G110), .Z(new_n673));
  XNOR2_X1  g487(.A(new_n672), .B(new_n673), .ZN(G12));
  AOI21_X1  g488(.A(new_n289), .B1(new_n288), .B2(new_n281), .ZN(new_n675));
  AND4_X1   g489(.A1(new_n289), .A2(new_n280), .A3(new_n281), .A4(new_n282), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n243), .B1(new_n270), .B2(new_n271), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT86), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n285), .A3(new_n295), .ZN(new_n680));
  AOI21_X1  g494(.A(G902), .B1(new_n680), .B2(new_n294), .ZN(new_n681));
  OAI22_X1  g495(.A1(new_n675), .A2(new_n676), .B1(new_n681), .B2(new_n281), .ZN(new_n682));
  INV_X1    g496(.A(new_n373), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n377), .B1(new_n683), .B2(new_n636), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n669), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n452), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n451), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NOR4_X1   g504(.A1(new_n499), .A2(new_n654), .A3(new_n433), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n189), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n682), .A2(new_n685), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n620), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  INV_X1    g510(.A(KEYINPUT106), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n602), .A2(new_n579), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n573), .A2(new_n575), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n282), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n700), .A2(G472), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n617), .A2(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n619), .A2(KEYINPUT32), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n702), .A2(new_n703), .A3(KEYINPUT105), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT105), .ZN(new_n705));
  INV_X1    g519(.A(new_n596), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n576), .B2(new_n589), .ZN(new_n707));
  INV_X1    g521(.A(G472), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n708), .B1(new_n699), .B2(new_n282), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n705), .B1(new_n594), .B2(new_n710), .ZN(new_n711));
  OAI21_X1  g525(.A(new_n697), .B1(new_n704), .B2(new_n711), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT105), .B1(new_n702), .B2(new_n703), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n594), .A2(new_n710), .A3(new_n705), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n713), .A2(KEYINPUT106), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n376), .A2(new_n379), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(KEYINPUT38), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(new_n449), .ZN(new_n720));
  INV_X1    g534(.A(new_n499), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n669), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n722), .A2(new_n635), .A3(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n689), .B(KEYINPUT39), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n301), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n726), .B(KEYINPUT40), .Z(new_n727));
  NAND4_X1  g541(.A1(new_n716), .A2(new_n719), .A3(new_n724), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G143), .ZN(G45));
  NOR3_X1   g543(.A1(new_n449), .A2(new_n645), .A3(new_n690), .ZN(new_n730));
  AND4_X1   g544(.A1(new_n692), .A2(new_n682), .A3(new_n730), .A4(new_n685), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n620), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G146), .ZN(G48));
  NAND2_X1  g547(.A1(new_n620), .A2(new_n621), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n735));
  OR2_X1    g549(.A1(new_n288), .A2(new_n281), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n291), .A2(new_n735), .A3(new_n692), .A4(new_n736), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n736), .B(new_n692), .C1(new_n675), .C2(new_n676), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT107), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n646), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n734), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g555(.A(KEYINPUT41), .B(G113), .Z(new_n742));
  XNOR2_X1  g556(.A(new_n741), .B(new_n742), .ZN(G15));
  NAND3_X1  g557(.A1(new_n655), .A2(new_n737), .A3(new_n739), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n734), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n313), .ZN(G18));
  NAND3_X1  g560(.A1(new_n739), .A2(new_n638), .A3(new_n737), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n670), .B1(new_n594), .B2(new_n614), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G119), .ZN(G21));
  NAND2_X1  g565(.A1(new_n576), .A2(new_n578), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n602), .A2(KEYINPUT28), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n604), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n602), .A2(KEYINPUT75), .A3(KEYINPUT28), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n569), .B1(new_n756), .B2(new_n598), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n591), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n630), .A2(new_n621), .A3(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n722), .A2(new_n639), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n739), .A3(new_n737), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n760), .A2(new_n763), .ZN(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(G122), .ZN(G24));
  NAND4_X1  g579(.A1(new_n630), .A2(new_n723), .A3(new_n758), .A4(new_n730), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n766), .A2(new_n747), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n343), .ZN(G27));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n290), .A2(new_n284), .B1(new_n299), .B2(G469), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(new_n189), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n682), .A2(KEYINPUT108), .A3(new_n692), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n635), .B1(new_n376), .B2(new_n379), .ZN(new_n773));
  AND3_X1   g587(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n547), .B1(new_n594), .B2(new_n614), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT109), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(KEYINPUT42), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n774), .A2(new_n775), .A3(new_n730), .A4(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n780));
  INV_X1    g594(.A(new_n730), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n734), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT109), .B(KEYINPUT42), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G131), .ZN(G33));
  NAND3_X1  g599(.A1(new_n774), .A2(new_n775), .A3(new_n691), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  INV_X1    g601(.A(new_n645), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n449), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT43), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT43), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n449), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n632), .A2(new_n592), .A3(new_n628), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n794), .A2(KEYINPUT111), .A3(new_n669), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT111), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n633), .B2(new_n723), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n793), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n281), .A2(new_n282), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n298), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n680), .A2(KEYINPUT45), .A3(new_n294), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(G469), .A3(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n803), .A2(new_n804), .A3(KEYINPUT110), .A4(G469), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n801), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n809), .A2(KEYINPUT46), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n291), .B1(new_n809), .B2(KEYINPUT46), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n812), .A2(new_n189), .ZN(new_n813));
  AND3_X1   g627(.A1(new_n813), .A2(new_n725), .A3(new_n773), .ZN(new_n814));
  OAI211_X1 g628(.A(KEYINPUT44), .B(new_n793), .C1(new_n795), .C2(new_n797), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n800), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G137), .ZN(G39));
  NAND3_X1  g631(.A1(new_n773), .A2(new_n547), .A3(new_n730), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT47), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n812), .B2(new_n189), .ZN(new_n820));
  OAI211_X1 g634(.A(KEYINPUT47), .B(new_n692), .C1(new_n810), .C2(new_n811), .ZN(new_n821));
  AOI211_X1 g635(.A(new_n620), .B(new_n818), .C1(new_n820), .C2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(new_n381), .ZN(G42));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n734), .B1(new_n740), .B2(new_n744), .ZN(new_n825));
  INV_X1    g639(.A(new_n670), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n620), .A2(new_n826), .ZN(new_n827));
  OAI22_X1  g641(.A1(new_n827), .A2(new_n747), .B1(new_n759), .B2(new_n762), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n496), .A2(new_n497), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n720), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n449), .A2(new_n645), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n833), .A2(new_n380), .A3(new_n454), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n794), .A2(new_n621), .A3(new_n301), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n829), .A2(new_n623), .A3(new_n672), .A4(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n630), .A2(new_n723), .A3(new_n730), .A4(new_n758), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n774), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n302), .A2(new_n690), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n654), .A2(new_n433), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n723), .A2(new_n830), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g655(.A1(new_n839), .A2(new_n620), .A3(new_n773), .A4(new_n841), .ZN(new_n842));
  AND3_X1   g656(.A1(new_n786), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n784), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n836), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n693), .B1(new_n594), .B2(new_n614), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n846), .B1(new_n837), .B2(new_n748), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n720), .A2(new_n638), .A3(new_n721), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n723), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n849), .A2(new_n301), .A3(new_n689), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n704), .B2(new_n711), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT52), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n847), .A2(new_n852), .A3(new_n853), .A4(new_n732), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n695), .B(new_n732), .C1(new_n766), .C2(new_n747), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n850), .B1(new_n713), .B2(new_n714), .ZN(new_n856));
  OAI21_X1  g670(.A(KEYINPUT52), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n847), .A2(new_n853), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n845), .B(new_n858), .C1(KEYINPUT53), .C2(new_n859), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n760), .A2(new_n763), .B1(new_n748), .B2(new_n749), .ZN(new_n861));
  AND2_X1   g675(.A1(new_n739), .A2(new_n737), .ZN(new_n862));
  OAI211_X1 g676(.A(new_n775), .B(new_n862), .C1(new_n646), .C2(new_n655), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n623), .A2(new_n861), .A3(new_n672), .A4(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n835), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n786), .A2(new_n838), .A3(new_n842), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n774), .A2(new_n775), .A3(new_n730), .ZN(new_n868));
  INV_X1    g682(.A(new_n783), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n870), .B2(new_n779), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n866), .A2(new_n858), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT53), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n824), .B1(new_n860), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n790), .A2(new_n451), .A3(new_n792), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT113), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n877), .B(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n879), .A2(new_n759), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n718), .A2(new_n635), .A3(new_n862), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT114), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT50), .ZN(new_n884));
  NAND4_X1  g698(.A1(new_n880), .A2(new_n882), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  NAND2_X1  g700(.A1(KEYINPUT114), .A2(KEYINPUT50), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n877), .B(KEYINPUT113), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(new_n760), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n886), .B(new_n887), .C1(new_n889), .C2(new_n881), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n885), .A2(new_n890), .A3(KEYINPUT115), .ZN(new_n891));
  AOI21_X1  g705(.A(KEYINPUT115), .B1(new_n885), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n862), .A2(new_n773), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n894), .A2(new_n547), .A3(new_n688), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n720), .A2(new_n788), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n895), .A2(new_n715), .A3(new_n712), .A4(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n879), .A2(new_n894), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n898), .A2(new_n630), .A3(new_n723), .A4(new_n758), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n291), .A2(new_n736), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT112), .Z(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n189), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n820), .A2(new_n821), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n717), .A2(new_n377), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n889), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n900), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  AOI21_X1  g721(.A(KEYINPUT51), .B1(new_n893), .B2(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n879), .A2(new_n894), .A3(new_n734), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT48), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n832), .A2(new_n895), .A3(new_n715), .A4(new_n712), .ZN(new_n911));
  OAI211_X1 g725(.A(G952), .B(new_n240), .C1(new_n889), .C2(new_n747), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n904), .A2(new_n906), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(new_n899), .A3(new_n897), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n885), .A2(new_n890), .A3(KEYINPUT51), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n908), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n859), .A2(new_n873), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n866), .A2(new_n858), .A3(new_n871), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n854), .A2(new_n857), .ZN(new_n921));
  NOR3_X1   g735(.A1(new_n836), .A2(new_n921), .A3(new_n844), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n824), .B(new_n920), .C1(new_n922), .C2(KEYINPUT53), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n876), .A2(new_n918), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(KEYINPUT116), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT116), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n876), .A2(new_n918), .A3(new_n926), .A4(new_n923), .ZN(new_n927));
  INV_X1    g741(.A(G952), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n928), .A2(new_n240), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n925), .A2(new_n927), .A3(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n902), .B(KEYINPUT49), .Z(new_n931));
  OR4_X1    g745(.A1(new_n547), .A2(new_n789), .A3(new_n635), .A4(new_n189), .ZN(new_n932));
  OR4_X1    g746(.A1(new_n716), .A2(new_n931), .A3(new_n719), .A4(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n933), .ZN(G75));
  NOR2_X1   g748(.A1(new_n240), .A2(G952), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n845), .B2(new_n858), .ZN(new_n937));
  AND4_X1   g751(.A1(new_n866), .A2(new_n858), .A3(new_n871), .A4(new_n919), .ZN(new_n938));
  OAI21_X1  g752(.A(G902), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(KEYINPUT56), .B1(new_n940), .B2(G210), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n340), .A2(new_n341), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(new_n349), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT55), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n936), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n939), .A2(KEYINPUT117), .ZN(new_n946));
  INV_X1    g760(.A(new_n303), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT117), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n948), .B(G902), .C1(new_n937), .C2(new_n938), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n946), .A2(KEYINPUT118), .A3(new_n947), .A4(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT56), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n944), .A2(new_n951), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n946), .A2(new_n947), .A3(new_n949), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT118), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n945), .B1(new_n953), .B2(new_n956), .ZN(G51));
  XNOR2_X1  g771(.A(new_n801), .B(KEYINPUT57), .ZN(new_n958));
  INV_X1    g772(.A(new_n923), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n824), .B1(new_n874), .B2(new_n920), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT119), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  OAI211_X1 g777(.A(KEYINPUT119), .B(new_n958), .C1(new_n959), .C2(new_n960), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n280), .A3(new_n964), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n946), .A2(new_n807), .A3(new_n808), .A4(new_n949), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n935), .B1(new_n965), .B2(new_n966), .ZN(G54));
  NAND2_X1  g781(.A1(KEYINPUT58), .A2(G475), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT120), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n946), .A2(new_n949), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n430), .A3(new_n440), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n946), .A2(new_n441), .A3(new_n949), .A4(new_n969), .ZN(new_n972));
  AND3_X1   g786(.A1(new_n971), .A2(new_n936), .A3(new_n972), .ZN(G60));
  INV_X1    g787(.A(KEYINPUT121), .ZN(new_n974));
  INV_X1    g788(.A(new_n641), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n643), .B(KEYINPUT59), .Z(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  INV_X1    g791(.A(new_n960), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n977), .B1(new_n978), .B2(new_n923), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n974), .B1(new_n979), .B2(new_n935), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n959), .A2(new_n960), .ZN(new_n981));
  OAI211_X1 g795(.A(KEYINPUT121), .B(new_n936), .C1(new_n981), .C2(new_n977), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n959), .B2(new_n875), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n641), .ZN(new_n984));
  AND3_X1   g798(.A1(new_n980), .A2(new_n982), .A3(new_n984), .ZN(G63));
  NAND2_X1  g799(.A1(new_n874), .A2(new_n920), .ZN(new_n986));
  NAND2_X1  g800(.A1(G217), .A2(G902), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT122), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT60), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n986), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n534), .A2(new_n537), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n664), .A2(new_n667), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n986), .A2(new_n993), .A3(new_n989), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n936), .A3(new_n994), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT61), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n995), .B(new_n996), .ZN(G66));
  OAI21_X1  g811(.A(G953), .B1(new_n453), .B2(new_n346), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT123), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n866), .B2(G953), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n942), .B1(G898), .B2(new_n240), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(G69));
  NOR2_X1   g816(.A1(new_n615), .A2(new_n622), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n833), .B(KEYINPUT124), .Z(new_n1004));
  NOR4_X1   g818(.A1(new_n1003), .A2(new_n1004), .A3(new_n726), .A4(new_n905), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n822), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(new_n855), .ZN(new_n1007));
  AOI21_X1  g821(.A(KEYINPUT62), .B1(new_n728), .B2(new_n1007), .ZN(new_n1008));
  AND3_X1   g822(.A1(new_n728), .A2(KEYINPUT62), .A3(new_n1007), .ZN(new_n1009));
  OAI211_X1 g823(.A(new_n1006), .B(new_n816), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n240), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n557), .A2(new_n560), .ZN(new_n1012));
  XOR2_X1   g826(.A(new_n1012), .B(new_n437), .Z(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1013), .B1(G900), .B2(G953), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n784), .A2(new_n786), .A3(new_n1007), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n822), .A2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n734), .A2(new_n848), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n813), .A2(new_n725), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g833(.A(new_n1019), .B(KEYINPUT126), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n1017), .A2(new_n1020), .A3(new_n816), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1015), .B1(new_n1021), .B2(G953), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1014), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n240), .B1(G227), .B2(G900), .ZN(new_n1024));
  INV_X1    g838(.A(KEYINPUT125), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1026));
  AND2_X1   g840(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1023), .A2(new_n1026), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n1027), .A2(new_n1028), .ZN(G72));
  NAND4_X1  g843(.A1(new_n1020), .A2(new_n1017), .A3(new_n816), .A4(new_n866), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  NAND2_X1  g846(.A1(new_n1030), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT127), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1030), .A2(KEYINPUT127), .A3(new_n1032), .ZN(new_n1036));
  AOI211_X1 g850(.A(new_n569), .B(new_n607), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1032), .B1(new_n1010), .B2(new_n836), .ZN(new_n1038));
  NAND3_X1  g852(.A1(new_n1038), .A2(new_n569), .A3(new_n607), .ZN(new_n1039));
  NAND2_X1  g853(.A1(new_n860), .A2(new_n874), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n573), .A2(new_n575), .ZN(new_n1041));
  AOI21_X1  g855(.A(new_n569), .B1(new_n563), .B2(new_n565), .ZN(new_n1042));
  OAI211_X1 g856(.A(new_n1040), .B(new_n1032), .C1(new_n1041), .C2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n1039), .A2(new_n936), .A3(new_n1043), .ZN(new_n1044));
  NOR2_X1   g858(.A1(new_n1037), .A2(new_n1044), .ZN(G57));
endmodule


