//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n763, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n807, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n190), .B1(new_n191), .B2(G146), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n188), .A2(KEYINPUT64), .A3(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n192), .B2(new_n193), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G146), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n189), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n194), .A2(new_n197), .B1(new_n200), .B2(new_n195), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT11), .ZN(new_n202));
  INV_X1    g016(.A(G134), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n202), .B1(new_n203), .B2(G137), .ZN(new_n204));
  INV_X1    g018(.A(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(KEYINPUT11), .A3(G134), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n203), .A2(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n206), .A3(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n204), .A2(new_n206), .A3(new_n210), .A4(new_n207), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n201), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT30), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(G137), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n205), .A2(G134), .ZN(new_n216));
  OAI21_X1  g030(.A(G131), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g031(.A1(new_n211), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n219), .A2(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n220), .A2(new_n189), .A3(new_n198), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n191), .A2(G146), .ZN(new_n222));
  OAI21_X1  g036(.A(KEYINPUT64), .B1(new_n188), .B2(G143), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n190), .A2(new_n191), .A3(G146), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n222), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n219), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n221), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n213), .A2(new_n214), .A3(new_n228), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n220), .A2(new_n189), .A3(new_n198), .ZN(new_n230));
  INV_X1    g044(.A(new_n226), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n230), .B1(new_n194), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n211), .A2(new_n217), .ZN(new_n233));
  OAI21_X1  g047(.A(KEYINPUT66), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT66), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n218), .A2(new_n227), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n213), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n229), .B1(KEYINPUT30), .B2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT65), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G116), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n242), .A3(G119), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n239), .A2(G119), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n247), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(new_n243), .A3(new_n245), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n187), .B1(new_n238), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n237), .A2(KEYINPUT30), .ZN(new_n254));
  INV_X1    g068(.A(new_n229), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n256), .A2(KEYINPUT67), .A3(new_n251), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n234), .A2(new_n252), .A3(new_n213), .A4(new_n236), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(KEYINPUT26), .B(G101), .ZN(new_n261));
  INV_X1    g075(.A(G210), .ZN(new_n262));
  NOR3_X1   g076(.A1(new_n262), .A2(G237), .A3(G953), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n261), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n260), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n213), .A2(new_n228), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n259), .B1(new_n269), .B2(new_n252), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT28), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n269), .A2(new_n252), .ZN(new_n272));
  INV_X1    g086(.A(KEYINPUT28), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(new_n267), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(KEYINPUT29), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n268), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n237), .A2(new_n251), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n259), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(KEYINPUT28), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n274), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  AND2_X1   g097(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n284));
  AOI21_X1  g098(.A(G902), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n278), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G472), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n266), .B1(new_n271), .B2(new_n274), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n259), .A2(new_n266), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT69), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT69), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n259), .A2(new_n292), .A3(new_n266), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n253), .B2(new_n257), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT31), .ZN(new_n296));
  OAI21_X1  g110(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT71), .ZN(new_n298));
  XOR2_X1   g112(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n291), .A2(new_n293), .ZN(new_n301));
  AOI21_X1  g115(.A(KEYINPUT67), .B1(new_n256), .B2(new_n251), .ZN(new_n302));
  AOI211_X1 g116(.A(new_n187), .B(new_n252), .C1(new_n254), .C2(new_n255), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n301), .B(new_n299), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(KEYINPUT71), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n297), .B1(new_n300), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g120(.A1(G472), .A2(G902), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n307), .B(KEYINPUT72), .ZN(new_n308));
  NOR3_X1   g122(.A1(new_n306), .A2(KEYINPUT32), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT32), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n301), .B1(new_n302), .B2(new_n303), .ZN(new_n311));
  AOI21_X1  g125(.A(new_n288), .B1(new_n311), .B2(KEYINPUT31), .ZN(new_n312));
  AND4_X1   g126(.A1(new_n298), .A2(new_n258), .A3(new_n301), .A4(new_n299), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n298), .B1(new_n295), .B2(new_n299), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n308), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n310), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n287), .B1(new_n309), .B2(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G137), .ZN(new_n319));
  INV_X1    g133(.A(G221), .ZN(new_n320));
  INV_X1    g134(.A(G234), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n320), .A2(new_n321), .A3(G953), .ZN(new_n322));
  XNOR2_X1  g136(.A(new_n319), .B(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G125), .ZN(new_n325));
  INV_X1    g139(.A(G125), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(G140), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT16), .ZN(new_n328));
  OR3_X1    g142(.A1(new_n326), .A2(KEYINPUT16), .A3(G140), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n328), .A2(G146), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n329), .A3(G146), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT75), .ZN(new_n334));
  AOI21_X1  g148(.A(G146), .B1(new_n328), .B2(new_n329), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  OR2_X1    g151(.A1(new_n219), .A2(G119), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n219), .A2(G119), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g155(.A(KEYINPUT24), .B(G110), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n341), .A2(new_n343), .A3(KEYINPUT74), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT74), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n345), .B1(new_n340), .B2(new_n342), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT23), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n339), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n348), .A2(new_n349), .A3(new_n338), .ZN(new_n350));
  AOI22_X1  g164(.A1(new_n344), .A2(new_n346), .B1(G110), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n337), .A2(new_n351), .ZN(new_n352));
  OAI22_X1  g166(.A1(new_n341), .A2(new_n343), .B1(new_n350), .B2(G110), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n325), .A2(new_n327), .A3(new_n188), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n353), .A2(new_n333), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n323), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n352), .A2(new_n355), .A3(new_n323), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G902), .ZN(new_n360));
  OAI21_X1  g174(.A(G217), .B1(new_n321), .B2(G902), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n361), .B(KEYINPUT73), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n360), .A3(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n363), .A2(KEYINPUT77), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(KEYINPUT77), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n358), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n367), .B2(new_n356), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT25), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT76), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(KEYINPUT25), .B1(new_n359), .B2(new_n360), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT76), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n373), .A3(new_n369), .ZN(new_n374));
  INV_X1    g188(.A(new_n362), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n372), .A2(new_n376), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n366), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g192(.A(KEYINPUT9), .B(G234), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n320), .B1(new_n380), .B2(new_n360), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n382));
  OAI211_X1 g196(.A(KEYINPUT82), .B(KEYINPUT1), .C1(new_n191), .C2(G146), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(KEYINPUT82), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n385));
  OAI21_X1  g199(.A(G128), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n230), .B1(new_n386), .B2(new_n199), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT80), .B(G101), .Z(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(G107), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT79), .B1(new_n390), .B2(G104), .ZN(new_n391));
  INV_X1    g205(.A(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT3), .B1(new_n392), .B2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT79), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n392), .A3(G107), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT3), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n390), .A3(G104), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n391), .A2(new_n393), .A3(new_n395), .A4(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT81), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(new_n390), .B2(G104), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n392), .A2(KEYINPUT81), .A3(G107), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n400), .A2(new_n401), .B1(G104), .B2(new_n390), .ZN(new_n402));
  INV_X1    g216(.A(G101), .ZN(new_n403));
  OAI22_X1  g217(.A1(new_n389), .A2(new_n398), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n382), .B1(new_n387), .B2(new_n404), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n391), .A2(new_n395), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n393), .A2(new_n397), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n388), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n398), .A2(G101), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(KEYINPUT4), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT4), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n398), .A2(new_n411), .A3(G101), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(new_n201), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n398), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n400), .A2(new_n401), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n390), .A2(G104), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g231(.A1(new_n414), .A2(new_n388), .B1(new_n417), .B2(G101), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(KEYINPUT10), .A3(new_n227), .ZN(new_n419));
  AND3_X1   g233(.A1(new_n209), .A2(KEYINPUT84), .A3(new_n211), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT84), .B1(new_n209), .B2(new_n211), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n405), .A2(new_n413), .A3(new_n419), .A4(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n219), .B1(new_n426), .B2(new_n383), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n221), .B1(new_n427), .B2(new_n200), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n418), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n404), .A2(new_n232), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT12), .B1(new_n212), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n431), .A2(new_n212), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n434), .B1(new_n431), .B2(new_n212), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n423), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(G110), .B(G140), .Z(new_n438));
  XNOR2_X1  g252(.A(new_n438), .B(KEYINPUT78), .ZN(new_n439));
  INV_X1    g253(.A(G953), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n440), .A2(G227), .ZN(new_n441));
  XOR2_X1   g255(.A(new_n439), .B(new_n441), .Z(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n423), .A2(new_n442), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n405), .A2(new_n413), .A3(new_n419), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n448));
  AND3_X1   g262(.A1(new_n447), .A2(new_n448), .A3(new_n212), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n448), .B1(new_n447), .B2(new_n212), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n446), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n444), .A2(new_n451), .A3(KEYINPUT87), .ZN(new_n452));
  AOI21_X1  g266(.A(KEYINPUT87), .B1(new_n444), .B2(new_n451), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n360), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(G469), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n423), .B1(new_n449), .B2(new_n450), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n443), .ZN(new_n457));
  INV_X1    g271(.A(new_n212), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n429), .B2(new_n430), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n434), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n446), .ZN(new_n461));
  AOI21_X1  g275(.A(G902), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  XOR2_X1   g276(.A(KEYINPUT88), .B(G469), .Z(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n381), .B1(new_n455), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT96), .ZN(new_n466));
  INV_X1    g280(.A(G237), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(new_n440), .A3(G214), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT93), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G143), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g285(.A1(G237), .A2(G953), .ZN(new_n472));
  OAI211_X1 g286(.A(new_n472), .B(G214), .C1(new_n469), .C2(G143), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G131), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT17), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n471), .A2(new_n473), .A3(new_n210), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n475), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n335), .B1(new_n330), .B2(new_n331), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n210), .B1(new_n471), .B2(new_n473), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT17), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n478), .A2(new_n479), .A3(new_n334), .A4(new_n481), .ZN(new_n482));
  XNOR2_X1  g296(.A(G113), .B(G122), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n483), .B(new_n392), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n474), .A2(KEYINPUT18), .A3(G131), .ZN(new_n485));
  NAND2_X1  g299(.A1(KEYINPUT18), .A2(G131), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n471), .A2(new_n473), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n325), .A2(new_n327), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G146), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n489), .A2(new_n354), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n482), .A2(new_n484), .A3(new_n491), .ZN(new_n492));
  AND3_X1   g306(.A1(new_n325), .A2(new_n327), .A3(KEYINPUT19), .ZN(new_n493));
  AOI21_X1  g307(.A(KEYINPUT19), .B1(new_n325), .B2(new_n327), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n188), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND3_X1   g309(.A1(new_n471), .A2(new_n473), .A3(new_n210), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n495), .B(new_n333), .C1(new_n496), .C2(new_n480), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n497), .A2(new_n491), .A3(KEYINPUT94), .ZN(new_n498));
  INV_X1    g312(.A(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT94), .B1(new_n497), .B2(new_n491), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n492), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(G475), .A2(G902), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n503), .B(KEYINPUT95), .Z(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT20), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT20), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n492), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n484), .B1(new_n482), .B2(new_n491), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n360), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G475), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n466), .B1(new_n509), .B2(new_n513), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n502), .A2(new_n507), .A3(new_n504), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n507), .B1(new_n502), .B2(new_n504), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n513), .B(new_n466), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n514), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT100), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT99), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n191), .A2(G128), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n191), .A2(G128), .ZN(new_n524));
  OR3_X1    g338(.A1(new_n523), .A2(new_n524), .A3(G134), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n240), .A2(new_n242), .A3(G122), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n239), .A2(G122), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n526), .A2(new_n390), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n528), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n390), .B1(new_n526), .B2(new_n527), .ZN(new_n530));
  OAI21_X1  g344(.A(new_n525), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n522), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n533), .A2(KEYINPUT97), .B1(KEYINPUT13), .B2(new_n523), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT97), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n532), .A2(new_n535), .A3(new_n522), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n203), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT14), .ZN(new_n539));
  NAND4_X1  g353(.A1(new_n240), .A2(new_n242), .A3(new_n539), .A4(G122), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(new_n527), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT65), .B(G116), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n539), .B1(new_n542), .B2(G122), .ZN(new_n543));
  OAI21_X1  g357(.A(G107), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT98), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT98), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(G107), .C1(new_n541), .C2(new_n543), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G134), .B1(new_n523), .B2(new_n524), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n529), .B1(new_n525), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n538), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n380), .A2(G217), .A3(new_n440), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n521), .B1(new_n551), .B2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n547), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n526), .A2(KEYINPUT14), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n527), .A3(new_n540), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n546), .B1(new_n557), .B2(G107), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n550), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  OR2_X1    g373(.A1(new_n531), .A2(new_n537), .ZN(new_n560));
  NAND4_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n521), .A4(new_n553), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n525), .A2(new_n549), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n528), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n545), .B2(new_n547), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n552), .B1(new_n564), .B2(new_n538), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n520), .B(new_n360), .C1(new_n554), .C2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(G478), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n559), .A2(new_n560), .A3(new_n553), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(KEYINPUT99), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n561), .A3(new_n565), .ZN(new_n573));
  INV_X1    g387(.A(new_n569), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n520), .A3(new_n360), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  XOR2_X1   g391(.A(KEYINPUT21), .B(G898), .Z(new_n578));
  OAI211_X1 g392(.A(G902), .B(G953), .C1(new_n321), .C2(new_n467), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G952), .ZN(new_n581));
  AOI211_X1 g395(.A(G953), .B(new_n581), .C1(G234), .C2(G237), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n519), .A2(new_n577), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n410), .A2(new_n251), .A3(new_n412), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n243), .A2(KEYINPUT5), .A3(new_n245), .ZN(new_n587));
  INV_X1    g401(.A(G113), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT5), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n588), .B1(new_n244), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n244), .B1(new_n542), .B2(G119), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n587), .A2(new_n590), .B1(new_n591), .B2(new_n249), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n418), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(G110), .B(G122), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n586), .A2(new_n595), .A3(new_n593), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n597), .A2(KEYINPUT6), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n201), .A2(G125), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(G125), .B2(new_n232), .ZN(new_n601));
  INV_X1    g415(.A(G224), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G953), .ZN(new_n603));
  INV_X1    g417(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n601), .B(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT6), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n594), .A2(new_n606), .A3(new_n596), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n599), .A2(new_n605), .A3(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT89), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n599), .A2(KEYINPUT89), .A3(new_n605), .A4(new_n607), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n601), .A2(KEYINPUT7), .A3(new_n604), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n604), .A2(KEYINPUT7), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n600), .B(new_n613), .C1(G125), .C2(new_n232), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n612), .A2(new_n598), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT90), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n418), .B2(new_n592), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n587), .A2(new_n590), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n250), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n619), .A2(KEYINPUT90), .A3(new_n404), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n617), .A2(new_n620), .A3(new_n593), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n595), .B(KEYINPUT8), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(KEYINPUT91), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g438(.A(KEYINPUT91), .B1(new_n621), .B2(new_n622), .ZN(new_n625));
  OAI21_X1  g439(.A(new_n615), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n610), .A2(new_n360), .A3(new_n611), .A4(new_n626), .ZN(new_n627));
  OAI21_X1  g441(.A(G210), .B1(G237), .B2(G902), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(KEYINPUT92), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n625), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n623), .ZN(new_n632));
  AOI21_X1  g446(.A(G902), .B1(new_n632), .B2(new_n615), .ZN(new_n633));
  INV_X1    g447(.A(new_n629), .ZN(new_n634));
  NAND4_X1  g448(.A1(new_n633), .A2(new_n611), .A3(new_n610), .A4(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  OAI21_X1  g450(.A(G214), .B1(G237), .B2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n585), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n318), .A2(new_n378), .A3(new_n465), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(new_n389), .ZN(G3));
  NAND2_X1  g455(.A1(new_n305), .A2(new_n300), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n308), .B1(new_n642), .B2(new_n312), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n315), .A2(new_n360), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n643), .B1(new_n644), .B2(G472), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT101), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n645), .A2(new_n646), .A3(new_n378), .A4(new_n465), .ZN(new_n647));
  AOI21_X1  g461(.A(G902), .B1(new_n642), .B2(new_n312), .ZN(new_n648));
  INV_X1    g462(.A(G472), .ZN(new_n649));
  OAI22_X1  g463(.A1(new_n648), .A2(new_n649), .B1(new_n308), .B2(new_n306), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT87), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n442), .B1(new_n460), .B2(new_n423), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n447), .A2(new_n212), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(KEYINPUT86), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n447), .A2(new_n448), .A3(new_n212), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n445), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n651), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n444), .A2(new_n451), .A3(KEYINPUT87), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G469), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n464), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n381), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n661), .A2(new_n378), .A3(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT101), .B1(new_n650), .B2(new_n663), .ZN(new_n664));
  INV_X1    g478(.A(new_n628), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n627), .A2(new_n665), .ZN(new_n666));
  NAND4_X1  g480(.A1(new_n633), .A2(new_n611), .A3(new_n610), .A4(new_n628), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(KEYINPUT96), .ZN(new_n670));
  INV_X1    g484(.A(KEYINPUT33), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n573), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n565), .A2(new_n571), .A3(KEYINPUT33), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n568), .A2(G902), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n672), .A2(new_n673), .A3(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n573), .A2(new_n360), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n568), .ZN(new_n677));
  AOI22_X1  g491(.A1(new_n670), .A2(new_n517), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n668), .A2(new_n678), .A3(new_n584), .A4(new_n637), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n637), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n666), .B2(new_n667), .ZN(new_n683));
  NAND4_X1  g497(.A1(new_n683), .A2(KEYINPUT102), .A3(new_n584), .A4(new_n678), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n647), .A2(new_n664), .A3(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT34), .B(G104), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G6));
  XNOR2_X1  g502(.A(new_n584), .B(KEYINPUT104), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n683), .A2(new_n689), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT103), .ZN(new_n691));
  AOI22_X1  g505(.A1(new_n506), .A2(new_n508), .B1(new_n513), .B2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n512), .A2(KEYINPUT103), .A3(G475), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n690), .A2(new_n577), .A3(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n647), .A2(new_n664), .A3(new_n695), .ZN(new_n696));
  XOR2_X1   g510(.A(KEYINPUT35), .B(G107), .Z(new_n697));
  XNOR2_X1  g511(.A(new_n696), .B(new_n697), .ZN(G9));
  NAND2_X1  g512(.A1(new_n352), .A2(new_n355), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(KEYINPUT36), .B2(new_n323), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n323), .A2(KEYINPUT36), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n352), .A2(new_n355), .A3(new_n701), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n360), .A3(new_n362), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(KEYINPUT105), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n377), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n645), .A2(new_n639), .A3(new_n465), .A4(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT106), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G12));
  OAI21_X1  g523(.A(new_n583), .B1(new_n579), .B2(G900), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT107), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n576), .A2(new_n693), .A3(new_n692), .A4(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n683), .A2(new_n713), .A3(KEYINPUT108), .ZN(new_n714));
  AND2_X1   g528(.A1(new_n714), .A2(new_n465), .ZN(new_n715));
  AOI21_X1  g529(.A(KEYINPUT108), .B1(new_n683), .B2(new_n713), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n715), .A2(new_n318), .A3(new_n705), .A4(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G128), .ZN(G30));
  XNOR2_X1  g533(.A(new_n636), .B(KEYINPUT38), .ZN(new_n720));
  INV_X1    g534(.A(new_n720), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n670), .A2(new_n517), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n576), .ZN(new_n723));
  NOR4_X1   g537(.A1(new_n721), .A2(new_n682), .A3(new_n705), .A4(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(KEYINPUT32), .B1(new_n306), .B2(new_n308), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n315), .A2(new_n310), .A3(new_n316), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n295), .B1(new_n267), .B2(new_n280), .ZN(new_n728));
  OAI21_X1  g542(.A(G472), .B1(new_n728), .B2(G902), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n727), .A2(KEYINPUT109), .A3(new_n729), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(KEYINPUT110), .B(KEYINPUT39), .Z(new_n735));
  XNOR2_X1  g549(.A(new_n711), .B(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT40), .B1(new_n465), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n465), .A2(new_n737), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT40), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n724), .B(new_n734), .C1(new_n738), .C2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT111), .B(G143), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G45));
  NAND2_X1  g558(.A1(new_n661), .A2(new_n662), .ZN(new_n745));
  INV_X1    g559(.A(new_n683), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n675), .A2(new_n677), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n748), .B(new_n712), .C1(new_n514), .C2(new_n518), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT112), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT112), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n678), .A2(new_n751), .A3(new_n712), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n318), .A2(new_n747), .A3(new_n753), .A4(new_n705), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G146), .ZN(G48));
  AND2_X1   g569(.A1(new_n457), .A2(new_n461), .ZN(new_n756));
  OAI21_X1  g570(.A(G469), .B1(new_n756), .B2(G902), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n757), .A2(new_n662), .A3(new_n464), .ZN(new_n758));
  INV_X1    g572(.A(new_n758), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n685), .A2(new_n318), .A3(new_n378), .A4(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT41), .B(G113), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(G15));
  NAND4_X1  g576(.A1(new_n695), .A2(new_n318), .A3(new_n378), .A4(new_n759), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G116), .ZN(G18));
  INV_X1    g578(.A(new_n585), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n746), .A2(new_n758), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n318), .A2(new_n765), .A3(new_n766), .A4(new_n705), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G119), .ZN(G21));
  NOR3_X1   g582(.A1(new_n690), .A2(new_n758), .A3(new_n723), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n311), .A2(KEYINPUT31), .B1(new_n267), .B2(new_n282), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n308), .B1(new_n642), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g585(.A(KEYINPUT113), .B(G472), .Z(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n771), .B1(new_n644), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n769), .A2(new_n378), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G122), .ZN(G24));
  OAI21_X1  g590(.A(new_n770), .B1(new_n313), .B2(new_n314), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n316), .ZN(new_n778));
  OAI211_X1 g592(.A(new_n778), .B(new_n705), .C1(new_n648), .C2(new_n772), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n780), .A2(new_n753), .A3(new_n766), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(G125), .ZN(G27));
  AOI22_X1  g596(.A1(new_n725), .A2(new_n726), .B1(G472), .B2(new_n286), .ZN(new_n783));
  INV_X1    g597(.A(new_n378), .ZN(new_n784));
  OAI21_X1  g598(.A(KEYINPUT116), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT116), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n318), .A2(new_n786), .A3(new_n378), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n750), .A2(new_n752), .A3(KEYINPUT42), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT114), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n630), .A2(new_n635), .A3(new_n662), .A4(new_n637), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n360), .B1(new_n652), .B2(new_n656), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n462), .A2(new_n463), .B1(G469), .B2(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n630), .A2(new_n637), .A3(new_n635), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n791), .A2(G469), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n464), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(KEYINPUT114), .A3(new_n662), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n788), .B1(new_n793), .B2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n785), .A2(new_n787), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n793), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n800), .A2(new_n318), .A3(new_n378), .A4(new_n753), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT42), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n803), .B1(new_n801), .B2(KEYINPUT115), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n799), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G131), .ZN(G33));
  NAND4_X1  g620(.A1(new_n800), .A2(new_n318), .A3(new_n378), .A4(new_n713), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(G134), .ZN(G36));
  NAND2_X1  g622(.A1(new_n519), .A2(new_n748), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n809), .A2(KEYINPUT43), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT43), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n519), .A2(new_n811), .A3(new_n748), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n810), .A2(new_n705), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  OR3_X1    g628(.A1(new_n813), .A2(new_n814), .A3(new_n645), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n814), .B1(new_n813), .B2(new_n645), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n815), .A2(new_n816), .A3(new_n794), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT117), .ZN(new_n819));
  AOI21_X1  g633(.A(KEYINPUT45), .B1(new_n657), .B2(new_n658), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n819), .B1(new_n820), .B2(new_n660), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT45), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n822), .B1(new_n452), .B2(new_n453), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(KEYINPUT117), .A3(G469), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n444), .A2(new_n451), .A3(KEYINPUT45), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n821), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(G469), .A2(G902), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT46), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n818), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n828), .A2(new_n829), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n826), .A2(KEYINPUT118), .A3(KEYINPUT46), .A4(new_n827), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n830), .A2(new_n831), .A3(new_n464), .A4(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n817), .A2(new_n662), .A3(new_n737), .A4(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(G137), .ZN(G39));
  NAND2_X1  g649(.A1(new_n750), .A2(new_n752), .ZN(new_n836));
  INV_X1    g650(.A(new_n794), .ZN(new_n837));
  NOR4_X1   g651(.A1(new_n318), .A2(new_n836), .A3(new_n378), .A4(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n833), .A2(KEYINPUT47), .A3(new_n662), .ZN(new_n839));
  AOI21_X1  g653(.A(KEYINPUT47), .B1(new_n833), .B2(new_n662), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(G140), .ZN(G42));
  NOR2_X1   g656(.A1(new_n648), .A2(new_n772), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n843), .A2(new_n784), .A3(new_n771), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n810), .A2(new_n582), .A3(new_n812), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n720), .A2(new_n637), .A3(new_n758), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(KEYINPUT50), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n844), .A3(new_n845), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT50), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n757), .A2(new_n464), .ZN(new_n853));
  AND4_X1   g667(.A1(new_n662), .A2(new_n845), .A3(new_n853), .A4(new_n794), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n849), .A2(new_n852), .B1(new_n780), .B2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n853), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n856), .A2(new_n784), .A3(new_n583), .A4(new_n790), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n732), .A2(new_n857), .A3(new_n733), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT122), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n732), .A2(new_n857), .A3(KEYINPUT122), .A4(new_n733), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n722), .A2(new_n748), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n853), .B(KEYINPUT119), .Z(new_n865));
  NOR2_X1   g679(.A1(new_n865), .A2(new_n662), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n839), .A2(new_n840), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n847), .A2(new_n794), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n864), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT51), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n785), .A2(new_n787), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n854), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT48), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n860), .A2(new_n678), .A3(new_n861), .ZN(new_n875));
  AOI211_X1 g689(.A(new_n581), .B(G953), .C1(new_n847), .C2(new_n766), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n874), .A2(new_n875), .A3(new_n876), .ZN(new_n877));
  OAI211_X1 g691(.A(new_n864), .B(KEYINPUT51), .C1(new_n867), .C2(new_n868), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n871), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT54), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n780), .A2(new_n800), .A3(new_n753), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n694), .A2(new_n576), .A3(new_n711), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n794), .A2(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n318), .A2(new_n465), .A3(new_n705), .A4(new_n883), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n807), .A2(new_n881), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT120), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n678), .B1(new_n576), .B2(new_n519), .ZN(new_n887));
  INV_X1    g701(.A(new_n689), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n887), .A2(new_n638), .A3(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n647), .A2(new_n664), .A3(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n890), .A2(new_n760), .A3(new_n763), .ZN(new_n891));
  AND4_X1   g705(.A1(new_n640), .A2(new_n767), .A3(new_n706), .A4(new_n775), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT120), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n807), .A2(new_n881), .A3(new_n884), .A4(new_n893), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n886), .A2(new_n891), .A3(new_n892), .A4(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(new_n799), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n784), .B1(new_n727), .B2(new_n287), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT115), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n898), .A3(new_n753), .A4(new_n800), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n899), .A2(new_n803), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n801), .A2(KEYINPUT115), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n896), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n895), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n377), .A2(new_n704), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n662), .B1(new_n711), .B2(KEYINPUT121), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n905), .B1(KEYINPUT121), .B2(new_n711), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n796), .A2(new_n904), .A3(new_n906), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n907), .A2(new_n746), .A3(new_n723), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n730), .A2(new_n908), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n718), .A2(new_n754), .A3(new_n781), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT52), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n783), .A2(new_n904), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n714), .A2(new_n465), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n914), .A2(new_n716), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n836), .A2(new_n745), .A3(new_n746), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n917), .A2(KEYINPUT52), .A3(new_n781), .A4(new_n909), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n912), .A2(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT53), .B1(new_n903), .B2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n890), .A2(new_n760), .A3(new_n763), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n640), .A2(new_n767), .A3(new_n706), .A4(new_n775), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n805), .A2(new_n923), .A3(new_n886), .A4(new_n894), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT53), .ZN(new_n925));
  AND2_X1   g739(.A1(new_n912), .A2(new_n918), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n880), .B1(new_n920), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n929));
  AND4_X1   g743(.A1(new_n892), .A2(new_n886), .A3(new_n891), .A4(new_n894), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n930), .A2(KEYINPUT53), .A3(new_n805), .A4(new_n919), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n929), .A2(new_n931), .A3(KEYINPUT54), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n879), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g747(.A1(G952), .A2(G953), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n865), .B(KEYINPUT49), .Z(new_n935));
  NOR4_X1   g749(.A1(new_n784), .A2(new_n809), .A3(new_n381), .A4(new_n682), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n935), .A2(new_n721), .A3(new_n936), .ZN(new_n937));
  OAI22_X1  g751(.A1(new_n933), .A2(new_n934), .B1(new_n734), .B2(new_n937), .ZN(G75));
  NAND2_X1  g752(.A1(new_n599), .A2(new_n607), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(new_n605), .Z(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT55), .Z(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI211_X1 g756(.A(new_n262), .B(new_n360), .C1(new_n929), .C2(new_n931), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(KEYINPUT56), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n360), .B1(new_n929), .B2(new_n931), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(G210), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT56), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n947), .A3(new_n941), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n581), .A2(G953), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT123), .Z(new_n950));
  AND3_X1   g764(.A1(new_n944), .A2(new_n948), .A3(new_n950), .ZN(G51));
  INV_X1    g765(.A(new_n950), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n929), .A2(new_n931), .ZN(new_n953));
  INV_X1    g767(.A(new_n826), .ZN(new_n954));
  AND4_X1   g768(.A1(KEYINPUT124), .A2(new_n953), .A3(G902), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT124), .B1(new_n945), .B2(new_n954), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n827), .B(KEYINPUT57), .Z(new_n958));
  NAND3_X1  g772(.A1(new_n928), .A2(new_n932), .A3(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(new_n756), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n952), .B1(new_n957), .B2(new_n961), .ZN(G54));
  NAND3_X1  g776(.A1(new_n945), .A2(KEYINPUT58), .A3(G475), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(new_n502), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n502), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n952), .B1(new_n964), .B2(new_n965), .ZN(G60));
  XNOR2_X1  g780(.A(KEYINPUT125), .B(KEYINPUT59), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n568), .A2(new_n360), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n928), .A2(new_n932), .A3(new_n969), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n672), .A2(new_n673), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n928), .A2(new_n971), .A3(new_n932), .A4(new_n969), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n973), .A2(new_n950), .A3(new_n974), .ZN(G63));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(G217), .A2(G902), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n977), .B(KEYINPUT60), .Z(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(new_n929), .B2(new_n931), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n980), .A2(new_n702), .A3(new_n700), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n950), .B1(new_n980), .B2(new_n359), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OR2_X1    g797(.A1(new_n980), .A2(new_n359), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n980), .A2(new_n702), .A3(new_n700), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(KEYINPUT61), .A3(new_n950), .A4(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(G66));
  NOR2_X1   g801(.A1(new_n602), .A2(new_n440), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n923), .A2(new_n440), .B1(new_n578), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n939), .B1(G898), .B2(new_n440), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  AOI21_X1  g805(.A(new_n440), .B1(G227), .B2(G900), .ZN(new_n992));
  AND2_X1   g806(.A1(new_n917), .A2(new_n781), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n805), .A2(new_n993), .A3(new_n807), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n833), .A2(new_n662), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n995), .A2(new_n736), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n785), .A2(new_n787), .ZN(new_n997));
  NOR3_X1   g811(.A1(new_n997), .A2(new_n746), .A3(new_n723), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n996), .B1(new_n998), .B2(new_n817), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n994), .A2(new_n841), .A3(new_n999), .ZN(new_n1000));
  OR2_X1    g814(.A1(new_n1000), .A2(G953), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n493), .A2(new_n494), .ZN(new_n1002));
  XNOR2_X1  g816(.A(new_n256), .B(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1003), .B1(G900), .B2(G953), .ZN(new_n1004));
  AND2_X1   g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1003), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n993), .A2(new_n742), .ZN(new_n1007));
  XOR2_X1   g821(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n1008));
  NAND2_X1  g822(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND4_X1  g823(.A1(new_n993), .A2(new_n742), .A3(KEYINPUT126), .A4(KEYINPUT62), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n739), .A2(new_n837), .A3(new_n887), .ZN(new_n1012));
  AOI22_X1  g826(.A1(new_n996), .A2(new_n817), .B1(new_n897), .B2(new_n1012), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1013), .A3(new_n841), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1006), .B1(new_n1014), .B2(new_n440), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n992), .B1(new_n1005), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1017));
  INV_X1    g831(.A(new_n992), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1016), .A2(new_n1019), .ZN(G72));
  NAND4_X1  g834(.A1(new_n1011), .A2(new_n1013), .A3(new_n841), .A4(new_n923), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  NAND2_X1  g837(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n267), .B1(new_n258), .B2(new_n259), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g840(.A(new_n923), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1023), .B1(new_n1000), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g842(.A1(new_n260), .A2(new_n266), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1026), .A2(new_n1030), .A3(new_n950), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n268), .A2(new_n311), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n953), .A2(new_n1023), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g847(.A(KEYINPUT127), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OR2_X1    g849(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n1031), .B1(new_n1035), .B2(new_n1036), .ZN(G57));
endmodule


