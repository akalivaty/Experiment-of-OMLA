

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589;

  XNOR2_X1 U325 ( .A(n477), .B(n476), .ZN(n545) );
  XNOR2_X1 U326 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n476) );
  XNOR2_X1 U327 ( .A(n395), .B(n394), .ZN(n398) );
  XNOR2_X1 U328 ( .A(KEYINPUT118), .B(KEYINPUT47), .ZN(n469) );
  NOR2_X1 U329 ( .A1(n547), .A2(n431), .ZN(n432) );
  XNOR2_X1 U330 ( .A(n470), .B(n469), .ZN(n475) );
  INV_X1 U331 ( .A(KEYINPUT99), .ZN(n392) );
  INV_X1 U332 ( .A(KEYINPUT31), .ZN(n319) );
  XNOR2_X1 U333 ( .A(n458), .B(KEYINPUT110), .ZN(n459) );
  XNOR2_X1 U334 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U335 ( .A(n320), .B(n319), .ZN(n321) );
  XNOR2_X1 U336 ( .A(n460), .B(n459), .ZN(n502) );
  XNOR2_X1 U337 ( .A(n322), .B(n321), .ZN(n323) );
  NOR2_X1 U338 ( .A1(n566), .A2(n565), .ZN(n575) );
  XNOR2_X1 U339 ( .A(n400), .B(n399), .ZN(n526) );
  XNOR2_X1 U340 ( .A(n462), .B(G106GAT), .ZN(n463) );
  XNOR2_X1 U341 ( .A(n464), .B(n463), .ZN(G1339GAT) );
  XOR2_X1 U342 ( .A(KEYINPUT22), .B(KEYINPUT91), .Z(n294) );
  XNOR2_X1 U343 ( .A(KEYINPUT90), .B(KEYINPUT24), .ZN(n293) );
  XNOR2_X1 U344 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U345 ( .A(G204GAT), .B(KEYINPUT23), .Z(n296) );
  XOR2_X1 U346 ( .A(G141GAT), .B(G22GAT), .Z(n330) );
  XOR2_X1 U347 ( .A(G50GAT), .B(G162GAT), .Z(n359) );
  XNOR2_X1 U348 ( .A(n330), .B(n359), .ZN(n295) );
  XNOR2_X1 U349 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U350 ( .A(n298), .B(n297), .Z(n300) );
  NAND2_X1 U351 ( .A1(G228GAT), .A2(G233GAT), .ZN(n299) );
  XNOR2_X1 U352 ( .A(n300), .B(n299), .ZN(n303) );
  XOR2_X1 U353 ( .A(G155GAT), .B(KEYINPUT2), .Z(n302) );
  XNOR2_X1 U354 ( .A(KEYINPUT3), .B(KEYINPUT94), .ZN(n301) );
  XNOR2_X1 U355 ( .A(n302), .B(n301), .ZN(n369) );
  XOR2_X1 U356 ( .A(n303), .B(n369), .Z(n310) );
  XNOR2_X1 U357 ( .A(G211GAT), .B(KEYINPUT21), .ZN(n304) );
  XNOR2_X1 U358 ( .A(n304), .B(KEYINPUT92), .ZN(n305) );
  XOR2_X1 U359 ( .A(n305), .B(KEYINPUT93), .Z(n307) );
  XNOR2_X1 U360 ( .A(G197GAT), .B(G218GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n390) );
  XNOR2_X1 U362 ( .A(G106GAT), .B(G78GAT), .ZN(n308) );
  XNOR2_X1 U363 ( .A(n308), .B(G148GAT), .ZN(n316) );
  XNOR2_X1 U364 ( .A(n390), .B(n316), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n561) );
  XOR2_X1 U366 ( .A(n561), .B(KEYINPUT28), .Z(n521) );
  XOR2_X1 U367 ( .A(G120GAT), .B(G71GAT), .Z(n413) );
  XOR2_X1 U368 ( .A(G99GAT), .B(G85GAT), .Z(n358) );
  XNOR2_X1 U369 ( .A(n413), .B(n358), .ZN(n324) );
  XOR2_X1 U370 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n312) );
  NAND2_X1 U371 ( .A1(G230GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U372 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U373 ( .A(n313), .B(KEYINPUT69), .Z(n318) );
  XOR2_X1 U374 ( .A(G64GAT), .B(G92GAT), .Z(n315) );
  XNOR2_X1 U375 ( .A(G176GAT), .B(G204GAT), .ZN(n314) );
  XNOR2_X1 U376 ( .A(n315), .B(n314), .ZN(n391) );
  XNOR2_X1 U377 ( .A(n391), .B(n316), .ZN(n317) );
  XNOR2_X1 U378 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT13), .Z(n438) );
  XNOR2_X1 U380 ( .A(n438), .B(KEYINPUT70), .ZN(n320) );
  XOR2_X1 U381 ( .A(n324), .B(n323), .Z(n584) );
  XOR2_X1 U382 ( .A(n584), .B(KEYINPUT41), .Z(n549) );
  XOR2_X1 U383 ( .A(KEYINPUT66), .B(KEYINPUT67), .Z(n326) );
  XNOR2_X1 U384 ( .A(G1GAT), .B(G8GAT), .ZN(n325) );
  XNOR2_X1 U385 ( .A(n326), .B(n325), .ZN(n343) );
  XOR2_X1 U386 ( .A(G113GAT), .B(G197GAT), .Z(n328) );
  XNOR2_X1 U387 ( .A(G36GAT), .B(G50GAT), .ZN(n327) );
  XNOR2_X1 U388 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U389 ( .A(n329), .B(G15GAT), .Z(n332) );
  XNOR2_X1 U390 ( .A(G169GAT), .B(n330), .ZN(n331) );
  XNOR2_X1 U391 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U392 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n334) );
  NAND2_X1 U393 ( .A1(G229GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U394 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U395 ( .A(n336), .B(n335), .Z(n341) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n338) );
  XNOR2_X1 U397 ( .A(G43GAT), .B(G29GAT), .ZN(n337) );
  XNOR2_X1 U398 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U399 ( .A(KEYINPUT7), .B(n339), .Z(n363) );
  XNOR2_X1 U400 ( .A(n363), .B(KEYINPUT65), .ZN(n340) );
  XNOR2_X1 U401 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U402 ( .A(n343), .B(n342), .ZN(n579) );
  INV_X1 U403 ( .A(n579), .ZN(n567) );
  NOR2_X1 U404 ( .A1(n549), .A2(n567), .ZN(n344) );
  XNOR2_X1 U405 ( .A(n344), .B(KEYINPUT114), .ZN(n514) );
  XOR2_X1 U406 ( .A(G92GAT), .B(G106GAT), .Z(n346) );
  XNOR2_X1 U407 ( .A(G134GAT), .B(G218GAT), .ZN(n345) );
  XNOR2_X1 U408 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U409 ( .A(KEYINPUT9), .B(KEYINPUT73), .Z(n348) );
  XNOR2_X1 U410 ( .A(KEYINPUT72), .B(KEYINPUT10), .ZN(n347) );
  XNOR2_X1 U411 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U412 ( .A(n350), .B(n349), .Z(n355) );
  XOR2_X1 U413 ( .A(KEYINPUT74), .B(KEYINPUT11), .Z(n352) );
  NAND2_X1 U414 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U416 ( .A(KEYINPUT76), .B(n353), .ZN(n354) );
  XNOR2_X1 U417 ( .A(n355), .B(n354), .ZN(n357) );
  XNOR2_X1 U418 ( .A(G36GAT), .B(G190GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n356), .B(KEYINPUT75), .ZN(n396) );
  XOR2_X1 U420 ( .A(n357), .B(n396), .Z(n361) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U423 ( .A(n363), .B(n362), .Z(n576) );
  XOR2_X1 U424 ( .A(KEYINPUT36), .B(n576), .Z(n484) );
  XOR2_X1 U425 ( .A(KEYINPUT6), .B(G57GAT), .Z(n365) );
  XNOR2_X1 U426 ( .A(G1GAT), .B(G120GAT), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n373) );
  XOR2_X1 U428 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n371) );
  XOR2_X1 U429 ( .A(KEYINPUT0), .B(G134GAT), .Z(n367) );
  XNOR2_X1 U430 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U432 ( .A(G113GAT), .B(n368), .Z(n417) );
  XNOR2_X1 U433 ( .A(n417), .B(n369), .ZN(n370) );
  XNOR2_X1 U434 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U435 ( .A(n373), .B(n372), .ZN(n385) );
  NAND2_X1 U436 ( .A1(G225GAT), .A2(G233GAT), .ZN(n379) );
  XOR2_X1 U437 ( .A(G162GAT), .B(G148GAT), .Z(n375) );
  XNOR2_X1 U438 ( .A(G141GAT), .B(G127GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U440 ( .A(G29GAT), .B(G85GAT), .Z(n376) );
  XNOR2_X1 U441 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n383) );
  XOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT97), .Z(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n380) );
  XNOR2_X1 U445 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U446 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n559) );
  INV_X1 U448 ( .A(n521), .ZN(n386) );
  NOR2_X1 U449 ( .A1(n559), .A2(n386), .ZN(n403) );
  XOR2_X1 U450 ( .A(KEYINPUT17), .B(KEYINPUT19), .Z(n388) );
  XNOR2_X1 U451 ( .A(KEYINPUT18), .B(G183GAT), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U453 ( .A(G169GAT), .B(n389), .Z(n410) );
  XNOR2_X1 U454 ( .A(n410), .B(n390), .ZN(n400) );
  XOR2_X1 U455 ( .A(G8GAT), .B(KEYINPUT77), .Z(n442) );
  XOR2_X1 U456 ( .A(n442), .B(n391), .Z(n395) );
  NAND2_X1 U457 ( .A1(G226GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n396), .B(KEYINPUT98), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U460 ( .A(n526), .B(KEYINPUT27), .Z(n401) );
  XOR2_X1 U461 ( .A(KEYINPUT100), .B(n401), .Z(n426) );
  INV_X1 U462 ( .A(n426), .ZN(n402) );
  NAND2_X1 U463 ( .A1(n403), .A2(n402), .ZN(n530) );
  XNOR2_X1 U464 ( .A(n530), .B(KEYINPUT101), .ZN(n422) );
  XOR2_X1 U465 ( .A(KEYINPUT89), .B(KEYINPUT20), .Z(n405) );
  XNOR2_X1 U466 ( .A(KEYINPUT87), .B(KEYINPUT84), .ZN(n404) );
  XNOR2_X1 U467 ( .A(n405), .B(n404), .ZN(n406) );
  XOR2_X1 U468 ( .A(G176GAT), .B(n406), .Z(n408) );
  NAND2_X1 U469 ( .A1(G227GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U470 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U471 ( .A(n409), .B(KEYINPUT85), .Z(n412) );
  XNOR2_X1 U472 ( .A(n410), .B(KEYINPUT88), .ZN(n411) );
  XNOR2_X1 U473 ( .A(n412), .B(n411), .ZN(n421) );
  XOR2_X1 U474 ( .A(KEYINPUT86), .B(G190GAT), .Z(n415) );
  XOR2_X1 U475 ( .A(G15GAT), .B(G127GAT), .Z(n452) );
  XNOR2_X1 U476 ( .A(n452), .B(n413), .ZN(n414) );
  XNOR2_X1 U477 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(n416), .B(G99GAT), .Z(n419) );
  XNOR2_X1 U479 ( .A(G43GAT), .B(n417), .ZN(n418) );
  XNOR2_X1 U480 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U481 ( .A(n421), .B(n420), .ZN(n532) );
  INV_X1 U482 ( .A(n532), .ZN(n566) );
  NAND2_X1 U483 ( .A1(n422), .A2(n566), .ZN(n423) );
  XNOR2_X1 U484 ( .A(n423), .B(KEYINPUT102), .ZN(n435) );
  XOR2_X1 U485 ( .A(KEYINPUT26), .B(KEYINPUT103), .Z(n425) );
  NAND2_X1 U486 ( .A1(n561), .A2(n566), .ZN(n424) );
  XNOR2_X1 U487 ( .A(n425), .B(n424), .ZN(n480) );
  NOR2_X1 U488 ( .A1(n480), .A2(n426), .ZN(n547) );
  XNOR2_X1 U489 ( .A(KEYINPUT25), .B(KEYINPUT105), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n427), .B(KEYINPUT104), .ZN(n430) );
  NOR2_X1 U491 ( .A1(n566), .A2(n526), .ZN(n428) );
  NOR2_X1 U492 ( .A1(n561), .A2(n428), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U494 ( .A(KEYINPUT106), .B(n432), .Z(n433) );
  NAND2_X1 U495 ( .A1(n559), .A2(n433), .ZN(n434) );
  NAND2_X1 U496 ( .A1(n435), .A2(n434), .ZN(n491) );
  XOR2_X1 U497 ( .A(G78GAT), .B(G211GAT), .Z(n437) );
  XNOR2_X1 U498 ( .A(G183GAT), .B(G71GAT), .ZN(n436) );
  XNOR2_X1 U499 ( .A(n437), .B(n436), .ZN(n439) );
  XOR2_X1 U500 ( .A(n439), .B(n438), .Z(n441) );
  XNOR2_X1 U501 ( .A(G22GAT), .B(G155GAT), .ZN(n440) );
  XNOR2_X1 U502 ( .A(n441), .B(n440), .ZN(n456) );
  XOR2_X1 U503 ( .A(n442), .B(KEYINPUT81), .Z(n444) );
  NAND2_X1 U504 ( .A1(G231GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U505 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U506 ( .A(KEYINPUT15), .B(KEYINPUT12), .Z(n446) );
  XNOR2_X1 U507 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n445) );
  XNOR2_X1 U508 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U509 ( .A(n448), .B(n447), .Z(n454) );
  XOR2_X1 U510 ( .A(KEYINPUT78), .B(KEYINPUT79), .Z(n450) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(KEYINPUT80), .ZN(n449) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U515 ( .A(n456), .B(n455), .ZN(n587) );
  NAND2_X1 U516 ( .A1(n491), .A2(n587), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n484), .A2(n457), .ZN(n460) );
  XNOR2_X1 U518 ( .A(KEYINPUT37), .B(KEYINPUT109), .ZN(n458) );
  NAND2_X1 U519 ( .A1(n514), .A2(n502), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT116), .ZN(n528) );
  NOR2_X1 U521 ( .A1(n521), .A2(n528), .ZN(n464) );
  XNOR2_X1 U522 ( .A(KEYINPUT117), .B(KEYINPUT44), .ZN(n462) );
  INV_X1 U523 ( .A(G218GAT), .ZN(n487) );
  OR2_X1 U524 ( .A1(n549), .A2(n579), .ZN(n466) );
  INV_X1 U525 ( .A(KEYINPUT46), .ZN(n465) );
  XNOR2_X1 U526 ( .A(n466), .B(n465), .ZN(n468) );
  INV_X1 U527 ( .A(n576), .ZN(n557) );
  NAND2_X1 U528 ( .A1(n557), .A2(n587), .ZN(n467) );
  OR2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n470) );
  NOR2_X1 U530 ( .A1(n484), .A2(n587), .ZN(n471) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT45), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n472), .A2(n584), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n473), .A2(n567), .ZN(n474) );
  NOR2_X1 U534 ( .A1(n475), .A2(n474), .ZN(n477) );
  XOR2_X1 U535 ( .A(KEYINPUT125), .B(n526), .Z(n478) );
  NOR2_X1 U536 ( .A1(n545), .A2(n478), .ZN(n479) );
  XNOR2_X1 U537 ( .A(n479), .B(KEYINPUT54), .ZN(n563) );
  INV_X1 U538 ( .A(n480), .ZN(n481) );
  AND2_X1 U539 ( .A1(n559), .A2(n481), .ZN(n482) );
  AND2_X1 U540 ( .A1(n563), .A2(n482), .ZN(n483) );
  XOR2_X1 U541 ( .A(n483), .B(KEYINPUT126), .Z(n588) );
  NOR2_X1 U542 ( .A1(n484), .A2(n588), .ZN(n485) );
  XNOR2_X1 U543 ( .A(KEYINPUT62), .B(n485), .ZN(n486) );
  XNOR2_X1 U544 ( .A(n487), .B(n486), .ZN(G1355GAT) );
  NAND2_X1 U545 ( .A1(n584), .A2(n567), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n488), .B(KEYINPUT71), .ZN(n501) );
  INV_X1 U547 ( .A(n587), .ZN(n573) );
  NAND2_X1 U548 ( .A1(n573), .A2(n557), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT16), .B(n489), .Z(n490) );
  AND2_X1 U550 ( .A1(n491), .A2(n490), .ZN(n515) );
  NAND2_X1 U551 ( .A1(n501), .A2(n515), .ZN(n492) );
  XOR2_X1 U552 ( .A(KEYINPUT107), .B(n492), .Z(n499) );
  NOR2_X1 U553 ( .A1(n559), .A2(n499), .ZN(n494) );
  XNOR2_X1 U554 ( .A(KEYINPUT34), .B(KEYINPUT108), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(n495) );
  XOR2_X1 U556 ( .A(G1GAT), .B(n495), .Z(G1324GAT) );
  NOR2_X1 U557 ( .A1(n526), .A2(n499), .ZN(n496) );
  XOR2_X1 U558 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U559 ( .A1(n566), .A2(n499), .ZN(n498) );
  XNOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n521), .A2(n499), .ZN(n500) );
  XOR2_X1 U563 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NAND2_X1 U564 ( .A1(n502), .A2(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT38), .ZN(n512) );
  NOR2_X1 U566 ( .A1(n512), .A2(n559), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(KEYINPUT39), .ZN(n505) );
  XNOR2_X1 U568 ( .A(G29GAT), .B(n505), .ZN(G1328GAT) );
  NOR2_X1 U569 ( .A1(n526), .A2(n512), .ZN(n506) );
  XOR2_X1 U570 ( .A(G36GAT), .B(n506), .Z(G1329GAT) );
  XOR2_X1 U571 ( .A(KEYINPUT40), .B(KEYINPUT113), .Z(n508) );
  XNOR2_X1 U572 ( .A(G43GAT), .B(KEYINPUT112), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT111), .B(n509), .ZN(n511) );
  NOR2_X1 U575 ( .A1(n566), .A2(n512), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1330GAT) );
  NOR2_X1 U577 ( .A1(n521), .A2(n512), .ZN(n513) );
  XOR2_X1 U578 ( .A(G50GAT), .B(n513), .Z(G1331GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n559), .A2(n520), .ZN(n516) );
  XOR2_X1 U581 ( .A(G57GAT), .B(n516), .Z(n517) );
  XNOR2_X1 U582 ( .A(KEYINPUT42), .B(n517), .ZN(G1332GAT) );
  NOR2_X1 U583 ( .A1(n526), .A2(n520), .ZN(n518) );
  XOR2_X1 U584 ( .A(G64GAT), .B(n518), .Z(G1333GAT) );
  NOR2_X1 U585 ( .A1(n566), .A2(n520), .ZN(n519) );
  XOR2_X1 U586 ( .A(G71GAT), .B(n519), .Z(G1334GAT) );
  NOR2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U588 ( .A(KEYINPUT43), .B(KEYINPUT115), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(n524) );
  XOR2_X1 U590 ( .A(G78GAT), .B(n524), .Z(G1335GAT) );
  NOR2_X1 U591 ( .A1(n559), .A2(n528), .ZN(n525) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n528), .ZN(n527) );
  XOR2_X1 U594 ( .A(G92GAT), .B(n527), .Z(G1337GAT) );
  NOR2_X1 U595 ( .A1(n566), .A2(n528), .ZN(n529) );
  XOR2_X1 U596 ( .A(G99GAT), .B(n529), .Z(G1338GAT) );
  NOR2_X1 U597 ( .A1(n545), .A2(n530), .ZN(n531) );
  NAND2_X1 U598 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n533), .B(KEYINPUT119), .ZN(n542) );
  NAND2_X1 U600 ( .A1(n567), .A2(n542), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G113GAT), .B(n534), .ZN(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT120), .Z(n536) );
  INV_X1 U603 ( .A(n549), .ZN(n569) );
  NAND2_X1 U604 ( .A1(n542), .A2(n569), .ZN(n535) );
  XNOR2_X1 U605 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n537), .ZN(G1341GAT) );
  XNOR2_X1 U607 ( .A(G127GAT), .B(KEYINPUT50), .ZN(n541) );
  XOR2_X1 U608 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n539) );
  NAND2_X1 U609 ( .A1(n542), .A2(n573), .ZN(n538) );
  XNOR2_X1 U610 ( .A(n539), .B(n538), .ZN(n540) );
  XNOR2_X1 U611 ( .A(n541), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(G134GAT), .B(KEYINPUT51), .Z(n544) );
  NAND2_X1 U613 ( .A1(n542), .A2(n576), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n544), .B(n543), .ZN(G1343GAT) );
  NOR2_X1 U615 ( .A1(n559), .A2(n545), .ZN(n546) );
  NAND2_X1 U616 ( .A1(n547), .A2(n546), .ZN(n556) );
  NOR2_X1 U617 ( .A1(n579), .A2(n556), .ZN(n548) );
  XOR2_X1 U618 ( .A(G141GAT), .B(n548), .Z(G1344GAT) );
  NOR2_X1 U619 ( .A1(n556), .A2(n549), .ZN(n553) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n551) );
  XNOR2_X1 U621 ( .A(G148GAT), .B(KEYINPUT123), .ZN(n550) );
  XNOR2_X1 U622 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U623 ( .A(n553), .B(n552), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n587), .A2(n556), .ZN(n554) );
  XOR2_X1 U625 ( .A(KEYINPUT124), .B(n554), .Z(n555) );
  XNOR2_X1 U626 ( .A(G155GAT), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n558), .Z(G1347GAT) );
  INV_X1 U629 ( .A(n559), .ZN(n560) );
  NOR2_X1 U630 ( .A1(n561), .A2(n560), .ZN(n562) );
  AND2_X1 U631 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n564), .B(KEYINPUT55), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n575), .A2(n567), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U635 ( .A1(n575), .A2(n569), .ZN(n571) );
  XOR2_X1 U636 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G176GAT), .ZN(G1349GAT) );
  NAND2_X1 U639 ( .A1(n575), .A2(n573), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U641 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1351GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n588), .ZN(n583) );
  XOR2_X1 U645 ( .A(KEYINPUT127), .B(KEYINPUT59), .Z(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n588), .A2(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n585) );
  XNOR2_X1 U651 ( .A(n586), .B(n585), .ZN(G1353GAT) );
  NOR2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n589) );
  XOR2_X1 U653 ( .A(G211GAT), .B(n589), .Z(G1354GAT) );
endmodule

