

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U552 ( .A1(G2104), .A2(n525), .ZN(n583) );
  XNOR2_X1 U553 ( .A(n719), .B(KEYINPUT30), .ZN(n720) );
  XNOR2_X1 U554 ( .A(n721), .B(n720), .ZN(n722) );
  INV_X1 U555 ( .A(KEYINPUT31), .ZN(n729) );
  XNOR2_X1 U556 ( .A(n763), .B(KEYINPUT97), .ZN(n764) );
  XNOR2_X1 U557 ( .A(n765), .B(n764), .ZN(n795) );
  XOR2_X1 U558 ( .A(KEYINPUT1), .B(n515), .Z(n635) );
  XOR2_X1 U559 ( .A(G543), .B(KEYINPUT0), .Z(n613) );
  NOR2_X1 U560 ( .A1(G651), .A2(n613), .ZN(n628) );
  NAND2_X1 U561 ( .A1(G52), .A2(n628), .ZN(n517) );
  INV_X1 U562 ( .A(G651), .ZN(n519) );
  NOR2_X1 U563 ( .A1(G543), .A2(n519), .ZN(n515) );
  NAND2_X1 U564 ( .A1(G64), .A2(n635), .ZN(n516) );
  NAND2_X1 U565 ( .A1(n517), .A2(n516), .ZN(n518) );
  XOR2_X1 U566 ( .A(KEYINPUT67), .B(n518), .Z(n524) );
  NOR2_X1 U567 ( .A1(G543), .A2(G651), .ZN(n627) );
  NAND2_X1 U568 ( .A1(G90), .A2(n627), .ZN(n521) );
  NOR2_X1 U569 ( .A1(n613), .A2(n519), .ZN(n631) );
  NAND2_X1 U570 ( .A1(G77), .A2(n631), .ZN(n520) );
  NAND2_X1 U571 ( .A1(n521), .A2(n520), .ZN(n522) );
  XOR2_X1 U572 ( .A(KEYINPUT9), .B(n522), .Z(n523) );
  NOR2_X1 U573 ( .A1(n524), .A2(n523), .ZN(G171) );
  AND2_X1 U574 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U575 ( .A(G57), .ZN(G237) );
  INV_X1 U576 ( .A(G132), .ZN(G219) );
  INV_X1 U577 ( .A(G82), .ZN(G220) );
  INV_X1 U578 ( .A(G2105), .ZN(n525) );
  NAND2_X1 U579 ( .A1(G125), .A2(n583), .ZN(n527) );
  AND2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n873) );
  NAND2_X1 U581 ( .A1(G113), .A2(n873), .ZN(n526) );
  NAND2_X1 U582 ( .A1(n527), .A2(n526), .ZN(n671) );
  NAND2_X1 U583 ( .A1(n525), .A2(G2104), .ZN(n528) );
  XNOR2_X1 U584 ( .A(n528), .B(KEYINPUT65), .ZN(n589) );
  NAND2_X1 U585 ( .A1(G101), .A2(n589), .ZN(n529) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(n529), .Z(n676) );
  NOR2_X1 U587 ( .A1(G2105), .A2(G2104), .ZN(n530) );
  XOR2_X1 U588 ( .A(KEYINPUT17), .B(n530), .Z(n585) );
  NAND2_X1 U589 ( .A1(n585), .A2(G137), .ZN(n674) );
  NAND2_X1 U590 ( .A1(n676), .A2(n674), .ZN(n531) );
  NOR2_X1 U591 ( .A1(n671), .A2(n531), .ZN(G160) );
  NAND2_X1 U592 ( .A1(G7), .A2(G661), .ZN(n532) );
  XNOR2_X1 U593 ( .A(n532), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U594 ( .A(G223), .ZN(n835) );
  NAND2_X1 U595 ( .A1(n835), .A2(G567), .ZN(n533) );
  XOR2_X1 U596 ( .A(KEYINPUT11), .B(n533), .Z(G234) );
  NAND2_X1 U597 ( .A1(G81), .A2(n627), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n534), .B(KEYINPUT12), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT70), .ZN(n537) );
  NAND2_X1 U600 ( .A1(G68), .A2(n631), .ZN(n536) );
  NAND2_X1 U601 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U602 ( .A(n538), .B(KEYINPUT13), .ZN(n540) );
  NAND2_X1 U603 ( .A1(G43), .A2(n628), .ZN(n539) );
  NAND2_X1 U604 ( .A1(n540), .A2(n539), .ZN(n543) );
  NAND2_X1 U605 ( .A1(n635), .A2(G56), .ZN(n541) );
  XOR2_X1 U606 ( .A(KEYINPUT14), .B(n541), .Z(n542) );
  NOR2_X1 U607 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(KEYINPUT71), .B(n544), .ZN(n992) );
  INV_X1 U609 ( .A(n992), .ZN(n545) );
  NAND2_X1 U610 ( .A1(n545), .A2(G860), .ZN(G153) );
  INV_X1 U611 ( .A(G171), .ZN(G301) );
  NAND2_X1 U612 ( .A1(G868), .A2(G301), .ZN(n556) );
  NAND2_X1 U613 ( .A1(G79), .A2(n631), .ZN(n546) );
  XNOR2_X1 U614 ( .A(n546), .B(KEYINPUT72), .ZN(n553) );
  NAND2_X1 U615 ( .A1(G92), .A2(n627), .ZN(n548) );
  NAND2_X1 U616 ( .A1(G66), .A2(n635), .ZN(n547) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U618 ( .A1(G54), .A2(n628), .ZN(n549) );
  XNOR2_X1 U619 ( .A(KEYINPUT73), .B(n549), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U622 ( .A(KEYINPUT15), .B(n554), .Z(n974) );
  INV_X1 U623 ( .A(G868), .ZN(n645) );
  NAND2_X1 U624 ( .A1(n974), .A2(n645), .ZN(n555) );
  NAND2_X1 U625 ( .A1(n556), .A2(n555), .ZN(G284) );
  NAND2_X1 U626 ( .A1(n627), .A2(G89), .ZN(n557) );
  XNOR2_X1 U627 ( .A(n557), .B(KEYINPUT4), .ZN(n559) );
  NAND2_X1 U628 ( .A1(G76), .A2(n631), .ZN(n558) );
  NAND2_X1 U629 ( .A1(n559), .A2(n558), .ZN(n560) );
  XNOR2_X1 U630 ( .A(n560), .B(KEYINPUT5), .ZN(n565) );
  NAND2_X1 U631 ( .A1(G51), .A2(n628), .ZN(n562) );
  NAND2_X1 U632 ( .A1(G63), .A2(n635), .ZN(n561) );
  NAND2_X1 U633 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U634 ( .A(KEYINPUT6), .B(n563), .Z(n564) );
  NAND2_X1 U635 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U636 ( .A(n566), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U637 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U638 ( .A1(n635), .A2(G65), .ZN(n573) );
  NAND2_X1 U639 ( .A1(G91), .A2(n627), .ZN(n568) );
  NAND2_X1 U640 ( .A1(G53), .A2(n628), .ZN(n567) );
  NAND2_X1 U641 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U642 ( .A1(n631), .A2(G78), .ZN(n569) );
  XOR2_X1 U643 ( .A(KEYINPUT68), .B(n569), .Z(n570) );
  NOR2_X1 U644 ( .A1(n571), .A2(n570), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U646 ( .A(KEYINPUT69), .B(n574), .Z(G299) );
  NAND2_X1 U647 ( .A1(G286), .A2(G868), .ZN(n576) );
  NAND2_X1 U648 ( .A1(G299), .A2(n645), .ZN(n575) );
  NAND2_X1 U649 ( .A1(n576), .A2(n575), .ZN(G297) );
  INV_X1 U650 ( .A(G559), .ZN(n579) );
  NOR2_X1 U651 ( .A1(G860), .A2(n579), .ZN(n577) );
  NOR2_X1 U652 ( .A1(n974), .A2(n577), .ZN(n578) );
  XOR2_X1 U653 ( .A(KEYINPUT16), .B(n578), .Z(G148) );
  INV_X1 U654 ( .A(n974), .ZN(n602) );
  NAND2_X1 U655 ( .A1(n579), .A2(n602), .ZN(n580) );
  NAND2_X1 U656 ( .A1(n580), .A2(G868), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n992), .A2(n645), .ZN(n581) );
  NAND2_X1 U658 ( .A1(n582), .A2(n581), .ZN(G282) );
  NAND2_X1 U659 ( .A1(n583), .A2(G123), .ZN(n584) );
  XNOR2_X1 U660 ( .A(n584), .B(KEYINPUT18), .ZN(n587) );
  BUF_X1 U661 ( .A(n585), .Z(n876) );
  NAND2_X1 U662 ( .A1(G135), .A2(n876), .ZN(n586) );
  NAND2_X1 U663 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U664 ( .A(KEYINPUT74), .B(n588), .ZN(n593) );
  BUF_X1 U665 ( .A(n589), .Z(n878) );
  NAND2_X1 U666 ( .A1(G99), .A2(n878), .ZN(n591) );
  NAND2_X1 U667 ( .A1(G111), .A2(n873), .ZN(n590) );
  NAND2_X1 U668 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U669 ( .A1(n593), .A2(n592), .ZN(n947) );
  XNOR2_X1 U670 ( .A(G2096), .B(n947), .ZN(n595) );
  INV_X1 U671 ( .A(G2100), .ZN(n594) );
  NAND2_X1 U672 ( .A1(n595), .A2(n594), .ZN(G156) );
  NAND2_X1 U673 ( .A1(G93), .A2(n627), .ZN(n597) );
  NAND2_X1 U674 ( .A1(G80), .A2(n631), .ZN(n596) );
  NAND2_X1 U675 ( .A1(n597), .A2(n596), .ZN(n601) );
  NAND2_X1 U676 ( .A1(G55), .A2(n628), .ZN(n599) );
  NAND2_X1 U677 ( .A1(G67), .A2(n635), .ZN(n598) );
  NAND2_X1 U678 ( .A1(n599), .A2(n598), .ZN(n600) );
  OR2_X1 U679 ( .A1(n601), .A2(n600), .ZN(n646) );
  NAND2_X1 U680 ( .A1(G559), .A2(n602), .ZN(n603) );
  XNOR2_X1 U681 ( .A(n603), .B(n992), .ZN(n643) );
  NOR2_X1 U682 ( .A1(G860), .A2(n643), .ZN(n604) );
  XOR2_X1 U683 ( .A(KEYINPUT75), .B(n604), .Z(n605) );
  XOR2_X1 U684 ( .A(n646), .B(n605), .Z(G145) );
  NAND2_X1 U685 ( .A1(G50), .A2(n628), .ZN(n607) );
  NAND2_X1 U686 ( .A1(G62), .A2(n635), .ZN(n606) );
  NAND2_X1 U687 ( .A1(n607), .A2(n606), .ZN(n608) );
  XNOR2_X1 U688 ( .A(KEYINPUT77), .B(n608), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G88), .A2(n627), .ZN(n610) );
  NAND2_X1 U690 ( .A1(G75), .A2(n631), .ZN(n609) );
  AND2_X1 U691 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U692 ( .A1(n612), .A2(n611), .ZN(G303) );
  INV_X1 U693 ( .A(G303), .ZN(G166) );
  NAND2_X1 U694 ( .A1(G49), .A2(n628), .ZN(n615) );
  NAND2_X1 U695 ( .A1(G87), .A2(n613), .ZN(n614) );
  NAND2_X1 U696 ( .A1(n615), .A2(n614), .ZN(n616) );
  NOR2_X1 U697 ( .A1(n635), .A2(n616), .ZN(n618) );
  NAND2_X1 U698 ( .A1(G651), .A2(G74), .ZN(n617) );
  NAND2_X1 U699 ( .A1(n618), .A2(n617), .ZN(G288) );
  XOR2_X1 U700 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n620) );
  NAND2_X1 U701 ( .A1(G73), .A2(n631), .ZN(n619) );
  XNOR2_X1 U702 ( .A(n620), .B(n619), .ZN(n624) );
  NAND2_X1 U703 ( .A1(G86), .A2(n627), .ZN(n622) );
  NAND2_X1 U704 ( .A1(G48), .A2(n628), .ZN(n621) );
  NAND2_X1 U705 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U706 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U707 ( .A1(n635), .A2(G61), .ZN(n625) );
  NAND2_X1 U708 ( .A1(n626), .A2(n625), .ZN(G305) );
  NAND2_X1 U709 ( .A1(G85), .A2(n627), .ZN(n630) );
  NAND2_X1 U710 ( .A1(G47), .A2(n628), .ZN(n629) );
  NAND2_X1 U711 ( .A1(n630), .A2(n629), .ZN(n634) );
  NAND2_X1 U712 ( .A1(n631), .A2(G72), .ZN(n632) );
  XOR2_X1 U713 ( .A(KEYINPUT66), .B(n632), .Z(n633) );
  NOR2_X1 U714 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n635), .A2(G60), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(G290) );
  INV_X1 U717 ( .A(G299), .ZN(n981) );
  XNOR2_X1 U718 ( .A(n981), .B(G166), .ZN(n642) );
  XNOR2_X1 U719 ( .A(KEYINPUT19), .B(G288), .ZN(n638) );
  XNOR2_X1 U720 ( .A(n638), .B(G305), .ZN(n639) );
  XOR2_X1 U721 ( .A(n646), .B(n639), .Z(n640) );
  XNOR2_X1 U722 ( .A(n640), .B(G290), .ZN(n641) );
  XNOR2_X1 U723 ( .A(n642), .B(n641), .ZN(n888) );
  XNOR2_X1 U724 ( .A(n643), .B(n888), .ZN(n644) );
  NAND2_X1 U725 ( .A1(n644), .A2(G868), .ZN(n648) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(n647) );
  NAND2_X1 U727 ( .A1(n648), .A2(n647), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n649) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n649), .Z(n650) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n650), .ZN(n651) );
  XNOR2_X1 U731 ( .A(KEYINPUT21), .B(n651), .ZN(n652) );
  NAND2_X1 U732 ( .A1(n652), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U733 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U734 ( .A1(G220), .A2(G219), .ZN(n653) );
  XOR2_X1 U735 ( .A(KEYINPUT22), .B(n653), .Z(n654) );
  NOR2_X1 U736 ( .A1(G218), .A2(n654), .ZN(n655) );
  XNOR2_X1 U737 ( .A(KEYINPUT78), .B(n655), .ZN(n656) );
  NAND2_X1 U738 ( .A1(n656), .A2(G96), .ZN(n839) );
  NAND2_X1 U739 ( .A1(G2106), .A2(n839), .ZN(n657) );
  XOR2_X1 U740 ( .A(KEYINPUT79), .B(n657), .Z(n662) );
  NAND2_X1 U741 ( .A1(G120), .A2(G69), .ZN(n658) );
  NOR2_X1 U742 ( .A1(G237), .A2(n658), .ZN(n659) );
  XNOR2_X1 U743 ( .A(KEYINPUT80), .B(n659), .ZN(n660) );
  NAND2_X1 U744 ( .A1(n660), .A2(G108), .ZN(n840) );
  NAND2_X1 U745 ( .A1(G567), .A2(n840), .ZN(n661) );
  NAND2_X1 U746 ( .A1(n662), .A2(n661), .ZN(n887) );
  NAND2_X1 U747 ( .A1(G661), .A2(G483), .ZN(n663) );
  NOR2_X1 U748 ( .A1(n887), .A2(n663), .ZN(n838) );
  NAND2_X1 U749 ( .A1(G36), .A2(n838), .ZN(n664) );
  XOR2_X1 U750 ( .A(KEYINPUT81), .B(n664), .Z(G176) );
  NAND2_X1 U751 ( .A1(G138), .A2(n876), .ZN(n666) );
  NAND2_X1 U752 ( .A1(G102), .A2(n878), .ZN(n665) );
  NAND2_X1 U753 ( .A1(n666), .A2(n665), .ZN(n670) );
  NAND2_X1 U754 ( .A1(G126), .A2(n583), .ZN(n668) );
  NAND2_X1 U755 ( .A1(G114), .A2(n873), .ZN(n667) );
  NAND2_X1 U756 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U757 ( .A1(n670), .A2(n669), .ZN(G164) );
  XNOR2_X1 U758 ( .A(G1986), .B(G290), .ZN(n984) );
  NOR2_X1 U759 ( .A1(G164), .A2(G1384), .ZN(n710) );
  INV_X1 U760 ( .A(G40), .ZN(n672) );
  NOR2_X1 U761 ( .A1(n672), .A2(n671), .ZN(n673) );
  AND2_X1 U762 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U763 ( .A1(n676), .A2(n675), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n677), .B(KEYINPUT82), .ZN(n709) );
  NOR2_X1 U765 ( .A1(n710), .A2(n709), .ZN(n678) );
  XNOR2_X1 U766 ( .A(KEYINPUT83), .B(n678), .ZN(n707) );
  INV_X1 U767 ( .A(n707), .ZN(n820) );
  NAND2_X1 U768 ( .A1(n984), .A2(n820), .ZN(n810) );
  XNOR2_X1 U769 ( .A(G2067), .B(KEYINPUT37), .ZN(n818) );
  NAND2_X1 U770 ( .A1(G140), .A2(n876), .ZN(n680) );
  NAND2_X1 U771 ( .A1(G104), .A2(n878), .ZN(n679) );
  NAND2_X1 U772 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U773 ( .A(KEYINPUT34), .B(n681), .ZN(n686) );
  NAND2_X1 U774 ( .A1(G128), .A2(n583), .ZN(n683) );
  NAND2_X1 U775 ( .A1(G116), .A2(n873), .ZN(n682) );
  NAND2_X1 U776 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U777 ( .A(KEYINPUT35), .B(n684), .Z(n685) );
  NOR2_X1 U778 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U779 ( .A(KEYINPUT36), .B(n687), .ZN(n867) );
  NOR2_X1 U780 ( .A1(n818), .A2(n867), .ZN(n953) );
  NAND2_X1 U781 ( .A1(n953), .A2(n820), .ZN(n816) );
  XNOR2_X1 U782 ( .A(KEYINPUT86), .B(G1991), .ZN(n924) );
  NAND2_X1 U783 ( .A1(G119), .A2(n583), .ZN(n689) );
  NAND2_X1 U784 ( .A1(G107), .A2(n873), .ZN(n688) );
  NAND2_X1 U785 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U786 ( .A(KEYINPUT84), .B(n690), .ZN(n695) );
  NAND2_X1 U787 ( .A1(n878), .A2(G95), .ZN(n691) );
  XOR2_X1 U788 ( .A(KEYINPUT85), .B(n691), .Z(n693) );
  NAND2_X1 U789 ( .A1(n876), .A2(G131), .ZN(n692) );
  NAND2_X1 U790 ( .A1(n693), .A2(n692), .ZN(n694) );
  OR2_X1 U791 ( .A1(n695), .A2(n694), .ZN(n866) );
  AND2_X1 U792 ( .A1(n924), .A2(n866), .ZN(n706) );
  NAND2_X1 U793 ( .A1(G141), .A2(n876), .ZN(n696) );
  XNOR2_X1 U794 ( .A(n696), .B(KEYINPUT88), .ZN(n704) );
  NAND2_X1 U795 ( .A1(n878), .A2(G105), .ZN(n697) );
  XNOR2_X1 U796 ( .A(n697), .B(KEYINPUT38), .ZN(n699) );
  NAND2_X1 U797 ( .A1(G129), .A2(n583), .ZN(n698) );
  NAND2_X1 U798 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U799 ( .A1(G117), .A2(n873), .ZN(n700) );
  XNOR2_X1 U800 ( .A(KEYINPUT87), .B(n700), .ZN(n701) );
  NOR2_X1 U801 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n865) );
  AND2_X1 U803 ( .A1(n865), .A2(G1996), .ZN(n705) );
  NOR2_X1 U804 ( .A1(n706), .A2(n705), .ZN(n946) );
  NOR2_X1 U805 ( .A1(n946), .A2(n707), .ZN(n813) );
  INV_X1 U806 ( .A(n813), .ZN(n708) );
  NAND2_X1 U807 ( .A1(n816), .A2(n708), .ZN(n808) );
  XNOR2_X1 U808 ( .A(KEYINPUT89), .B(n709), .ZN(n711) );
  NAND2_X1 U809 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X2 U810 ( .A(n712), .B(KEYINPUT64), .ZN(n742) );
  NOR2_X1 U811 ( .A1(n742), .A2(G2090), .ZN(n714) );
  NAND2_X1 U812 ( .A1(n742), .A2(G8), .ZN(n791) );
  NOR2_X1 U813 ( .A1(G1971), .A2(n791), .ZN(n713) );
  NOR2_X1 U814 ( .A1(n714), .A2(n713), .ZN(n715) );
  NAND2_X1 U815 ( .A1(n715), .A2(G303), .ZN(n716) );
  XNOR2_X1 U816 ( .A(KEYINPUT96), .B(n716), .ZN(n761) );
  NOR2_X1 U817 ( .A1(n742), .A2(G2084), .ZN(n770) );
  NOR2_X1 U818 ( .A1(G1966), .A2(n791), .ZN(n768) );
  NOR2_X1 U819 ( .A1(n770), .A2(n768), .ZN(n717) );
  XNOR2_X1 U820 ( .A(n717), .B(KEYINPUT92), .ZN(n718) );
  NAND2_X1 U821 ( .A1(n718), .A2(G8), .ZN(n721) );
  INV_X1 U822 ( .A(KEYINPUT93), .ZN(n719) );
  NOR2_X1 U823 ( .A1(n722), .A2(G168), .ZN(n728) );
  INV_X1 U824 ( .A(n742), .ZN(n741) );
  NOR2_X1 U825 ( .A1(G1961), .A2(n741), .ZN(n725) );
  XOR2_X1 U826 ( .A(G2078), .B(KEYINPUT25), .Z(n919) );
  NOR2_X1 U827 ( .A1(n742), .A2(n919), .ZN(n723) );
  XNOR2_X1 U828 ( .A(n723), .B(KEYINPUT90), .ZN(n724) );
  NOR2_X1 U829 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U830 ( .A(KEYINPUT91), .B(n726), .ZN(n731) );
  NOR2_X1 U831 ( .A1(G171), .A2(n731), .ZN(n727) );
  NOR2_X1 U832 ( .A1(n728), .A2(n727), .ZN(n730) );
  XNOR2_X1 U833 ( .A(n730), .B(n729), .ZN(n758) );
  NAND2_X1 U834 ( .A1(n731), .A2(G171), .ZN(n756) );
  NAND2_X1 U835 ( .A1(G2072), .A2(n741), .ZN(n732) );
  XNOR2_X1 U836 ( .A(n732), .B(KEYINPUT27), .ZN(n734) );
  INV_X1 U837 ( .A(G1956), .ZN(n998) );
  NOR2_X1 U838 ( .A1(n741), .A2(n998), .ZN(n733) );
  NOR2_X1 U839 ( .A1(n734), .A2(n733), .ZN(n736) );
  NOR2_X1 U840 ( .A1(n981), .A2(n736), .ZN(n735) );
  XOR2_X1 U841 ( .A(n735), .B(KEYINPUT28), .Z(n753) );
  NAND2_X1 U842 ( .A1(n981), .A2(n736), .ZN(n751) );
  AND2_X1 U843 ( .A1(n741), .A2(G1996), .ZN(n737) );
  XOR2_X1 U844 ( .A(n737), .B(KEYINPUT26), .Z(n739) );
  NAND2_X1 U845 ( .A1(n742), .A2(G1341), .ZN(n738) );
  NAND2_X1 U846 ( .A1(n739), .A2(n738), .ZN(n740) );
  NOR2_X1 U847 ( .A1(n992), .A2(n740), .ZN(n746) );
  NAND2_X1 U848 ( .A1(G2067), .A2(n741), .ZN(n744) );
  NAND2_X1 U849 ( .A1(n742), .A2(G1348), .ZN(n743) );
  NAND2_X1 U850 ( .A1(n744), .A2(n743), .ZN(n747) );
  NOR2_X1 U851 ( .A1(n974), .A2(n747), .ZN(n745) );
  OR2_X1 U852 ( .A1(n746), .A2(n745), .ZN(n749) );
  NAND2_X1 U853 ( .A1(n974), .A2(n747), .ZN(n748) );
  NAND2_X1 U854 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U855 ( .A1(n751), .A2(n750), .ZN(n752) );
  NAND2_X1 U856 ( .A1(n753), .A2(n752), .ZN(n754) );
  XOR2_X1 U857 ( .A(KEYINPUT29), .B(n754), .Z(n755) );
  NAND2_X1 U858 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U859 ( .A1(n758), .A2(n757), .ZN(n766) );
  NAND2_X1 U860 ( .A1(G286), .A2(n766), .ZN(n759) );
  XOR2_X1 U861 ( .A(KEYINPUT95), .B(n759), .Z(n760) );
  NAND2_X1 U862 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U863 ( .A1(n762), .A2(G8), .ZN(n765) );
  XOR2_X1 U864 ( .A(KEYINPUT32), .B(KEYINPUT98), .Z(n763) );
  INV_X1 U865 ( .A(n766), .ZN(n767) );
  NOR2_X1 U866 ( .A1(n768), .A2(n767), .ZN(n769) );
  XNOR2_X1 U867 ( .A(n769), .B(KEYINPUT94), .ZN(n772) );
  NAND2_X1 U868 ( .A1(n770), .A2(G8), .ZN(n771) );
  NAND2_X1 U869 ( .A1(n772), .A2(n771), .ZN(n793) );
  XOR2_X1 U870 ( .A(G1981), .B(G305), .Z(n971) );
  NOR2_X1 U871 ( .A1(G1976), .A2(G288), .ZN(n773) );
  XOR2_X1 U872 ( .A(KEYINPUT99), .B(n773), .Z(n796) );
  INV_X1 U873 ( .A(n796), .ZN(n979) );
  NOR2_X1 U874 ( .A1(n791), .A2(n979), .ZN(n774) );
  NAND2_X1 U875 ( .A1(KEYINPUT33), .A2(n774), .ZN(n775) );
  AND2_X1 U876 ( .A1(n971), .A2(n775), .ZN(n788) );
  NAND2_X1 U877 ( .A1(n788), .A2(KEYINPUT33), .ZN(n781) );
  INV_X1 U878 ( .A(n781), .ZN(n776) );
  OR2_X1 U879 ( .A1(n776), .A2(n791), .ZN(n778) );
  AND2_X1 U880 ( .A1(n793), .A2(n778), .ZN(n777) );
  NAND2_X1 U881 ( .A1(n795), .A2(n777), .ZN(n786) );
  INV_X1 U882 ( .A(n778), .ZN(n784) );
  NOR2_X1 U883 ( .A1(G2090), .A2(G303), .ZN(n779) );
  NAND2_X1 U884 ( .A1(G8), .A2(n779), .ZN(n780) );
  XNOR2_X1 U885 ( .A(n780), .B(KEYINPUT100), .ZN(n782) );
  AND2_X1 U886 ( .A1(n782), .A2(n781), .ZN(n783) );
  OR2_X1 U887 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U888 ( .A1(n786), .A2(n785), .ZN(n806) );
  NOR2_X1 U889 ( .A1(G1981), .A2(G305), .ZN(n787) );
  XNOR2_X1 U890 ( .A(KEYINPUT24), .B(n787), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G1976), .A2(G288), .ZN(n980) );
  AND2_X1 U892 ( .A1(n788), .A2(n980), .ZN(n789) );
  NOR2_X1 U893 ( .A1(n798), .A2(n789), .ZN(n790) );
  OR2_X1 U894 ( .A1(n791), .A2(n790), .ZN(n802) );
  INV_X1 U895 ( .A(n802), .ZN(n792) );
  AND2_X1 U896 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U897 ( .A1(n795), .A2(n794), .ZN(n804) );
  NOR2_X1 U898 ( .A1(G1971), .A2(G303), .ZN(n797) );
  NOR2_X1 U899 ( .A1(n797), .A2(n796), .ZN(n800) );
  INV_X1 U900 ( .A(n798), .ZN(n799) );
  AND2_X1 U901 ( .A1(n800), .A2(n799), .ZN(n801) );
  OR2_X1 U902 ( .A1(n802), .A2(n801), .ZN(n803) );
  NAND2_X1 U903 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U904 ( .A1(n806), .A2(n805), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  NAND2_X1 U906 ( .A1(n810), .A2(n809), .ZN(n823) );
  NOR2_X1 U907 ( .A1(G1996), .A2(n865), .ZN(n958) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n811) );
  NOR2_X1 U909 ( .A1(n924), .A2(n866), .ZN(n948) );
  NOR2_X1 U910 ( .A1(n811), .A2(n948), .ZN(n812) );
  NOR2_X1 U911 ( .A1(n813), .A2(n812), .ZN(n814) );
  NOR2_X1 U912 ( .A1(n958), .A2(n814), .ZN(n815) );
  XNOR2_X1 U913 ( .A(n815), .B(KEYINPUT39), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n818), .A2(n867), .ZN(n945) );
  NAND2_X1 U916 ( .A1(n819), .A2(n945), .ZN(n821) );
  NAND2_X1 U917 ( .A1(n821), .A2(n820), .ZN(n822) );
  NAND2_X1 U918 ( .A1(n823), .A2(n822), .ZN(n824) );
  XNOR2_X1 U919 ( .A(KEYINPUT40), .B(n824), .ZN(G329) );
  XOR2_X1 U920 ( .A(G2454), .B(G2435), .Z(n826) );
  XNOR2_X1 U921 ( .A(G2438), .B(G2427), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n826), .B(n825), .ZN(n833) );
  XOR2_X1 U923 ( .A(KEYINPUT101), .B(G2446), .Z(n828) );
  XNOR2_X1 U924 ( .A(G2443), .B(G2430), .ZN(n827) );
  XNOR2_X1 U925 ( .A(n828), .B(n827), .ZN(n829) );
  XOR2_X1 U926 ( .A(n829), .B(G2451), .Z(n831) );
  XNOR2_X1 U927 ( .A(G1341), .B(G1348), .ZN(n830) );
  XNOR2_X1 U928 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n834), .A2(G14), .ZN(n913) );
  XOR2_X1 U931 ( .A(KEYINPUT102), .B(n913), .Z(G401) );
  NAND2_X1 U932 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U934 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G188) );
  XNOR2_X1 U937 ( .A(G108), .B(KEYINPUT113), .ZN(G238) );
  INV_X1 U939 ( .A(G120), .ZN(G236) );
  INV_X1 U940 ( .A(G96), .ZN(G221) );
  INV_X1 U941 ( .A(G69), .ZN(G235) );
  NOR2_X1 U942 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U943 ( .A(G325), .ZN(G261) );
  NAND2_X1 U944 ( .A1(n583), .A2(G124), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n841), .B(KEYINPUT44), .ZN(n843) );
  NAND2_X1 U946 ( .A1(G112), .A2(n873), .ZN(n842) );
  NAND2_X1 U947 ( .A1(n843), .A2(n842), .ZN(n847) );
  NAND2_X1 U948 ( .A1(G136), .A2(n876), .ZN(n845) );
  NAND2_X1 U949 ( .A1(G100), .A2(n878), .ZN(n844) );
  NAND2_X1 U950 ( .A1(n845), .A2(n844), .ZN(n846) );
  NOR2_X1 U951 ( .A1(n847), .A2(n846), .ZN(G162) );
  XNOR2_X1 U952 ( .A(KEYINPUT47), .B(KEYINPUT107), .ZN(n851) );
  NAND2_X1 U953 ( .A1(G127), .A2(n583), .ZN(n849) );
  NAND2_X1 U954 ( .A1(G115), .A2(n873), .ZN(n848) );
  NAND2_X1 U955 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U956 ( .A(n851), .B(n850), .ZN(n856) );
  NAND2_X1 U957 ( .A1(n878), .A2(G103), .ZN(n852) );
  XNOR2_X1 U958 ( .A(n852), .B(KEYINPUT106), .ZN(n854) );
  NAND2_X1 U959 ( .A1(G139), .A2(n876), .ZN(n853) );
  NAND2_X1 U960 ( .A1(n854), .A2(n853), .ZN(n855) );
  NOR2_X1 U961 ( .A1(n856), .A2(n855), .ZN(n940) );
  XNOR2_X1 U962 ( .A(G162), .B(n940), .ZN(n863) );
  XOR2_X1 U963 ( .A(KEYINPUT111), .B(KEYINPUT109), .Z(n858) );
  XNOR2_X1 U964 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n857) );
  XNOR2_X1 U965 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U966 ( .A(n859), .B(KEYINPUT108), .Z(n861) );
  XNOR2_X1 U967 ( .A(KEYINPUT110), .B(KEYINPUT112), .ZN(n860) );
  XNOR2_X1 U968 ( .A(n861), .B(n860), .ZN(n862) );
  XNOR2_X1 U969 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U970 ( .A(n865), .B(n864), .Z(n869) );
  XOR2_X1 U971 ( .A(n867), .B(n866), .Z(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XOR2_X1 U973 ( .A(n870), .B(n947), .Z(n872) );
  XNOR2_X1 U974 ( .A(G164), .B(G160), .ZN(n871) );
  XNOR2_X1 U975 ( .A(n872), .B(n871), .ZN(n885) );
  NAND2_X1 U976 ( .A1(G130), .A2(n583), .ZN(n875) );
  NAND2_X1 U977 ( .A1(G118), .A2(n873), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n883) );
  NAND2_X1 U979 ( .A1(n876), .A2(G142), .ZN(n877) );
  XOR2_X1 U980 ( .A(KEYINPUT105), .B(n877), .Z(n880) );
  NAND2_X1 U981 ( .A1(n878), .A2(G106), .ZN(n879) );
  NAND2_X1 U982 ( .A1(n880), .A2(n879), .ZN(n881) );
  XOR2_X1 U983 ( .A(n881), .B(KEYINPUT45), .Z(n882) );
  NOR2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XOR2_X1 U985 ( .A(n885), .B(n884), .Z(n886) );
  NOR2_X1 U986 ( .A1(G37), .A2(n886), .ZN(G395) );
  XNOR2_X1 U987 ( .A(KEYINPUT103), .B(n887), .ZN(G319) );
  XNOR2_X1 U988 ( .A(G171), .B(n974), .ZN(n889) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n891) );
  XNOR2_X1 U990 ( .A(n992), .B(G286), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  NOR2_X1 U992 ( .A1(G37), .A2(n892), .ZN(G397) );
  XOR2_X1 U993 ( .A(G2096), .B(KEYINPUT43), .Z(n894) );
  XNOR2_X1 U994 ( .A(G2072), .B(G2678), .ZN(n893) );
  XNOR2_X1 U995 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(n895), .B(KEYINPUT42), .Z(n897) );
  XNOR2_X1 U997 ( .A(G2067), .B(G2090), .ZN(n896) );
  XNOR2_X1 U998 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U999 ( .A(KEYINPUT104), .B(G2100), .Z(n899) );
  XNOR2_X1 U1000 ( .A(G2078), .B(G2084), .ZN(n898) );
  XNOR2_X1 U1001 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U1002 ( .A(n901), .B(n900), .ZN(G227) );
  XOR2_X1 U1003 ( .A(G1986), .B(G1976), .Z(n903) );
  XNOR2_X1 U1004 ( .A(G1956), .B(G1971), .ZN(n902) );
  XNOR2_X1 U1005 ( .A(n903), .B(n902), .ZN(n904) );
  XOR2_X1 U1006 ( .A(n904), .B(G2474), .Z(n906) );
  XNOR2_X1 U1007 ( .A(G1996), .B(G1991), .ZN(n905) );
  XNOR2_X1 U1008 ( .A(n906), .B(n905), .ZN(n910) );
  XOR2_X1 U1009 ( .A(KEYINPUT41), .B(G1981), .Z(n908) );
  XNOR2_X1 U1010 ( .A(G1961), .B(G1966), .ZN(n907) );
  XNOR2_X1 U1011 ( .A(n908), .B(n907), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n910), .B(n909), .ZN(G229) );
  NOR2_X1 U1013 ( .A1(G227), .A2(G229), .ZN(n911) );
  XOR2_X1 U1014 ( .A(KEYINPUT49), .B(n911), .Z(n912) );
  NAND2_X1 U1015 ( .A1(n913), .A2(n912), .ZN(n914) );
  NOR2_X1 U1016 ( .A1(G397), .A2(n914), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(G319), .A2(n915), .ZN(n916) );
  NOR2_X1 U1018 ( .A1(G395), .A2(n916), .ZN(G308) );
  INV_X1 U1019 ( .A(G308), .ZN(G225) );
  XOR2_X1 U1020 ( .A(G2090), .B(G35), .Z(n932) );
  XNOR2_X1 U1021 ( .A(G1996), .B(G32), .ZN(n918) );
  XNOR2_X1 U1022 ( .A(G2067), .B(G26), .ZN(n917) );
  NOR2_X1 U1023 ( .A1(n918), .A2(n917), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n919), .B(G27), .ZN(n921) );
  XNOR2_X1 U1025 ( .A(G2072), .B(G33), .ZN(n920) );
  NOR2_X1 U1026 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1027 ( .A1(n923), .A2(n922), .ZN(n928) );
  XOR2_X1 U1028 ( .A(n924), .B(G25), .Z(n925) );
  NAND2_X1 U1029 ( .A1(n925), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1030 ( .A(n926), .B(KEYINPUT118), .ZN(n927) );
  NOR2_X1 U1031 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1032 ( .A(n929), .B(KEYINPUT119), .ZN(n930) );
  XNOR2_X1 U1033 ( .A(n930), .B(KEYINPUT53), .ZN(n931) );
  NAND2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(G34), .B(G2084), .ZN(n933) );
  XNOR2_X1 U1036 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NOR2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1038 ( .A(KEYINPUT55), .B(n936), .Z(n937) );
  XNOR2_X1 U1039 ( .A(KEYINPUT120), .B(n937), .ZN(n938) );
  NOR2_X1 U1040 ( .A1(G29), .A2(n938), .ZN(n939) );
  XNOR2_X1 U1041 ( .A(n939), .B(KEYINPUT121), .ZN(n969) );
  XNOR2_X1 U1042 ( .A(KEYINPUT52), .B(KEYINPUT117), .ZN(n965) );
  XNOR2_X1 U1043 ( .A(G164), .B(G2078), .ZN(n943) );
  XNOR2_X1 U1044 ( .A(G2072), .B(n940), .ZN(n941) );
  XNOR2_X1 U1045 ( .A(n941), .B(KEYINPUT116), .ZN(n942) );
  NAND2_X1 U1046 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1047 ( .A(n944), .B(KEYINPUT50), .ZN(n963) );
  NAND2_X1 U1048 ( .A1(n946), .A2(n945), .ZN(n956) );
  XNOR2_X1 U1049 ( .A(G160), .B(G2084), .ZN(n950) );
  NOR2_X1 U1050 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1051 ( .A1(n950), .A2(n949), .ZN(n951) );
  XNOR2_X1 U1052 ( .A(KEYINPUT114), .B(n951), .ZN(n952) );
  NOR2_X1 U1053 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1054 ( .A(KEYINPUT115), .B(n954), .ZN(n955) );
  NOR2_X1 U1055 ( .A1(n956), .A2(n955), .ZN(n961) );
  XOR2_X1 U1056 ( .A(G2090), .B(G162), .Z(n957) );
  NOR2_X1 U1057 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1058 ( .A(KEYINPUT51), .B(n959), .Z(n960) );
  NAND2_X1 U1059 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1060 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1061 ( .A(n965), .B(n964), .ZN(n966) );
  OR2_X1 U1062 ( .A1(KEYINPUT55), .A2(n966), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(G29), .A2(n967), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n1026) );
  INV_X1 U1065 ( .A(G16), .ZN(n1021) );
  XOR2_X1 U1066 ( .A(KEYINPUT56), .B(KEYINPUT122), .Z(n970) );
  XNOR2_X1 U1067 ( .A(n1021), .B(n970), .ZN(n996) );
  XNOR2_X1 U1068 ( .A(G168), .B(G1966), .ZN(n972) );
  NAND2_X1 U1069 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n973), .B(KEYINPUT57), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(G301), .B(G1961), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(n974), .B(G1348), .ZN(n975) );
  NOR2_X1 U1073 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1074 ( .A1(n978), .A2(n977), .ZN(n991) );
  NAND2_X1 U1075 ( .A1(n980), .A2(n979), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(n998), .B(n981), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(n982), .B(KEYINPUT123), .ZN(n986) );
  XNOR2_X1 U1078 ( .A(G1971), .B(G303), .ZN(n983) );
  NOR2_X1 U1079 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1082 ( .A(KEYINPUT124), .B(n989), .Z(n990) );
  NOR2_X1 U1083 ( .A1(n991), .A2(n990), .ZN(n994) );
  XOR2_X1 U1084 ( .A(G1341), .B(n992), .Z(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n1023) );
  XNOR2_X1 U1087 ( .A(KEYINPUT125), .B(G1966), .ZN(n997) );
  XNOR2_X1 U1088 ( .A(n997), .B(G21), .ZN(n1010) );
  XNOR2_X1 U1089 ( .A(G20), .B(n998), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1341), .B(G19), .ZN(n1000) );
  XNOR2_X1 U1091 ( .A(G6), .B(G1981), .ZN(n999) );
  NOR2_X1 U1092 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1005) );
  XOR2_X1 U1094 ( .A(KEYINPUT59), .B(G1348), .Z(n1003) );
  XNOR2_X1 U1095 ( .A(G4), .B(n1003), .ZN(n1004) );
  NOR2_X1 U1096 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1097 ( .A(KEYINPUT60), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1098 ( .A(G1961), .B(G5), .ZN(n1007) );
  NOR2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1012) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1011) );
  NOR2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1013) );
  NAND2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1015), .ZN(n1016) );
  NOR2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1108 ( .A(n1018), .B(KEYINPUT61), .ZN(n1019) );
  XNOR2_X1 U1109 ( .A(n1019), .B(KEYINPUT126), .ZN(n1020) );
  NAND2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1111 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1024), .Z(n1025) );
  NOR2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1114 ( .A1(n1027), .A2(G11), .ZN(n1028) );
  XOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1028), .Z(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

