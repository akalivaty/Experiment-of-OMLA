//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:40 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1269, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(G13), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G68), .A2(G238), .B1(G116), .B2(G270), .ZN(new_n217));
  INV_X1    g0017(.A(G226), .ZN(new_n218));
  OAI21_X1  g0018(.A(new_n217), .B1(new_n202), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g0019(.A(KEYINPUT64), .B(G77), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g0021(.A(new_n219), .B1(G244), .B2(new_n221), .ZN(new_n222));
  INV_X1    g0022(.A(KEYINPUT65), .ZN(new_n223));
  AOI22_X1  g0023(.A1(new_n222), .A2(new_n223), .B1(G107), .B2(G264), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n224), .B1(new_n223), .B2(new_n222), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(G87), .B2(G250), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G97), .A2(G257), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n211), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  XOR2_X1   g0030(.A(new_n230), .B(KEYINPUT1), .Z(new_n231));
  NAND2_X1  g0031(.A1(G1), .A2(G13), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n232), .A2(new_n210), .ZN(new_n233));
  INV_X1    g0033(.A(new_n201), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n234), .A2(G50), .ZN(new_n235));
  INV_X1    g0035(.A(new_n235), .ZN(new_n236));
  AOI211_X1 g0036(.A(new_n216), .B(new_n231), .C1(new_n233), .C2(new_n236), .ZN(G361));
  XOR2_X1   g0037(.A(G250), .B(G257), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G270), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT66), .B(G264), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(new_n226), .ZN(new_n243));
  XOR2_X1   g0043(.A(KEYINPUT2), .B(G226), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n241), .B(new_n245), .ZN(G358));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  INV_X1    g0047(.A(G116), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(KEYINPUT67), .B(G107), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G50), .B(G58), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XOR2_X1   g0054(.A(new_n251), .B(new_n254), .Z(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n232), .ZN(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G77), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NOR2_X1   g0062(.A1(G20), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n264), .A2(new_n202), .B1(new_n210), .B2(G68), .ZN(new_n265));
  OAI21_X1  g0065(.A(new_n257), .B1(new_n262), .B2(new_n265), .ZN(new_n266));
  XOR2_X1   g0066(.A(KEYINPUT77), .B(KEYINPUT11), .Z(new_n267));
  XNOR2_X1  g0067(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT12), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(new_n271), .B2(G68), .ZN(new_n272));
  INV_X1    g0072(.A(new_n271), .ZN(new_n273));
  INV_X1    g0073(.A(G68), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n273), .A2(KEYINPUT12), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n257), .B1(new_n209), .B2(G20), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n272), .B(new_n275), .C1(new_n277), .C2(new_n274), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n226), .A2(G1698), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  OAI221_X1 g0084(.A(new_n282), .B1(G226), .B2(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT75), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G97), .ZN(new_n287));
  AND3_X1   g0087(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(new_n285), .B2(new_n287), .ZN(new_n289));
  AND2_X1   g0089(.A1(G1), .A2(G13), .ZN(new_n290));
  NAND2_X1  g0090(.A1(G33), .A2(G41), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NOR3_X1   g0092(.A1(new_n288), .A2(new_n289), .A3(new_n292), .ZN(new_n293));
  AND2_X1   g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  OAI21_X1  g0094(.A(KEYINPUT68), .B1(new_n294), .B2(new_n232), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT68), .ZN(new_n296));
  NAND3_X1  g0096(.A1(new_n290), .A2(new_n296), .A3(new_n291), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G41), .ZN(new_n299));
  INV_X1    g0099(.A(G45), .ZN(new_n300));
  AOI21_X1  g0100(.A(G1), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n298), .A2(G274), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n301), .B1(new_n295), .B2(new_n297), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(G238), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n302), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(KEYINPUT13), .B1(new_n293), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n289), .ZN(new_n308));
  INV_X1    g0108(.A(new_n292), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n285), .A2(new_n286), .A3(new_n287), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n308), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  INV_X1    g0112(.A(G274), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n313), .B1(new_n295), .B2(new_n297), .ZN(new_n314));
  AOI22_X1  g0114(.A1(G238), .A2(new_n303), .B1(new_n314), .B2(new_n301), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n311), .A2(new_n312), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n281), .B1(new_n307), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT14), .ZN(new_n318));
  XNOR2_X1  g0118(.A(new_n317), .B(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(G179), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n307), .A2(new_n316), .A3(KEYINPUT76), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT76), .ZN(new_n322));
  OAI211_X1 g0122(.A(new_n322), .B(KEYINPUT13), .C1(new_n293), .C2(new_n306), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n320), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n280), .B1(new_n319), .B2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT78), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n321), .A2(new_n323), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n280), .B1(new_n327), .B2(G190), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n307), .A2(new_n316), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n329), .A2(G200), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n325), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  XOR2_X1   g0132(.A(KEYINPUT8), .B(G58), .Z(new_n333));
  AOI22_X1  g0133(.A1(new_n221), .A2(G20), .B1(new_n333), .B2(new_n263), .ZN(new_n334));
  XOR2_X1   g0134(.A(KEYINPUT15), .B(G87), .Z(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n334), .B1(new_n260), .B2(new_n336), .ZN(new_n337));
  AOI22_X1  g0137(.A1(new_n337), .A2(new_n257), .B1(new_n220), .B2(new_n273), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n276), .A2(G77), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  XNOR2_X1  g0141(.A(KEYINPUT3), .B(G33), .ZN(new_n342));
  INV_X1    g0142(.A(G1698), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n342), .A2(G232), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n342), .A2(G238), .A3(G1698), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n283), .A2(new_n284), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G107), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n309), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n303), .A2(G244), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(new_n302), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT71), .ZN(new_n352));
  XOR2_X1   g0152(.A(KEYINPUT73), .B(G200), .Z(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT71), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n349), .A2(new_n355), .A3(new_n302), .A4(new_n350), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n354), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n352), .A2(new_n356), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT72), .B1(new_n358), .B2(G190), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT72), .ZN(new_n360));
  INV_X1    g0160(.A(G190), .ZN(new_n361));
  AOI211_X1 g0161(.A(new_n360), .B(new_n361), .C1(new_n352), .C2(new_n356), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n341), .B(new_n357), .C1(new_n359), .C2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT16), .ZN(new_n364));
  OR2_X1    g0164(.A1(KEYINPUT3), .A2(G33), .ZN(new_n365));
  NAND2_X1  g0165(.A1(KEYINPUT3), .A2(G33), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n210), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT7), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n365), .A2(KEYINPUT7), .A3(new_n210), .A4(new_n366), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n274), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n225), .A2(new_n274), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n372), .B2(new_n201), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n263), .A2(G159), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n364), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT80), .ZN(new_n377));
  INV_X1    g0177(.A(new_n375), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT79), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n369), .A2(new_n379), .A3(new_n370), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g0181(.A(G68), .B1(new_n369), .B2(new_n379), .ZN(new_n382));
  OAI211_X1 g0182(.A(KEYINPUT16), .B(new_n378), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  OAI211_X1 g0184(.A(new_n384), .B(new_n364), .C1(new_n371), .C2(new_n375), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n377), .A2(new_n383), .A3(new_n257), .A4(new_n385), .ZN(new_n386));
  OR2_X1    g0186(.A1(G223), .A2(G1698), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n218), .A2(G1698), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n388), .C1(new_n283), .C2(new_n284), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G33), .A2(G87), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(new_n309), .ZN(new_n392));
  INV_X1    g0192(.A(new_n301), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n298), .A2(G232), .A3(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n392), .A2(new_n302), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(KEYINPUT82), .B1(new_n395), .B2(G190), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n301), .A2(new_n314), .B1(new_n391), .B2(new_n309), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT82), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n397), .A2(new_n398), .A3(new_n361), .A4(new_n394), .ZN(new_n399));
  INV_X1    g0199(.A(G200), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n396), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT70), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(G58), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT8), .ZN(new_n405));
  XNOR2_X1  g0205(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n277), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n407), .B1(new_n273), .B2(new_n406), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n386), .A2(new_n402), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(KEYINPUT83), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n409), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g0212(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NAND4_X1  g0214(.A1(new_n386), .A2(new_n402), .A3(new_n408), .A4(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n386), .A2(new_n408), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n397), .A2(G179), .A3(new_n394), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n395), .A2(G169), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT18), .B1(new_n417), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT81), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  AOI221_X4 g0224(.A(new_n424), .B1(new_n419), .B2(new_n418), .C1(new_n386), .C2(new_n408), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n422), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n417), .A2(KEYINPUT18), .A3(new_n421), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT81), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n416), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n332), .A2(new_n363), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n203), .A2(G20), .ZN(new_n431));
  INV_X1    g0231(.A(G150), .ZN(new_n432));
  OAI221_X1 g0232(.A(new_n431), .B1(new_n432), .B2(new_n264), .C1(new_n406), .C2(new_n260), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n257), .B1(new_n202), .B2(new_n273), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(new_n202), .B2(new_n277), .ZN(new_n435));
  INV_X1    g0235(.A(KEYINPUT9), .ZN(new_n436));
  OR2_X1    g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n436), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT10), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n346), .A2(new_n220), .ZN(new_n441));
  NOR2_X1   g0241(.A1(G222), .A2(G1698), .ZN(new_n442));
  XOR2_X1   g0242(.A(KEYINPUT69), .B(G223), .Z(new_n443));
  AOI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(G1698), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n309), .B(new_n441), .C1(new_n444), .C2(new_n346), .ZN(new_n445));
  OAI211_X1 g0245(.A(new_n445), .B(new_n302), .C1(new_n218), .C2(new_n304), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n446), .A2(new_n361), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n446), .A2(new_n354), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT74), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n439), .A2(new_n440), .A3(new_n447), .A4(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(new_n447), .A3(new_n438), .ZN(new_n451));
  INV_X1    g0251(.A(new_n449), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT10), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  OR2_X1    g0254(.A1(new_n446), .A2(G179), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n446), .A2(new_n281), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n455), .A2(new_n435), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n358), .A2(new_n320), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n458), .B(new_n340), .C1(G169), .C2(new_n358), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n326), .B1(new_n325), .B2(new_n331), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT88), .ZN(new_n462));
  OAI211_X1 g0262(.A(G244), .B(new_n343), .C1(new_n283), .C2(new_n284), .ZN(new_n463));
  INV_X1    g0263(.A(KEYINPUT4), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n342), .A2(KEYINPUT4), .A3(G244), .A4(new_n343), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G283), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n342), .A2(G250), .A3(G1698), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n465), .A2(new_n466), .A3(new_n467), .A4(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n309), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT87), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n209), .B(G45), .C1(new_n299), .C2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT86), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n300), .A2(G1), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT5), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(KEYINPUT86), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n471), .B1(new_n474), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n299), .A2(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n472), .A2(new_n473), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n475), .A2(KEYINPUT86), .A3(new_n477), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(KEYINPUT87), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n479), .A2(new_n314), .A3(new_n480), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(new_n482), .A3(new_n480), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G257), .A3(new_n298), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n470), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n400), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n470), .A2(new_n484), .A3(new_n361), .A4(new_n486), .ZN(new_n489));
  AND2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n271), .A2(G97), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n209), .A2(G33), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n271), .A2(new_n493), .A3(new_n232), .A4(new_n256), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(new_n205), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n369), .A2(new_n370), .ZN(new_n497));
  AOI21_X1  g0297(.A(KEYINPUT85), .B1(new_n497), .B2(G107), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT85), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n499), .B(new_n206), .C1(new_n369), .C2(new_n370), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n263), .A2(G77), .ZN(new_n501));
  NAND2_X1  g0301(.A1(KEYINPUT6), .A2(G97), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT84), .B1(new_n502), .B2(G107), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT84), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n504), .A2(new_n206), .A3(KEYINPUT6), .A4(G97), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G97), .A2(G107), .ZN(new_n507));
  AOI21_X1  g0307(.A(KEYINPUT6), .B1(new_n207), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n501), .B1(new_n509), .B2(new_n210), .ZN(new_n510));
  NOR3_X1   g0310(.A1(new_n498), .A2(new_n500), .A3(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n257), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n492), .B(new_n496), .C1(new_n511), .C2(new_n512), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n462), .B1(new_n490), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT7), .B1(new_n346), .B2(new_n210), .ZN(new_n515));
  NOR4_X1   g0315(.A1(new_n283), .A2(new_n284), .A3(new_n368), .A4(G20), .ZN(new_n516));
  OAI21_X1  g0316(.A(G107), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n499), .ZN(new_n518));
  INV_X1    g0318(.A(new_n507), .ZN(new_n519));
  NOR2_X1   g0319(.A1(G97), .A2(G107), .ZN(new_n520));
  NOR2_X1   g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(new_n503), .B(new_n505), .C1(new_n521), .C2(KEYINPUT6), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(G20), .B1(G77), .B2(new_n263), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n497), .A2(KEYINPUT85), .A3(G107), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n491), .B(new_n495), .C1(new_n525), .C2(new_n257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n488), .A2(new_n489), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT88), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n491), .B1(new_n525), .B2(new_n257), .ZN(new_n529));
  AOI22_X1  g0329(.A1(new_n529), .A2(new_n496), .B1(new_n281), .B2(new_n487), .ZN(new_n530));
  INV_X1    g0330(.A(new_n487), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n320), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n514), .A2(new_n528), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n273), .A2(KEYINPUT25), .A3(new_n206), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(KEYINPUT25), .B1(new_n273), .B2(new_n206), .ZN(new_n536));
  OAI22_X1  g0336(.A1(new_n535), .A2(new_n536), .B1(new_n206), .B2(new_n494), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT94), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n210), .B(G87), .C1(new_n283), .C2(new_n284), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND4_X1  g0342(.A1(new_n342), .A2(KEYINPUT22), .A3(new_n210), .A4(G87), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT23), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n210), .B2(G107), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n546));
  AOI22_X1  g0346(.A1(new_n545), .A2(new_n546), .B1(new_n259), .B2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT24), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT24), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n542), .A2(new_n543), .A3(new_n550), .A4(new_n547), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(new_n539), .B1(new_n552), .B2(new_n257), .ZN(new_n553));
  AOI211_X1 g0353(.A(KEYINPUT94), .B(new_n512), .C1(new_n549), .C2(new_n551), .ZN(new_n554));
  OAI21_X1  g0354(.A(new_n538), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI211_X1 g0355(.A(G257), .B(G1698), .C1(new_n283), .C2(new_n284), .ZN(new_n556));
  OAI211_X1 g0356(.A(G250), .B(new_n343), .C1(new_n283), .C2(new_n284), .ZN(new_n557));
  NAND2_X1  g0357(.A1(G33), .A2(G294), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n309), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n485), .A2(G264), .A3(new_n298), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n484), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n281), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n483), .A2(new_n314), .A3(new_n480), .ZN(new_n564));
  AOI21_X1  g0364(.A(KEYINPUT87), .B1(new_n481), .B2(new_n482), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n561), .A2(new_n560), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n320), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n555), .A2(new_n563), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n342), .A2(G257), .A3(new_n343), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n342), .A2(G264), .A3(G1698), .ZN(new_n572));
  INV_X1    g0372(.A(G303), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n342), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n309), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n485), .A2(G270), .A3(new_n298), .ZN(new_n576));
  AND3_X1   g0376(.A1(new_n575), .A2(new_n484), .A3(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n467), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT90), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(G20), .B1(new_n258), .B2(G97), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n581), .A2(KEYINPUT90), .A3(new_n467), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT91), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT20), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n256), .A2(new_n232), .B1(G20), .B2(new_n248), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n580), .A2(new_n582), .A3(new_n585), .A4(new_n586), .ZN(new_n587));
  NOR2_X1   g0387(.A1(new_n583), .A2(new_n584), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n587), .A2(new_n588), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n273), .A2(new_n248), .ZN(new_n591));
  INV_X1    g0391(.A(new_n494), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G116), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n589), .A2(new_n590), .A3(new_n591), .A4(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n577), .A2(new_n594), .A3(G179), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT92), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n575), .A2(new_n484), .A3(G179), .A4(new_n576), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT92), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n594), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n575), .A2(new_n484), .A3(new_n576), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n594), .A2(G169), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(KEYINPUT21), .ZN(new_n604));
  INV_X1    g0404(.A(KEYINPUT21), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n594), .A2(new_n602), .A3(new_n605), .A4(G169), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n570), .A2(new_n601), .A3(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT93), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n594), .B1(G200), .B2(new_n602), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n577), .A2(G190), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n610), .A2(new_n609), .A3(new_n611), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n305), .A2(new_n343), .ZN(new_n616));
  INV_X1    g0416(.A(G244), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G1698), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n616), .B(new_n618), .C1(new_n283), .C2(new_n284), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G33), .A2(G116), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n621), .A2(new_n309), .ZN(new_n622));
  AOI21_X1  g0422(.A(G250), .B1(new_n209), .B2(G45), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n300), .A2(G1), .A3(G274), .ZN(new_n625));
  INV_X1    g0425(.A(new_n625), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n298), .A2(new_n624), .A3(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(G169), .B1(new_n622), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n335), .A2(new_n271), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT19), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n210), .B1(new_n287), .B2(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G87), .ZN(new_n632));
  AND4_X1   g0432(.A1(KEYINPUT89), .A2(new_n632), .A3(new_n205), .A4(new_n206), .ZN(new_n633));
  AOI21_X1  g0433(.A(KEYINPUT89), .B1(new_n520), .B2(new_n632), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n342), .A2(new_n210), .A3(G68), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n630), .B1(new_n260), .B2(new_n205), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n629), .B1(new_n638), .B2(new_n257), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n592), .A2(new_n335), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n628), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  AOI211_X1 g0441(.A(new_n623), .B(new_n625), .C1(new_n295), .C2(new_n297), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n292), .B1(new_n619), .B2(new_n620), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n320), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  NOR3_X1   g0446(.A1(new_n642), .A2(new_n643), .A3(new_n361), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n353), .B1(new_n622), .B2(new_n627), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n494), .A2(new_n632), .ZN(new_n650));
  AOI211_X1 g0450(.A(new_n629), .B(new_n650), .C1(new_n638), .C2(new_n257), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n552), .A2(new_n257), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(KEYINPUT94), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n552), .A2(new_n539), .A3(new_n257), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n537), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n400), .B1(new_n566), .B2(new_n567), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(KEYINPUT95), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n568), .A2(new_n361), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT95), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n562), .A2(new_n661), .A3(new_n400), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n659), .A2(new_n660), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n653), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n533), .A2(new_n608), .A3(new_n615), .A4(new_n664), .ZN(new_n665));
  NOR4_X1   g0465(.A1(new_n430), .A2(new_n460), .A3(new_n461), .A4(new_n665), .ZN(G372));
  INV_X1    g0466(.A(new_n457), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT96), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n318), .B1(new_n329), .B2(G169), .ZN(new_n669));
  AOI211_X1 g0469(.A(KEYINPUT14), .B(new_n281), .C1(new_n307), .C2(new_n316), .ZN(new_n670));
  NOR3_X1   g0470(.A1(new_n324), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(new_n279), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n459), .B1(new_n328), .B2(new_n330), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n668), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n328), .A2(new_n330), .ZN(new_n675));
  OAI211_X1 g0475(.A(new_n325), .B(KEYINPUT96), .C1(new_n675), .C2(new_n459), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n412), .A2(new_n415), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n417), .A2(new_n421), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n424), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n427), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n678), .A2(KEYINPUT97), .A3(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n454), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT97), .B1(new_n678), .B2(new_n681), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n667), .B1(new_n683), .B2(new_n685), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n430), .A2(new_n460), .A3(new_n461), .ZN(new_n687));
  INV_X1    g0487(.A(new_n646), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n641), .A2(new_n645), .B1(new_n649), .B2(new_n651), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n487), .A2(new_n281), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(new_n513), .A3(new_n690), .A4(new_n532), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT26), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n530), .A2(KEYINPUT26), .A3(new_n689), .A4(new_n532), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n688), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n530), .A2(new_n532), .ZN(new_n696));
  AOI21_X1  g0496(.A(KEYINPUT88), .B1(new_n526), .B2(new_n527), .ZN(new_n697));
  AND3_X1   g0497(.A1(new_n526), .A2(KEYINPUT88), .A3(new_n527), .ZN(new_n698));
  OAI211_X1 g0498(.A(new_n664), .B(new_n696), .C1(new_n697), .C2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n695), .B1(new_n699), .B2(new_n608), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n687), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n686), .A2(new_n701), .ZN(G369));
  NAND2_X1  g0502(.A1(new_n657), .A2(new_n663), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n212), .A2(G20), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(new_n209), .ZN(new_n705));
  OR2_X1    g0505(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(KEYINPUT27), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n706), .A2(G213), .A3(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(G343), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n555), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n703), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n570), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n570), .B2(new_n710), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND3_X1   g0515(.A1(new_n610), .A2(new_n609), .A3(new_n611), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n601), .B(new_n607), .C1(new_n716), .C2(new_n612), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n594), .A2(new_n710), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n601), .A2(new_n607), .A3(new_n718), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n720), .A2(G330), .A3(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(KEYINPUT98), .ZN(new_n724));
  INV_X1    g0524(.A(KEYINPUT98), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n721), .B1(new_n719), .B2(new_n717), .ZN(new_n726));
  AOI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(G330), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n715), .B1(new_n724), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n570), .A2(new_n710), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n710), .B1(new_n601), .B2(new_n607), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n729), .B1(new_n713), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n731), .ZN(G399));
  NOR2_X1   g0532(.A1(new_n633), .A2(new_n634), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n248), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n213), .A2(G41), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n735), .A2(G1), .A3(new_n737), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n738), .B1(new_n235), .B2(new_n737), .ZN(new_n739));
  XNOR2_X1  g0539(.A(new_n739), .B(KEYINPUT28), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n567), .B1(new_n597), .B2(KEYINPUT99), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n531), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n644), .B1(new_n597), .B2(KEYINPUT99), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n744), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n531), .A4(new_n742), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n487), .A2(new_n602), .A3(new_n562), .ZN(new_n748));
  OR3_X1    g0548(.A1(new_n748), .A2(G179), .A3(new_n644), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(new_n710), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n696), .B1(new_n698), .B2(new_n697), .ZN(new_n753));
  INV_X1    g0553(.A(new_n664), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n710), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n755), .A2(new_n615), .A3(new_n608), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n752), .B1(new_n757), .B2(KEYINPUT31), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n710), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(G330), .B1(new_n758), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n570), .A2(new_n601), .A3(new_n607), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n533), .A2(new_n664), .A3(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n710), .B1(new_n763), .B2(new_n695), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT29), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT29), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  AND2_X1   g0567(.A1(new_n761), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n740), .B1(new_n768), .B2(G1), .ZN(G364));
  NAND2_X1  g0569(.A1(new_n704), .A2(G45), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n737), .A2(G1), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  INV_X1    g0572(.A(new_n726), .ZN(new_n773));
  INV_X1    g0573(.A(G330), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(new_n773), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g0575(.A1(new_n726), .A2(new_n725), .A3(G330), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n723), .A2(KEYINPUT98), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n232), .B1(G20), .B2(new_n281), .ZN(new_n779));
  XOR2_X1   g0579(.A(new_n779), .B(KEYINPUT101), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n210), .A2(G179), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n354), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n361), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n342), .B1(new_n783), .B2(G303), .ZN(new_n784));
  XOR2_X1   g0584(.A(new_n784), .B(KEYINPUT103), .Z(new_n785));
  INV_X1    g0585(.A(G283), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n782), .A2(G190), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n785), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(G20), .A2(G179), .ZN(new_n790));
  XOR2_X1   g0590(.A(new_n790), .B(KEYINPUT102), .Z(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G190), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(G200), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n791), .A2(new_n361), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n400), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G322), .A2(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT104), .Z(new_n798));
  NAND3_X1  g0598(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G326), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n791), .A2(new_n361), .A3(new_n400), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n781), .A2(new_n361), .A3(new_n400), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  AOI22_X1  g0605(.A1(new_n803), .A2(G311), .B1(G329), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n798), .A2(new_n801), .A3(new_n806), .ZN(new_n807));
  NOR3_X1   g0607(.A1(new_n361), .A2(G179), .A3(G200), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n210), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g0610(.A(new_n789), .B(new_n807), .C1(G294), .C2(new_n810), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n346), .B1(new_n803), .B2(new_n221), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT32), .ZN(new_n813));
  INV_X1    g0613(.A(G159), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n804), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n783), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n812), .B1(new_n813), .B2(new_n815), .C1(new_n816), .C2(new_n632), .ZN(new_n817));
  AOI22_X1  g0617(.A1(G58), .A2(new_n793), .B1(new_n800), .B2(G50), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n813), .A2(new_n815), .B1(new_n810), .B2(G97), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(new_n206), .C2(new_n788), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n817), .B(new_n820), .C1(G68), .C2(new_n795), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n780), .B1(new_n811), .B2(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(G13), .A2(G33), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n824), .A2(G20), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n773), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n254), .A2(G45), .ZN(new_n827));
  XNOR2_X1  g0627(.A(new_n827), .B(KEYINPUT100), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n213), .A2(new_n342), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G45), .C2(new_n235), .ZN(new_n830));
  INV_X1    g0630(.A(G355), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n214), .A2(new_n342), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n830), .B1(G116), .B2(new_n214), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n780), .A2(new_n825), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND4_X1  g0635(.A1(new_n822), .A2(new_n826), .A3(new_n772), .A4(new_n835), .ZN(new_n836));
  AND2_X1   g0636(.A1(new_n778), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(G396));
  NOR2_X1   g0638(.A1(new_n459), .A2(new_n710), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n340), .A2(new_n710), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n363), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n839), .B1(new_n841), .B2(new_n459), .ZN(new_n842));
  OR2_X1    g0642(.A1(new_n764), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n700), .A2(new_n756), .A3(new_n842), .ZN(new_n844));
  AND2_X1   g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(KEYINPUT31), .B1(new_n665), .B2(new_n710), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n751), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n774), .B1(new_n847), .B2(new_n759), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n849), .B(KEYINPUT105), .Z(new_n850));
  OAI211_X1 g0650(.A(new_n850), .B(new_n771), .C1(new_n848), .C2(new_n845), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n787), .A2(G68), .B1(G132), .B2(new_n805), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n852), .B(new_n342), .C1(new_n202), .C2(new_n816), .ZN(new_n853));
  AOI22_X1  g0653(.A1(G143), .A2(new_n793), .B1(new_n795), .B2(G150), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n800), .A2(G137), .ZN(new_n855));
  OAI211_X1 g0655(.A(new_n854), .B(new_n855), .C1(new_n814), .C2(new_n802), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT34), .Z(new_n857));
  AOI211_X1 g0657(.A(new_n853), .B(new_n857), .C1(G58), .C2(new_n810), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n342), .B1(new_n805), .B2(G311), .ZN(new_n859));
  OAI221_X1 g0659(.A(new_n859), .B1(new_n205), .B2(new_n809), .C1(new_n788), .C2(new_n632), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G294), .A2(new_n793), .B1(new_n800), .B2(G303), .ZN(new_n861));
  INV_X1    g0661(.A(new_n795), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n861), .B1(new_n786), .B2(new_n862), .C1(new_n206), .C2(new_n816), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n860), .B(new_n863), .C1(G116), .C2(new_n803), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n780), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n842), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n823), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n780), .A2(new_n823), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(new_n261), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n865), .A2(new_n772), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n851), .A2(new_n870), .ZN(G384));
  INV_X1    g0671(.A(KEYINPUT108), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n759), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g0673(.A1(new_n750), .A2(KEYINPUT108), .A3(KEYINPUT31), .A4(new_n710), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n847), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n876), .A2(new_n687), .A3(G330), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n325), .A2(new_n331), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n279), .A2(new_n756), .ZN(new_n880));
  OAI22_X1  g0680(.A1(new_n879), .A2(new_n880), .B1(new_n325), .B2(new_n756), .ZN(new_n881));
  INV_X1    g0681(.A(new_n875), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n842), .B(new_n881), .C1(new_n758), .C2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(new_n708), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n383), .A2(new_n257), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n380), .B(G68), .C1(new_n379), .C2(new_n369), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n886), .B2(new_n378), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n408), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n420), .B1(new_n386), .B2(new_n408), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n891), .A2(new_n423), .A3(KEYINPUT18), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n428), .A2(new_n680), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n890), .B1(new_n893), .B2(new_n677), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT38), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n386), .A2(new_n402), .A3(new_n408), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n896), .A2(new_n891), .A3(KEYINPUT37), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n417), .A2(new_n884), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n421), .B1(new_n888), .B2(new_n889), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n890), .A2(new_n899), .A3(new_n409), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n897), .A2(new_n898), .B1(new_n900), .B2(KEYINPUT37), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n681), .A2(new_n677), .ZN(new_n903));
  INV_X1    g0703(.A(new_n898), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT37), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n896), .A2(new_n891), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n904), .B1(new_n907), .B2(KEYINPUT106), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n679), .A2(new_n409), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT106), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n906), .B1(new_n908), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n897), .A2(KEYINPUT107), .A3(new_n898), .ZN(new_n913));
  NAND4_X1  g0713(.A1(new_n679), .A2(new_n898), .A3(new_n906), .A4(new_n409), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT107), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n905), .B1(new_n912), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n902), .B1(new_n895), .B2(new_n918), .ZN(new_n919));
  OAI21_X1  g0719(.A(KEYINPUT40), .B1(new_n883), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n895), .B1(new_n894), .B2(new_n901), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n900), .A2(KEYINPUT37), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n914), .ZN(new_n923));
  OAI211_X1 g0723(.A(KEYINPUT38), .B(new_n923), .C1(new_n429), .C2(new_n890), .ZN(new_n924));
  AOI21_X1  g0724(.A(KEYINPUT40), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND4_X1  g0725(.A1(new_n876), .A2(new_n925), .A3(new_n842), .A4(new_n881), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n878), .B1(new_n927), .B2(G330), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n876), .A2(new_n687), .ZN(new_n929));
  INV_X1    g0729(.A(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n928), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n681), .A2(new_n884), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT39), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n914), .B(KEYINPUT107), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n898), .B1(new_n909), .B2(new_n910), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n907), .A2(KEYINPUT106), .ZN(new_n936));
  OAI21_X1  g0736(.A(KEYINPUT37), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI22_X1  g0737(.A1(new_n934), .A2(new_n937), .B1(new_n904), .B2(new_n903), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n933), .B(new_n924), .C1(new_n938), .C2(KEYINPUT38), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n921), .A2(new_n924), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(KEYINPUT39), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n672), .A2(new_n756), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n932), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n839), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n844), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n940), .A2(new_n947), .A3(new_n881), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n931), .B(new_n949), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n687), .A2(new_n765), .A3(new_n766), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n682), .A2(new_n454), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n951), .B(new_n457), .C1(new_n952), .C2(new_n684), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n950), .B(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n209), .B2(new_n704), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n248), .B1(new_n522), .B2(KEYINPUT35), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n956), .B(new_n233), .C1(KEYINPUT35), .C2(new_n522), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n957), .B(KEYINPUT36), .ZN(new_n958));
  OR2_X1    g0758(.A1(new_n235), .A2(new_n372), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n959), .A2(new_n220), .B1(G50), .B2(new_n274), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n960), .A2(G1), .A3(new_n212), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n955), .A2(new_n958), .A3(new_n961), .ZN(G367));
  INV_X1    g0762(.A(new_n730), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n714), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n533), .B1(new_n526), .B2(new_n756), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n530), .A2(new_n532), .A3(new_n710), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT42), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n968), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n696), .B1(new_n965), .B2(new_n570), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n756), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OR3_X1    g0773(.A1(new_n646), .A2(new_n651), .A3(new_n756), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n689), .B1(new_n651), .B2(new_n756), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT43), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n973), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n970), .A2(new_n978), .A3(new_n977), .A4(new_n972), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n714), .B1(new_n777), .B2(new_n776), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n984), .A2(new_n967), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n983), .B(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n736), .B(KEYINPUT41), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n724), .A2(new_n727), .A3(new_n715), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n963), .B1(new_n989), .B2(new_n984), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n777), .A2(new_n776), .A3(new_n714), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n728), .A2(new_n730), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n990), .A2(new_n761), .A3(new_n992), .A4(new_n767), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT110), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n967), .A2(new_n731), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(KEYINPUT109), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT109), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n967), .A2(new_n998), .A3(new_n731), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT45), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n967), .A2(new_n731), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n997), .A2(KEYINPUT45), .A3(new_n999), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1002), .A2(new_n1004), .A3(new_n728), .A4(new_n1005), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n768), .A2(KEYINPUT110), .A3(new_n992), .A4(new_n990), .ZN(new_n1007));
  NAND3_X1  g0807(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n984), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n995), .A2(new_n1006), .A3(new_n1007), .A4(new_n1009), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n988), .B1(new_n1010), .B2(new_n768), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n770), .A2(G1), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n1012), .B(KEYINPUT111), .Z(new_n1013));
  OAI21_X1  g0813(.A(new_n986), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n788), .A2(new_n205), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n342), .B1(new_n805), .B2(G317), .ZN(new_n1016));
  INV_X1    g0816(.A(G294), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1016), .B1(new_n862), .B2(new_n1017), .ZN(new_n1018));
  AOI211_X1 g0818(.A(new_n1015), .B(new_n1018), .C1(G283), .C2(new_n803), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n800), .A2(G311), .B1(G107), .B2(new_n810), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n793), .A2(G303), .ZN(new_n1021));
  AOI21_X1  g0821(.A(KEYINPUT112), .B1(new_n783), .B2(G116), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT46), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n783), .A2(G58), .B1(G137), .B2(new_n805), .ZN(new_n1025));
  XOR2_X1   g0825(.A(new_n1025), .B(KEYINPUT114), .Z(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(G50), .B2(new_n803), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n793), .A2(G150), .B1(G68), .B2(new_n810), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n800), .A2(G143), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n795), .A2(G159), .ZN(new_n1030));
  NAND4_X1  g0830(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .A4(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n346), .B1(new_n787), .B2(new_n221), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT113), .Z(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1035), .A2(new_n780), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n977), .A2(new_n825), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n829), .ZN(new_n1038));
  OAI221_X1 g0838(.A(new_n834), .B1(new_n214), .B2(new_n336), .C1(new_n241), .C2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1036), .A2(new_n772), .A3(new_n1037), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1014), .A2(new_n1040), .ZN(G387));
  INV_X1    g0841(.A(new_n768), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n990), .A2(new_n992), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1044), .A2(new_n736), .A3(new_n993), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(G311), .A2(new_n795), .B1(new_n793), .B2(G317), .ZN(new_n1046));
  INV_X1    g0846(.A(G322), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1046), .B1(new_n573), .B2(new_n802), .C1(new_n1047), .C2(new_n799), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT48), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1049), .B1(new_n786), .B2(new_n809), .C1(new_n1017), .C2(new_n816), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT49), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n342), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n805), .A2(G326), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n787), .A2(G116), .ZN(new_n1055));
  NAND4_X1  g0855(.A1(new_n1052), .A2(new_n1053), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n810), .A2(new_n335), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1057), .B1(new_n432), .B2(new_n804), .C1(new_n862), .C2(new_n406), .ZN(new_n1058));
  AOI211_X1 g0858(.A(new_n346), .B(new_n1058), .C1(G50), .C2(new_n793), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n783), .A2(new_n221), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n803), .A2(G68), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1015), .B1(G159), .B2(new_n800), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1060), .A3(new_n1061), .A4(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1056), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n829), .B1(new_n245), .B2(new_n300), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1065), .B1(new_n735), .B2(new_n832), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n333), .A2(new_n202), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1067), .B(KEYINPUT50), .Z(new_n1068));
  AOI21_X1  g0868(.A(new_n734), .B1(G68), .B2(G77), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1068), .A2(new_n300), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1066), .A2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n213), .A2(new_n206), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n1064), .A2(new_n780), .B1(new_n834), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n825), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n772), .C1(new_n715), .C2(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1013), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1045), .B(new_n1076), .C1(new_n1043), .C2(new_n1077), .ZN(G393));
  NAND2_X1  g0878(.A1(new_n1009), .A2(new_n1006), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1079), .A2(new_n1077), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n967), .A2(new_n1075), .ZN(new_n1081));
  XOR2_X1   g0881(.A(new_n1081), .B(KEYINPUT115), .Z(new_n1082));
  AOI22_X1  g0882(.A1(G311), .A2(new_n793), .B1(new_n800), .B2(G317), .ZN(new_n1083));
  XNOR2_X1  g0883(.A(new_n1083), .B(KEYINPUT52), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n816), .A2(new_n786), .B1(new_n1047), .B2(new_n804), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  OAI22_X1  g0886(.A1(new_n1085), .A2(new_n1086), .B1(new_n206), .B2(new_n788), .ZN(new_n1087));
  NOR3_X1   g0887(.A1(new_n1084), .A2(new_n1087), .A3(new_n342), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n862), .A2(new_n573), .B1(new_n248), .B2(new_n809), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1089), .A2(KEYINPUT118), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n1089), .A2(KEYINPUT118), .B1(G294), .B2(new_n803), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(G50), .A2(new_n795), .B1(new_n803), .B2(new_n333), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n1094), .A2(KEYINPUT116), .B1(new_n274), .B2(new_n816), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G87), .B2(new_n787), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n793), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n1097), .A2(new_n814), .B1(new_n432), .B2(new_n799), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT51), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n809), .A2(new_n261), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n805), .A2(G143), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n1094), .C2(KEYINPUT116), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1096), .A2(new_n1099), .A3(new_n342), .A4(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1093), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(new_n780), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n834), .B1(new_n205), .B2(new_n214), .C1(new_n251), .C2(new_n1038), .ZN(new_n1106));
  AND4_X1   g0906(.A1(new_n772), .A2(new_n1082), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1080), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1079), .A2(new_n993), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1109), .A2(new_n1010), .A3(new_n736), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1108), .A2(new_n1110), .ZN(G390));
  NAND2_X1  g0911(.A1(new_n947), .A2(new_n881), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n941), .A2(new_n939), .B1(new_n1112), .B2(new_n943), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n839), .B1(new_n764), .B2(new_n842), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n672), .A2(new_n675), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n880), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1115), .A2(new_n1116), .B1(new_n672), .B2(new_n710), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n943), .B1(new_n1114), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n924), .B1(new_n938), .B2(KEYINPUT38), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n848), .A2(new_n842), .ZN(new_n1121));
  OAI22_X1  g0921(.A1(new_n1113), .A2(new_n1120), .B1(new_n1117), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT120), .ZN(new_n1123));
  OAI21_X1  g0923(.A(KEYINPUT119), .B1(new_n1113), .B2(new_n1120), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT119), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n944), .B1(new_n947), .B2(new_n881), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n919), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n933), .B1(new_n921), .B2(new_n924), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n919), .B2(new_n933), .ZN(new_n1129));
  OAI211_X1 g0929(.A(new_n1125), .B(new_n1127), .C1(new_n1129), .C2(new_n1126), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  AOI22_X1  g0931(.A1(new_n846), .A2(new_n751), .B1(new_n873), .B2(new_n874), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(new_n866), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1133), .A2(G330), .A3(new_n881), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1123), .B1(new_n1131), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(KEYINPUT120), .B(new_n1134), .C1(new_n1124), .C2(new_n1130), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1122), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n686), .A2(KEYINPUT121), .A3(new_n951), .A4(new_n877), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT121), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1140), .B1(new_n953), .B2(new_n878), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1142));
  AND4_X1   g0942(.A1(new_n848), .A2(new_n842), .A3(new_n1112), .A4(new_n1142), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n1133), .A2(G330), .B1(new_n1112), .B2(new_n1142), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1139), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1138), .A2(new_n1146), .ZN(new_n1147));
  AND3_X1   g0947(.A1(new_n1139), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1122), .B(new_n1148), .C1(new_n1136), .C2(new_n1137), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1147), .A2(new_n736), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1129), .A2(new_n823), .ZN(new_n1151));
  XOR2_X1   g0951(.A(KEYINPUT54), .B(G143), .Z(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  OAI221_X1 g0953(.A(new_n342), .B1(new_n814), .B2(new_n809), .C1(new_n802), .C2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n793), .A2(G132), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n788), .B2(new_n202), .ZN(new_n1156));
  AOI211_X1 g0956(.A(new_n1154), .B(new_n1156), .C1(G125), .C2(new_n805), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n783), .A2(G150), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT53), .Z(new_n1159));
  AOI22_X1  g0959(.A1(G137), .A2(new_n795), .B1(new_n800), .B2(G128), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT122), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G116), .A2(new_n793), .B1(new_n800), .B2(G283), .ZN(new_n1163));
  OAI221_X1 g0963(.A(new_n1163), .B1(new_n205), .B2(new_n802), .C1(new_n206), .C2(new_n862), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G68), .B2(new_n787), .ZN(new_n1165));
  AOI22_X1  g0965(.A1(new_n783), .A2(G87), .B1(G294), .B2(new_n805), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1167), .A2(new_n342), .A3(new_n1100), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n780), .B1(new_n1162), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n868), .A2(new_n406), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1151), .A2(new_n772), .A3(new_n1169), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1138), .B2(new_n1077), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1150), .A2(new_n1173), .ZN(G378));
  NAND2_X1  g0974(.A1(new_n454), .A2(new_n457), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n435), .A2(new_n884), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n454), .A2(new_n457), .A3(new_n1176), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1180), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1183), .A2(new_n823), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n787), .A2(G58), .ZN(new_n1185));
  OAI211_X1 g0985(.A(new_n1185), .B(new_n346), .C1(new_n248), .C2(new_n799), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n795), .A2(G97), .B1(G68), .B2(new_n810), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n206), .B2(new_n1097), .ZN(new_n1188));
  AOI211_X1 g0988(.A(G41), .B(new_n1188), .C1(new_n335), .C2(new_n803), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1060), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1186), .B(new_n1190), .C1(G283), .C2(new_n805), .ZN(new_n1191));
  OR2_X1    g0991(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT58), .ZN(new_n1193));
  INV_X1    g0993(.A(G124), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n258), .B1(new_n804), .B2(new_n1194), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G132), .A2(new_n795), .B1(new_n800), .B2(G125), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n783), .A2(new_n1152), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n793), .A2(G128), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n803), .A2(G137), .B1(G150), .B2(new_n810), .ZN(new_n1199));
  NAND4_X1  g0999(.A1(new_n1196), .A2(new_n1197), .A3(new_n1198), .A4(new_n1199), .ZN(new_n1200));
  AOI211_X1 g1000(.A(G41), .B(new_n1195), .C1(new_n1200), .C2(KEYINPUT59), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(KEYINPUT59), .B2(new_n1200), .C1(new_n814), .C2(new_n788), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n202), .B1(new_n283), .B2(G41), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1192), .A2(new_n1193), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n780), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n868), .A2(new_n202), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1184), .A2(new_n772), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1183), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1208), .B1(new_n927), .B2(G330), .ZN(new_n1209));
  AOI211_X1 g1009(.A(new_n774), .B(new_n1183), .C1(new_n920), .C2(new_n926), .ZN(new_n1210));
  NOR3_X1   g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n949), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n949), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1119), .A2(new_n876), .A3(new_n842), .A4(new_n881), .ZN(new_n1213));
  NOR3_X1   g1013(.A1(new_n1132), .A2(new_n866), .A3(new_n1117), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1213), .A2(KEYINPUT40), .B1(new_n1214), .B2(new_n925), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1183), .B1(new_n1215), .B2(new_n774), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n927), .A2(G330), .A3(new_n1208), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1212), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1211), .A2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1207), .B1(new_n1219), .B2(new_n1077), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1219), .B1(new_n1149), .B2(new_n1223), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n736), .B1(new_n1224), .B2(KEYINPUT57), .ZN(new_n1225));
  INV_X1    g1025(.A(KEYINPUT57), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1226), .B(new_n1219), .C1(new_n1223), .C2(new_n1149), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1221), .B1(new_n1225), .B2(new_n1227), .ZN(G375));
  NAND2_X1  g1028(.A1(new_n1117), .A2(new_n823), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n342), .B1(new_n805), .B2(G303), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1057), .B(new_n1230), .C1(new_n816), .C2(new_n205), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G283), .A2(new_n793), .B1(new_n800), .B2(G294), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n248), .B2(new_n862), .C1(new_n261), .C2(new_n788), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G107), .C2(new_n803), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(G137), .A2(new_n793), .B1(new_n800), .B2(G132), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n805), .A2(G128), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1235), .A2(new_n1185), .A3(new_n1236), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n342), .B1(new_n202), .B2(new_n809), .C1(new_n862), .C2(new_n1153), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n816), .A2(new_n814), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n802), .A2(new_n432), .ZN(new_n1240));
  NOR4_X1   g1040(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1240), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n780), .B1(new_n1234), .B2(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n868), .A2(new_n274), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1229), .A2(new_n772), .A3(new_n1242), .A4(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1145), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1244), .B1(new_n1245), .B2(new_n1077), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT123), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT123), .ZN(new_n1248));
  OAI211_X1 g1048(.A(new_n1248), .B(new_n1244), .C1(new_n1245), .C2(new_n1077), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1222), .A2(new_n1245), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1251), .A2(new_n987), .A3(new_n1146), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(G381));
  NAND2_X1  g1053(.A1(new_n1149), .A2(new_n1223), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1219), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1226), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1224), .A2(KEYINPUT57), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1257), .A2(new_n736), .A3(new_n1258), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1149), .A2(new_n736), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1172), .B1(new_n1260), .B2(new_n1147), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1261), .A3(new_n1221), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(G390), .ZN(new_n1264));
  OR3_X1    g1064(.A1(G384), .A2(G393), .A3(G396), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G387), .ZN(new_n1268));
  AOI21_X1  g1068(.A(G381), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1263), .A2(new_n1264), .A3(new_n1268), .A4(new_n1269), .ZN(G407));
  OAI211_X1 g1070(.A(G407), .B(G213), .C1(G343), .C2(new_n1262), .ZN(G409));
  AOI21_X1  g1071(.A(new_n1220), .B1(new_n1224), .B2(new_n987), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1272), .A2(new_n1261), .B1(G213), .B2(new_n709), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1222), .A2(KEYINPUT60), .A3(new_n1245), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1274), .A2(new_n736), .A3(new_n1146), .ZN(new_n1275));
  AOI21_X1  g1075(.A(KEYINPUT60), .B1(new_n1222), .B2(new_n1245), .ZN(new_n1276));
  OAI211_X1 g1076(.A(new_n1250), .B(G384), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1251), .A2(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1280), .A2(new_n736), .A3(new_n1146), .A4(new_n1274), .ZN(new_n1281));
  AOI21_X1  g1081(.A(G384), .B1(new_n1281), .B2(new_n1250), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1278), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n737), .B1(new_n1256), .B2(new_n1226), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1220), .B1(new_n1284), .B2(new_n1258), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1273), .B(new_n1283), .C1(new_n1285), .C2(new_n1261), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT61), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1281), .A2(new_n1250), .ZN(new_n1289));
  INV_X1    g1089(.A(G384), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n709), .A2(G213), .A3(G2897), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1291), .A2(new_n1277), .A3(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(new_n1292), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n1278), .B2(new_n1282), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1293), .A2(new_n1295), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1261), .B1(new_n1259), .B2(new_n1221), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n709), .A2(G213), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1254), .A2(new_n987), .A3(new_n1255), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1300), .A2(new_n1221), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1301), .B2(G378), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1297), .B1(new_n1298), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(G375), .A2(G378), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT62), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1304), .A2(new_n1305), .A3(new_n1273), .A4(new_n1283), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1287), .A2(new_n1288), .A3(new_n1303), .A4(new_n1306), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(G393), .B(new_n837), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(G387), .A2(new_n1264), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1014), .A2(new_n1040), .A3(G390), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1309), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT125), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1311), .A2(new_n1313), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1014), .A2(KEYINPUT125), .A3(new_n1040), .A4(G390), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1314), .A2(new_n1310), .A3(new_n1309), .A4(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1316), .A2(KEYINPUT126), .ZN(new_n1317));
  AOI21_X1  g1117(.A(G390), .B1(new_n1014), .B2(new_n1040), .ZN(new_n1318));
  AND3_X1   g1118(.A1(new_n1014), .A2(new_n1040), .A3(G390), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1318), .B1(new_n1319), .B2(KEYINPUT125), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT126), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1308), .B1(new_n1311), .B2(new_n1313), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  AOI21_X1  g1123(.A(new_n1312), .B1(new_n1317), .B2(new_n1323), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1307), .A2(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1296), .B1(new_n1304), .B2(new_n1273), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT63), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1286), .B1(new_n1326), .B2(new_n1327), .ZN(new_n1328));
  NOR2_X1   g1128(.A1(new_n1324), .A2(KEYINPUT61), .ZN(new_n1329));
  OAI21_X1  g1129(.A(KEYINPUT127), .B1(new_n1286), .B2(new_n1327), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1302), .B1(G378), .B2(G375), .ZN(new_n1331));
  INV_X1    g1131(.A(KEYINPUT127), .ZN(new_n1332));
  NAND4_X1  g1132(.A1(new_n1331), .A2(new_n1332), .A3(KEYINPUT63), .A4(new_n1283), .ZN(new_n1333));
  NAND4_X1  g1133(.A1(new_n1328), .A2(new_n1329), .A3(new_n1330), .A4(new_n1333), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1325), .A2(new_n1334), .ZN(G405));
  AND2_X1   g1135(.A1(new_n1304), .A2(new_n1262), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1312), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1316), .A2(KEYINPUT126), .ZN(new_n1338));
  AOI21_X1  g1138(.A(new_n1321), .B1(new_n1320), .B2(new_n1322), .ZN(new_n1339));
  OAI21_X1  g1139(.A(new_n1337), .B1(new_n1338), .B2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1324), .B1(new_n1263), .B2(new_n1298), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1341), .A2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1283), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND3_X1  g1145(.A1(new_n1341), .A2(new_n1342), .A3(new_n1283), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1345), .A2(new_n1346), .ZN(G402));
endmodule


