

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XNOR2_X1 U323 ( .A(n347), .B(n346), .ZN(n377) );
  INV_X1 U324 ( .A(G204GAT), .ZN(n344) );
  XNOR2_X1 U325 ( .A(n345), .B(n344), .ZN(n346) );
  INV_X1 U326 ( .A(KEYINPUT55), .ZN(n451) );
  XNOR2_X1 U327 ( .A(n451), .B(KEYINPUT121), .ZN(n452) );
  XNOR2_X1 U328 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U329 ( .A(n574), .B(KEYINPUT41), .Z(n558) );
  XNOR2_X1 U330 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n455) );
  XNOR2_X1 U331 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XOR2_X1 U332 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n292) );
  XNOR2_X1 U333 ( .A(G218GAT), .B(G92GAT), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n296) );
  XOR2_X1 U335 ( .A(KEYINPUT80), .B(KEYINPUT10), .Z(n294) );
  XNOR2_X1 U336 ( .A(G134GAT), .B(G162GAT), .ZN(n293) );
  XNOR2_X1 U337 ( .A(n294), .B(n293), .ZN(n295) );
  XOR2_X1 U338 ( .A(n296), .B(n295), .Z(n305) );
  XOR2_X1 U339 ( .A(G99GAT), .B(G85GAT), .Z(n372) );
  XNOR2_X1 U340 ( .A(G190GAT), .B(KEYINPUT81), .ZN(n297) );
  NAND2_X1 U341 ( .A1(KEYINPUT78), .A2(n297), .ZN(n300) );
  INV_X1 U342 ( .A(KEYINPUT78), .ZN(n298) );
  XOR2_X1 U343 ( .A(G190GAT), .B(KEYINPUT81), .Z(n412) );
  NAND2_X1 U344 ( .A1(n298), .A2(n412), .ZN(n299) );
  NAND2_X1 U345 ( .A1(n300), .A2(n299), .ZN(n302) );
  NAND2_X1 U346 ( .A1(G232GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U347 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U348 ( .A(n372), .B(n303), .ZN(n304) );
  XNOR2_X1 U349 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U350 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n307) );
  XNOR2_X1 U351 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n306) );
  XNOR2_X1 U352 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U353 ( .A(n309), .B(n308), .ZN(n314) );
  XOR2_X1 U354 ( .A(G29GAT), .B(KEYINPUT7), .Z(n311) );
  XNOR2_X1 U355 ( .A(G43GAT), .B(G36GAT), .ZN(n310) );
  XNOR2_X1 U356 ( .A(n311), .B(n310), .ZN(n313) );
  XOR2_X1 U357 ( .A(G50GAT), .B(KEYINPUT8), .Z(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n364) );
  XNOR2_X1 U359 ( .A(n314), .B(n364), .ZN(n551) );
  XOR2_X1 U360 ( .A(G183GAT), .B(KEYINPUT17), .Z(n316) );
  XNOR2_X1 U361 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n422) );
  XOR2_X1 U363 ( .A(G120GAT), .B(G71GAT), .Z(n378) );
  XOR2_X1 U364 ( .A(n422), .B(n378), .Z(n318) );
  XNOR2_X1 U365 ( .A(G99GAT), .B(G190GAT), .ZN(n317) );
  XNOR2_X1 U366 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U367 ( .A(G15GAT), .B(G176GAT), .Z(n320) );
  NAND2_X1 U368 ( .A1(G227GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U369 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U370 ( .A(n322), .B(n321), .Z(n327) );
  XOR2_X1 U371 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n324) );
  XNOR2_X1 U372 ( .A(G43GAT), .B(KEYINPUT85), .ZN(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(n325), .ZN(n326) );
  XNOR2_X1 U375 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U376 ( .A(KEYINPUT84), .B(G134GAT), .Z(n329) );
  XNOR2_X1 U377 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n328) );
  XNOR2_X1 U378 ( .A(n329), .B(n328), .ZN(n330) );
  XOR2_X1 U379 ( .A(G113GAT), .B(n330), .Z(n446) );
  XOR2_X2 U380 ( .A(n331), .B(n446), .Z(n528) );
  XOR2_X1 U381 ( .A(KEYINPUT22), .B(KEYINPUT90), .Z(n333) );
  XNOR2_X1 U382 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n332) );
  XNOR2_X1 U383 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U384 ( .A(n334), .B(KEYINPUT87), .Z(n336) );
  XOR2_X1 U385 ( .A(G141GAT), .B(G22GAT), .Z(n356) );
  XNOR2_X1 U386 ( .A(G50GAT), .B(n356), .ZN(n335) );
  XNOR2_X1 U387 ( .A(n336), .B(n335), .ZN(n342) );
  XOR2_X1 U388 ( .A(G211GAT), .B(KEYINPUT21), .Z(n338) );
  XNOR2_X1 U389 ( .A(G197GAT), .B(G218GAT), .ZN(n337) );
  XNOR2_X1 U390 ( .A(n338), .B(n337), .ZN(n414) );
  XOR2_X1 U391 ( .A(KEYINPUT88), .B(n414), .Z(n340) );
  NAND2_X1 U392 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U393 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U394 ( .A(n342), .B(n341), .Z(n352) );
  XNOR2_X1 U395 ( .A(G148GAT), .B(KEYINPUT73), .ZN(n343) );
  XNOR2_X1 U396 ( .A(n343), .B(KEYINPUT74), .ZN(n347) );
  XNOR2_X1 U397 ( .A(G78GAT), .B(G106GAT), .ZN(n345) );
  XOR2_X1 U398 ( .A(KEYINPUT89), .B(G162GAT), .Z(n349) );
  XNOR2_X1 U399 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U401 ( .A(KEYINPUT2), .B(n350), .Z(n436) );
  XNOR2_X1 U402 ( .A(n377), .B(n436), .ZN(n351) );
  XNOR2_X1 U403 ( .A(n352), .B(n351), .ZN(n467) );
  XOR2_X1 U404 ( .A(KEYINPUT67), .B(KEYINPUT68), .Z(n354) );
  XNOR2_X1 U405 ( .A(KEYINPUT30), .B(KEYINPUT29), .ZN(n353) );
  XNOR2_X1 U406 ( .A(n354), .B(n353), .ZN(n363) );
  XNOR2_X1 U407 ( .A(G15GAT), .B(G1GAT), .ZN(n355) );
  XNOR2_X1 U408 ( .A(n355), .B(KEYINPUT69), .ZN(n396) );
  XOR2_X1 U409 ( .A(n356), .B(n396), .Z(n358) );
  NAND2_X1 U410 ( .A1(G229GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U411 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U412 ( .A(G169GAT), .B(G8GAT), .Z(n413) );
  XOR2_X1 U413 ( .A(n359), .B(n413), .Z(n361) );
  XNOR2_X1 U414 ( .A(G197GAT), .B(G113GAT), .ZN(n360) );
  XNOR2_X1 U415 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U416 ( .A(n363), .B(n362), .ZN(n365) );
  XNOR2_X1 U417 ( .A(n365), .B(n364), .ZN(n571) );
  XNOR2_X1 U418 ( .A(KEYINPUT31), .B(KEYINPUT33), .ZN(n371) );
  XOR2_X1 U419 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n367) );
  XNOR2_X1 U420 ( .A(KEYINPUT72), .B(KEYINPUT71), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n369) );
  XNOR2_X1 U422 ( .A(G176GAT), .B(G92GAT), .ZN(n368) );
  XNOR2_X1 U423 ( .A(n368), .B(G64GAT), .ZN(n421) );
  XNOR2_X1 U424 ( .A(n369), .B(n421), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n376) );
  XOR2_X1 U426 ( .A(G57GAT), .B(KEYINPUT13), .Z(n392) );
  XOR2_X1 U427 ( .A(n372), .B(n392), .Z(n374) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n380) );
  XNOR2_X1 U431 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U432 ( .A(n380), .B(n379), .Z(n574) );
  NAND2_X1 U433 ( .A1(n571), .A2(n558), .ZN(n382) );
  INV_X1 U434 ( .A(KEYINPUT46), .ZN(n381) );
  XOR2_X1 U435 ( .A(n382), .B(n381), .Z(n401) );
  XOR2_X1 U436 ( .A(G64GAT), .B(G183GAT), .Z(n384) );
  XNOR2_X1 U437 ( .A(G127GAT), .B(G71GAT), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n388) );
  XOR2_X1 U439 ( .A(KEYINPUT83), .B(KEYINPUT15), .Z(n386) );
  XNOR2_X1 U440 ( .A(G8GAT), .B(KEYINPUT14), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n400) );
  XOR2_X1 U443 ( .A(G211GAT), .B(G155GAT), .Z(n390) );
  XNOR2_X1 U444 ( .A(G22GAT), .B(G78GAT), .ZN(n389) );
  XNOR2_X1 U445 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U446 ( .A(n392), .B(n391), .Z(n394) );
  NAND2_X1 U447 ( .A1(G231GAT), .A2(G233GAT), .ZN(n393) );
  XNOR2_X1 U448 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U449 ( .A(n395), .B(KEYINPUT82), .Z(n398) );
  XNOR2_X1 U450 ( .A(n396), .B(KEYINPUT12), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U452 ( .A(n400), .B(n399), .Z(n534) );
  INV_X1 U453 ( .A(n534), .ZN(n549) );
  NAND2_X1 U454 ( .A1(n401), .A2(n549), .ZN(n402) );
  NOR2_X1 U455 ( .A1(n551), .A2(n402), .ZN(n403) );
  XNOR2_X1 U456 ( .A(n403), .B(KEYINPUT47), .ZN(n409) );
  INV_X1 U457 ( .A(n571), .ZN(n503) );
  XOR2_X1 U458 ( .A(KEYINPUT70), .B(n503), .Z(n556) );
  XNOR2_X1 U459 ( .A(KEYINPUT36), .B(n551), .ZN(n579) );
  NAND2_X1 U460 ( .A1(n534), .A2(n579), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n404), .B(KEYINPUT112), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n405), .B(KEYINPUT45), .ZN(n406) );
  NOR2_X1 U463 ( .A1(n556), .A2(n406), .ZN(n407) );
  INV_X1 U464 ( .A(n574), .ZN(n457) );
  NAND2_X1 U465 ( .A1(n407), .A2(n457), .ZN(n408) );
  NAND2_X1 U466 ( .A1(n409), .A2(n408), .ZN(n411) );
  XNOR2_X1 U467 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n410) );
  XNOR2_X1 U468 ( .A(n411), .B(n410), .ZN(n525) );
  XNOR2_X1 U469 ( .A(n413), .B(n412), .ZN(n426) );
  XOR2_X1 U470 ( .A(n414), .B(KEYINPUT96), .Z(n416) );
  NAND2_X1 U471 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U473 ( .A(KEYINPUT95), .B(KEYINPUT97), .Z(n418) );
  XNOR2_X1 U474 ( .A(G36GAT), .B(G204GAT), .ZN(n417) );
  XNOR2_X1 U475 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U476 ( .A(n420), .B(n419), .Z(n424) );
  XNOR2_X1 U477 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(n426), .B(n425), .Z(n518) );
  INV_X1 U480 ( .A(n518), .ZN(n427) );
  NAND2_X1 U481 ( .A1(n525), .A2(n427), .ZN(n429) );
  XOR2_X1 U482 ( .A(KEYINPUT120), .B(KEYINPUT54), .Z(n428) );
  XNOR2_X1 U483 ( .A(n429), .B(n428), .ZN(n449) );
  XOR2_X1 U484 ( .A(KEYINPUT91), .B(KEYINPUT6), .Z(n431) );
  XNOR2_X1 U485 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n430) );
  XNOR2_X1 U486 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U487 ( .A(KEYINPUT4), .B(n432), .Z(n434) );
  NAND2_X1 U488 ( .A1(G225GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U490 ( .A(n435), .B(KEYINPUT94), .Z(n438) );
  XNOR2_X1 U491 ( .A(n436), .B(KEYINPUT92), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U493 ( .A(G85GAT), .B(G148GAT), .Z(n440) );
  XNOR2_X1 U494 ( .A(G29GAT), .B(G141GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U496 ( .A(n442), .B(n441), .Z(n448) );
  XOR2_X1 U497 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n444) );
  XNOR2_X1 U498 ( .A(G1GAT), .B(G120GAT), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U501 ( .A(n448), .B(n447), .ZN(n516) );
  NAND2_X1 U502 ( .A1(n449), .A2(n516), .ZN(n450) );
  XOR2_X1 U503 ( .A(n450), .B(KEYINPUT65), .Z(n569) );
  NOR2_X1 U504 ( .A1(n467), .A2(n569), .ZN(n453) );
  NOR2_X1 U505 ( .A1(n528), .A2(n454), .ZN(n563) );
  NAND2_X1 U506 ( .A1(n551), .A2(n563), .ZN(n456) );
  NAND2_X1 U507 ( .A1(n556), .A2(n457), .ZN(n491) );
  NOR2_X1 U508 ( .A1(n549), .A2(n551), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(KEYINPUT16), .ZN(n474) );
  NAND2_X1 U510 ( .A1(n467), .A2(n528), .ZN(n459) );
  XNOR2_X1 U511 ( .A(n459), .B(KEYINPUT26), .ZN(n570) );
  XNOR2_X1 U512 ( .A(n518), .B(KEYINPUT27), .ZN(n469) );
  NOR2_X1 U513 ( .A1(n570), .A2(n469), .ZN(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT99), .B(n460), .ZN(n464) );
  NOR2_X1 U515 ( .A1(n528), .A2(n518), .ZN(n461) );
  NOR2_X1 U516 ( .A1(n467), .A2(n461), .ZN(n462) );
  XNOR2_X1 U517 ( .A(KEYINPUT25), .B(n462), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n464), .A2(n463), .ZN(n465) );
  NAND2_X1 U519 ( .A1(n516), .A2(n465), .ZN(n466) );
  XNOR2_X1 U520 ( .A(KEYINPUT100), .B(n466), .ZN(n473) );
  XNOR2_X1 U521 ( .A(n467), .B(KEYINPUT66), .ZN(n468) );
  XOR2_X1 U522 ( .A(n468), .B(KEYINPUT28), .Z(n522) );
  INV_X1 U523 ( .A(n522), .ZN(n527) );
  NOR2_X1 U524 ( .A1(n516), .A2(n469), .ZN(n526) );
  NAND2_X1 U525 ( .A1(n528), .A2(n526), .ZN(n470) );
  NOR2_X1 U526 ( .A1(n527), .A2(n470), .ZN(n471) );
  XOR2_X1 U527 ( .A(KEYINPUT98), .B(n471), .Z(n472) );
  NAND2_X1 U528 ( .A1(n473), .A2(n472), .ZN(n487) );
  NAND2_X1 U529 ( .A1(n474), .A2(n487), .ZN(n504) );
  NOR2_X1 U530 ( .A1(n491), .A2(n504), .ZN(n475) );
  XNOR2_X1 U531 ( .A(KEYINPUT101), .B(n475), .ZN(n485) );
  NOR2_X1 U532 ( .A1(n516), .A2(n485), .ZN(n477) );
  XNOR2_X1 U533 ( .A(KEYINPUT34), .B(KEYINPUT102), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U535 ( .A(G1GAT), .B(n478), .Z(G1324GAT) );
  NOR2_X1 U536 ( .A1(n518), .A2(n485), .ZN(n480) );
  XNOR2_X1 U537 ( .A(G8GAT), .B(KEYINPUT103), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n480), .B(n479), .ZN(G1325GAT) );
  NOR2_X1 U539 ( .A1(n485), .A2(n528), .ZN(n484) );
  XOR2_X1 U540 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n482) );
  XNOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n481) );
  XNOR2_X1 U542 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U544 ( .A1(n522), .A2(n485), .ZN(n486) );
  XOR2_X1 U545 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  NAND2_X1 U546 ( .A1(n579), .A2(n487), .ZN(n488) );
  NOR2_X1 U547 ( .A1(n534), .A2(n488), .ZN(n490) );
  XNOR2_X1 U548 ( .A(KEYINPUT37), .B(KEYINPUT106), .ZN(n489) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(n515) );
  NOR2_X1 U550 ( .A1(n515), .A2(n491), .ZN(n493) );
  XNOR2_X1 U551 ( .A(KEYINPUT107), .B(KEYINPUT38), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n500) );
  NOR2_X1 U553 ( .A1(n516), .A2(n500), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(KEYINPUT39), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G29GAT), .B(n495), .ZN(G1328GAT) );
  NOR2_X1 U556 ( .A1(n500), .A2(n518), .ZN(n496) );
  XOR2_X1 U557 ( .A(G36GAT), .B(n496), .Z(G1329GAT) );
  XNOR2_X1 U558 ( .A(KEYINPUT40), .B(KEYINPUT108), .ZN(n498) );
  NOR2_X1 U559 ( .A1(n528), .A2(n500), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U561 ( .A(G43GAT), .B(n499), .Z(G1330GAT) );
  NOR2_X1 U562 ( .A1(n500), .A2(n522), .ZN(n502) );
  XNOR2_X1 U563 ( .A(G50GAT), .B(KEYINPUT109), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(G1331GAT) );
  NAND2_X1 U565 ( .A1(n503), .A2(n558), .ZN(n514) );
  OR2_X1 U566 ( .A1(n504), .A2(n514), .ZN(n510) );
  NOR2_X1 U567 ( .A1(n516), .A2(n510), .ZN(n505) );
  XOR2_X1 U568 ( .A(n505), .B(KEYINPUT42), .Z(n506) );
  XNOR2_X1 U569 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U570 ( .A1(n518), .A2(n510), .ZN(n507) );
  XOR2_X1 U571 ( .A(KEYINPUT110), .B(n507), .Z(n508) );
  XNOR2_X1 U572 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U573 ( .A1(n528), .A2(n510), .ZN(n509) );
  XOR2_X1 U574 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U575 ( .A1(n522), .A2(n510), .ZN(n512) );
  XNOR2_X1 U576 ( .A(KEYINPUT111), .B(KEYINPUT43), .ZN(n511) );
  XNOR2_X1 U577 ( .A(n512), .B(n511), .ZN(n513) );
  XOR2_X1 U578 ( .A(G78GAT), .B(n513), .Z(G1335GAT) );
  OR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n521) );
  NOR2_X1 U580 ( .A1(n516), .A2(n521), .ZN(n517) );
  XOR2_X1 U581 ( .A(G85GAT), .B(n517), .Z(G1336GAT) );
  NOR2_X1 U582 ( .A1(n518), .A2(n521), .ZN(n519) );
  XOR2_X1 U583 ( .A(G92GAT), .B(n519), .Z(G1337GAT) );
  NOR2_X1 U584 ( .A1(n528), .A2(n521), .ZN(n520) );
  XOR2_X1 U585 ( .A(G99GAT), .B(n520), .Z(G1338GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n523) );
  XOR2_X1 U587 ( .A(KEYINPUT44), .B(n523), .Z(n524) );
  XNOR2_X1 U588 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n542) );
  OR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n529) );
  NOR2_X1 U591 ( .A1(n542), .A2(n529), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n556), .A2(n537), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G113GAT), .B(n530), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT113), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U595 ( .A1(n537), .A2(n558), .ZN(n531) );
  XNOR2_X1 U596 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  NAND2_X1 U598 ( .A1(n534), .A2(n537), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n535), .B(KEYINPUT50), .ZN(n536) );
  XNOR2_X1 U600 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT114), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U602 ( .A1(n537), .A2(n551), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT115), .Z(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n570), .A2(n542), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n552), .A2(n571), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n543), .ZN(G1344GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT53), .B(KEYINPUT117), .Z(n545) );
  XNOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n544) );
  XNOR2_X1 U611 ( .A(n545), .B(n544), .ZN(n546) );
  XOR2_X1 U612 ( .A(KEYINPUT116), .B(n546), .Z(n548) );
  NAND2_X1 U613 ( .A1(n552), .A2(n558), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n534), .A2(n552), .ZN(n550) );
  XNOR2_X1 U616 ( .A(n550), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT119), .Z(n554) );
  NAND2_X1 U618 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  NAND2_X1 U621 ( .A1(n563), .A2(n556), .ZN(n557) );
  XNOR2_X1 U622 ( .A(n557), .B(G169GAT), .ZN(G1348GAT) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n562) );
  NAND2_X1 U624 ( .A1(n563), .A2(n558), .ZN(n560) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(n562), .B(n561), .ZN(G1349GAT) );
  XOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT123), .Z(n565) );
  NAND2_X1 U629 ( .A1(n563), .A2(n534), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n565), .B(n564), .ZN(G1350GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n567) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(n568) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(n568), .Z(n573) );
  NOR2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n580) );
  NAND2_X1 U636 ( .A1(n580), .A2(n571), .ZN(n572) );
  XNOR2_X1 U637 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U639 ( .A1(n580), .A2(n574), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U642 ( .A1(n534), .A2(n580), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n582) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n583), .ZN(G1355GAT) );
endmodule

