

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U554 ( .A1(n739), .A2(n933), .ZN(n708) );
  NOR2_X2 U555 ( .A1(G164), .A2(G1384), .ZN(n695) );
  INV_X1 U556 ( .A(KEYINPUT98), .ZN(n722) );
  XNOR2_X1 U557 ( .A(n753), .B(KEYINPUT100), .ZN(n754) );
  XOR2_X1 U558 ( .A(KEYINPUT17), .B(n518), .Z(n865) );
  NOR2_X1 U559 ( .A1(G651), .A2(n620), .ZN(n635) );
  NOR2_X1 U560 ( .A1(n525), .A2(n524), .ZN(G164) );
  INV_X1 U561 ( .A(G2105), .ZN(n521) );
  NOR2_X2 U562 ( .A1(G2104), .A2(n521), .ZN(n869) );
  NAND2_X1 U563 ( .A1(n869), .A2(G126), .ZN(n517) );
  XNOR2_X1 U564 ( .A(n517), .B(KEYINPUT82), .ZN(n520) );
  NOR2_X1 U565 ( .A1(G2105), .A2(G2104), .ZN(n518) );
  NAND2_X1 U566 ( .A1(G138), .A2(n865), .ZN(n519) );
  NAND2_X1 U567 ( .A1(n520), .A2(n519), .ZN(n525) );
  AND2_X1 U568 ( .A1(n521), .A2(G2104), .ZN(n864) );
  NAND2_X1 U569 ( .A1(G102), .A2(n864), .ZN(n523) );
  AND2_X1 U570 ( .A1(G2105), .A2(G2104), .ZN(n872) );
  NAND2_X1 U571 ( .A1(G114), .A2(n872), .ZN(n522) );
  NAND2_X1 U572 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n620) );
  INV_X1 U574 ( .A(G651), .ZN(n529) );
  NOR2_X1 U575 ( .A1(n620), .A2(n529), .ZN(n631) );
  NAND2_X1 U576 ( .A1(n631), .A2(G78), .ZN(n528) );
  NOR2_X1 U577 ( .A1(G651), .A2(G543), .ZN(n526) );
  XNOR2_X1 U578 ( .A(n526), .B(KEYINPUT66), .ZN(n632) );
  NAND2_X1 U579 ( .A1(G91), .A2(n632), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n528), .A2(n527), .ZN(n534) );
  NAND2_X1 U581 ( .A1(G53), .A2(n635), .ZN(n532) );
  NOR2_X1 U582 ( .A1(G543), .A2(n529), .ZN(n530) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n530), .Z(n636) );
  NAND2_X1 U584 ( .A1(G65), .A2(n636), .ZN(n531) );
  NAND2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n533) );
  OR2_X1 U586 ( .A1(n534), .A2(n533), .ZN(G299) );
  NAND2_X1 U587 ( .A1(G52), .A2(n635), .ZN(n536) );
  NAND2_X1 U588 ( .A1(G64), .A2(n636), .ZN(n535) );
  NAND2_X1 U589 ( .A1(n536), .A2(n535), .ZN(n542) );
  NAND2_X1 U590 ( .A1(n631), .A2(G77), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G90), .A2(n632), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U593 ( .A(KEYINPUT68), .B(n539), .Z(n540) );
  XNOR2_X1 U594 ( .A(KEYINPUT9), .B(n540), .ZN(n541) );
  NOR2_X1 U595 ( .A1(n542), .A2(n541), .ZN(G171) );
  AND2_X1 U596 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U597 ( .A(G57), .ZN(G237) );
  NAND2_X1 U598 ( .A1(n872), .A2(G113), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G101), .A2(n864), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT23), .B(n543), .Z(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U602 ( .A1(G125), .A2(n869), .ZN(n547) );
  NAND2_X1 U603 ( .A1(G137), .A2(n865), .ZN(n546) );
  NAND2_X1 U604 ( .A1(n547), .A2(n546), .ZN(n548) );
  NOR2_X1 U605 ( .A1(n549), .A2(n548), .ZN(G160) );
  NAND2_X1 U606 ( .A1(G7), .A2(G661), .ZN(n550) );
  XNOR2_X1 U607 ( .A(n550), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U608 ( .A(G223), .ZN(n820) );
  NAND2_X1 U609 ( .A1(n820), .A2(G567), .ZN(n551) );
  XNOR2_X1 U610 ( .A(n551), .B(KEYINPUT71), .ZN(n552) );
  XNOR2_X1 U611 ( .A(KEYINPUT11), .B(n552), .ZN(G234) );
  NAND2_X1 U612 ( .A1(G81), .A2(n632), .ZN(n553) );
  XNOR2_X1 U613 ( .A(n553), .B(KEYINPUT12), .ZN(n555) );
  NAND2_X1 U614 ( .A1(G68), .A2(n631), .ZN(n554) );
  NAND2_X1 U615 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U616 ( .A(n556), .B(KEYINPUT13), .ZN(n558) );
  NAND2_X1 U617 ( .A1(G43), .A2(n635), .ZN(n557) );
  NAND2_X1 U618 ( .A1(n558), .A2(n557), .ZN(n561) );
  NAND2_X1 U619 ( .A1(n636), .A2(G56), .ZN(n559) );
  XOR2_X1 U620 ( .A(KEYINPUT14), .B(n559), .Z(n560) );
  NOR2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n975) );
  NAND2_X1 U622 ( .A1(n975), .A2(G860), .ZN(G153) );
  INV_X1 U623 ( .A(G171), .ZN(G301) );
  NAND2_X1 U624 ( .A1(G868), .A2(G301), .ZN(n571) );
  NAND2_X1 U625 ( .A1(n636), .A2(G66), .ZN(n568) );
  NAND2_X1 U626 ( .A1(G79), .A2(n631), .ZN(n563) );
  NAND2_X1 U627 ( .A1(G54), .A2(n635), .ZN(n562) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U629 ( .A1(n632), .A2(G92), .ZN(n564) );
  XOR2_X1 U630 ( .A(KEYINPUT72), .B(n564), .Z(n565) );
  NOR2_X1 U631 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT15), .B(n569), .Z(n954) );
  INV_X1 U634 ( .A(G868), .ZN(n651) );
  NAND2_X1 U635 ( .A1(n954), .A2(n651), .ZN(n570) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(G284) );
  NAND2_X1 U637 ( .A1(G89), .A2(n632), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(KEYINPUT4), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G76), .A2(n631), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n575), .B(KEYINPUT5), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G51), .A2(n635), .ZN(n577) );
  NAND2_X1 U643 ( .A1(G63), .A2(n636), .ZN(n576) );
  NAND2_X1 U644 ( .A1(n577), .A2(n576), .ZN(n578) );
  XOR2_X1 U645 ( .A(KEYINPUT6), .B(n578), .Z(n579) );
  NAND2_X1 U646 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U647 ( .A(n581), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U648 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NOR2_X1 U649 ( .A1(G286), .A2(n651), .ZN(n583) );
  NOR2_X1 U650 ( .A1(G868), .A2(G299), .ZN(n582) );
  NOR2_X1 U651 ( .A1(n583), .A2(n582), .ZN(G297) );
  INV_X1 U652 ( .A(G860), .ZN(n584) );
  NAND2_X1 U653 ( .A1(n584), .A2(G559), .ZN(n585) );
  INV_X1 U654 ( .A(n954), .ZN(n607) );
  NAND2_X1 U655 ( .A1(n585), .A2(n607), .ZN(n586) );
  XNOR2_X1 U656 ( .A(n586), .B(KEYINPUT73), .ZN(n587) );
  XOR2_X1 U657 ( .A(KEYINPUT16), .B(n587), .Z(G148) );
  NAND2_X1 U658 ( .A1(n607), .A2(G868), .ZN(n588) );
  NOR2_X1 U659 ( .A1(G559), .A2(n588), .ZN(n590) );
  AND2_X1 U660 ( .A1(n651), .A2(n975), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(G282) );
  NAND2_X1 U662 ( .A1(G99), .A2(n864), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G111), .A2(n872), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n592), .A2(n591), .ZN(n593) );
  XNOR2_X1 U665 ( .A(KEYINPUT74), .B(n593), .ZN(n598) );
  NAND2_X1 U666 ( .A1(n869), .A2(G123), .ZN(n594) );
  XNOR2_X1 U667 ( .A(n594), .B(KEYINPUT18), .ZN(n596) );
  NAND2_X1 U668 ( .A1(G135), .A2(n865), .ZN(n595) );
  NAND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n597) );
  NOR2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n903) );
  XNOR2_X1 U671 ( .A(n903), .B(G2096), .ZN(n600) );
  INV_X1 U672 ( .A(G2100), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(G156) );
  NAND2_X1 U674 ( .A1(n631), .A2(G80), .ZN(n602) );
  NAND2_X1 U675 ( .A1(G93), .A2(n632), .ZN(n601) );
  NAND2_X1 U676 ( .A1(n602), .A2(n601), .ZN(n606) );
  NAND2_X1 U677 ( .A1(G55), .A2(n635), .ZN(n604) );
  NAND2_X1 U678 ( .A1(G67), .A2(n636), .ZN(n603) );
  NAND2_X1 U679 ( .A1(n604), .A2(n603), .ZN(n605) );
  OR2_X1 U680 ( .A1(n606), .A2(n605), .ZN(n652) );
  NAND2_X1 U681 ( .A1(G559), .A2(n607), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(n975), .ZN(n649) );
  XNOR2_X1 U683 ( .A(KEYINPUT75), .B(n649), .ZN(n609) );
  NOR2_X1 U684 ( .A1(G860), .A2(n609), .ZN(n610) );
  XOR2_X1 U685 ( .A(n652), .B(n610), .Z(G145) );
  NAND2_X1 U686 ( .A1(n631), .A2(G75), .ZN(n612) );
  NAND2_X1 U687 ( .A1(G88), .A2(n632), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G50), .A2(n635), .ZN(n614) );
  NAND2_X1 U690 ( .A1(G62), .A2(n636), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n616), .A2(n615), .ZN(G166) );
  NAND2_X1 U693 ( .A1(G49), .A2(n635), .ZN(n618) );
  NAND2_X1 U694 ( .A1(G74), .A2(G651), .ZN(n617) );
  NAND2_X1 U695 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U696 ( .A1(n636), .A2(n619), .ZN(n622) );
  NAND2_X1 U697 ( .A1(n620), .A2(G87), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(G288) );
  NAND2_X1 U699 ( .A1(n636), .A2(G61), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G86), .A2(n632), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U702 ( .A1(n631), .A2(G73), .ZN(n625) );
  XOR2_X1 U703 ( .A(KEYINPUT2), .B(n625), .Z(n626) );
  NOR2_X1 U704 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT76), .ZN(n630) );
  NAND2_X1 U706 ( .A1(G48), .A2(n635), .ZN(n629) );
  NAND2_X1 U707 ( .A1(n630), .A2(n629), .ZN(G305) );
  NAND2_X1 U708 ( .A1(n631), .A2(G72), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G85), .A2(n632), .ZN(n633) );
  NAND2_X1 U710 ( .A1(n634), .A2(n633), .ZN(n640) );
  NAND2_X1 U711 ( .A1(G47), .A2(n635), .ZN(n638) );
  NAND2_X1 U712 ( .A1(G60), .A2(n636), .ZN(n637) );
  NAND2_X1 U713 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U714 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U715 ( .A(KEYINPUT67), .B(n641), .ZN(G290) );
  XOR2_X1 U716 ( .A(KEYINPUT78), .B(KEYINPUT77), .Z(n643) );
  XNOR2_X1 U717 ( .A(G166), .B(KEYINPUT19), .ZN(n642) );
  XNOR2_X1 U718 ( .A(n643), .B(n642), .ZN(n646) );
  XOR2_X1 U719 ( .A(G299), .B(G305), .Z(n644) );
  XNOR2_X1 U720 ( .A(G288), .B(n644), .ZN(n645) );
  XNOR2_X1 U721 ( .A(n646), .B(n645), .ZN(n648) );
  XOR2_X1 U722 ( .A(G290), .B(n652), .Z(n647) );
  XNOR2_X1 U723 ( .A(n648), .B(n647), .ZN(n887) );
  XOR2_X1 U724 ( .A(n887), .B(n649), .Z(n650) );
  NOR2_X1 U725 ( .A1(n651), .A2(n650), .ZN(n654) );
  NOR2_X1 U726 ( .A1(G868), .A2(n652), .ZN(n653) );
  NOR2_X1 U727 ( .A1(n654), .A2(n653), .ZN(G295) );
  NAND2_X1 U728 ( .A1(G2078), .A2(G2084), .ZN(n655) );
  XOR2_X1 U729 ( .A(KEYINPUT20), .B(n655), .Z(n656) );
  NAND2_X1 U730 ( .A1(G2090), .A2(n656), .ZN(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT21), .B(n657), .ZN(n658) );
  NAND2_X1 U732 ( .A1(n658), .A2(G2072), .ZN(G158) );
  XOR2_X1 U733 ( .A(KEYINPUT79), .B(G44), .Z(n659) );
  XNOR2_X1 U734 ( .A(KEYINPUT3), .B(n659), .ZN(G218) );
  XOR2_X1 U735 ( .A(KEYINPUT70), .B(G82), .Z(G220) );
  XNOR2_X1 U736 ( .A(KEYINPUT69), .B(G132), .ZN(G219) );
  NOR2_X1 U737 ( .A1(G220), .A2(G219), .ZN(n660) );
  XOR2_X1 U738 ( .A(KEYINPUT22), .B(n660), .Z(n661) );
  XNOR2_X1 U739 ( .A(n661), .B(KEYINPUT80), .ZN(n662) );
  NOR2_X1 U740 ( .A1(G218), .A2(n662), .ZN(n663) );
  NAND2_X1 U741 ( .A1(G96), .A2(n663), .ZN(n824) );
  NAND2_X1 U742 ( .A1(G2106), .A2(n824), .ZN(n667) );
  NAND2_X1 U743 ( .A1(G108), .A2(G120), .ZN(n664) );
  NOR2_X1 U744 ( .A1(G237), .A2(n664), .ZN(n665) );
  NAND2_X1 U745 ( .A1(G69), .A2(n665), .ZN(n825) );
  NAND2_X1 U746 ( .A1(G567), .A2(n825), .ZN(n666) );
  NAND2_X1 U747 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U748 ( .A(KEYINPUT81), .B(n668), .ZN(G319) );
  INV_X1 U749 ( .A(G319), .ZN(n670) );
  NAND2_X1 U750 ( .A1(G661), .A2(G483), .ZN(n669) );
  NOR2_X1 U751 ( .A1(n670), .A2(n669), .ZN(n823) );
  NAND2_X1 U752 ( .A1(n823), .A2(G36), .ZN(G176) );
  XNOR2_X1 U753 ( .A(KEYINPUT83), .B(G166), .ZN(G303) );
  XNOR2_X1 U754 ( .A(KEYINPUT104), .B(KEYINPUT40), .ZN(n808) );
  NAND2_X1 U755 ( .A1(G117), .A2(n872), .ZN(n677) );
  NAND2_X1 U756 ( .A1(G129), .A2(n869), .ZN(n672) );
  NAND2_X1 U757 ( .A1(G141), .A2(n865), .ZN(n671) );
  NAND2_X1 U758 ( .A1(n672), .A2(n671), .ZN(n675) );
  NAND2_X1 U759 ( .A1(n864), .A2(G105), .ZN(n673) );
  XOR2_X1 U760 ( .A(KEYINPUT38), .B(n673), .Z(n674) );
  NOR2_X1 U761 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U762 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U763 ( .A(n678), .B(KEYINPUT90), .ZN(n882) );
  NAND2_X1 U764 ( .A1(G1996), .A2(n882), .ZN(n688) );
  NAND2_X1 U765 ( .A1(n869), .A2(G119), .ZN(n679) );
  XNOR2_X1 U766 ( .A(n679), .B(KEYINPUT88), .ZN(n681) );
  NAND2_X1 U767 ( .A1(G107), .A2(n872), .ZN(n680) );
  NAND2_X1 U768 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U769 ( .A(KEYINPUT89), .B(n682), .ZN(n686) );
  NAND2_X1 U770 ( .A1(G95), .A2(n864), .ZN(n684) );
  NAND2_X1 U771 ( .A1(G131), .A2(n865), .ZN(n683) );
  AND2_X1 U772 ( .A1(n684), .A2(n683), .ZN(n685) );
  NAND2_X1 U773 ( .A1(n686), .A2(n685), .ZN(n863) );
  NAND2_X1 U774 ( .A1(G1991), .A2(n863), .ZN(n687) );
  NAND2_X1 U775 ( .A1(n688), .A2(n687), .ZN(n922) );
  NAND2_X1 U776 ( .A1(G160), .A2(G40), .ZN(n693) );
  NOR2_X1 U777 ( .A1(n695), .A2(n693), .ZN(n804) );
  NAND2_X1 U778 ( .A1(n922), .A2(n804), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n689), .B(KEYINPUT91), .ZN(n794) );
  XOR2_X1 U780 ( .A(KEYINPUT92), .B(n794), .Z(n692) );
  XNOR2_X1 U781 ( .A(G1986), .B(G290), .ZN(n966) );
  NAND2_X1 U782 ( .A1(n966), .A2(n804), .ZN(n690) );
  XNOR2_X1 U783 ( .A(n690), .B(KEYINPUT84), .ZN(n691) );
  NAND2_X1 U784 ( .A1(n692), .A2(n691), .ZN(n778) );
  INV_X1 U785 ( .A(n693), .ZN(n694) );
  NAND2_X2 U786 ( .A1(n695), .A2(n694), .ZN(n739) );
  NAND2_X1 U787 ( .A1(G8), .A2(n739), .ZN(n773) );
  NOR2_X1 U788 ( .A1(G1966), .A2(n773), .ZN(n749) );
  NOR2_X1 U789 ( .A1(G2084), .A2(n739), .ZN(n750) );
  NOR2_X1 U790 ( .A1(n749), .A2(n750), .ZN(n696) );
  NAND2_X1 U791 ( .A1(G8), .A2(n696), .ZN(n697) );
  XNOR2_X1 U792 ( .A(KEYINPUT30), .B(n697), .ZN(n698) );
  NOR2_X1 U793 ( .A1(G168), .A2(n698), .ZN(n704) );
  INV_X1 U794 ( .A(n739), .ZN(n718) );
  NOR2_X1 U795 ( .A1(n718), .A2(G1961), .ZN(n699) );
  XOR2_X1 U796 ( .A(KEYINPUT94), .B(n699), .Z(n701) );
  XNOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .ZN(n939) );
  NAND2_X1 U798 ( .A1(n718), .A2(n939), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n701), .A2(n700), .ZN(n734) );
  NOR2_X1 U800 ( .A1(G171), .A2(n734), .ZN(n702) );
  XOR2_X1 U801 ( .A(KEYINPUT99), .B(n702), .Z(n703) );
  NOR2_X1 U802 ( .A1(n704), .A2(n703), .ZN(n705) );
  XOR2_X1 U803 ( .A(KEYINPUT31), .B(n705), .Z(n738) );
  XNOR2_X1 U804 ( .A(G1996), .B(KEYINPUT95), .ZN(n933) );
  XOR2_X1 U805 ( .A(KEYINPUT26), .B(KEYINPUT96), .Z(n706) );
  XNOR2_X1 U806 ( .A(KEYINPUT64), .B(n706), .ZN(n707) );
  XNOR2_X1 U807 ( .A(n708), .B(n707), .ZN(n710) );
  NAND2_X1 U808 ( .A1(n739), .A2(G1341), .ZN(n709) );
  NAND2_X1 U809 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U810 ( .A(KEYINPUT97), .B(n711), .ZN(n712) );
  NAND2_X1 U811 ( .A1(n712), .A2(n975), .ZN(n713) );
  XNOR2_X1 U812 ( .A(n713), .B(KEYINPUT65), .ZN(n717) );
  NOR2_X1 U813 ( .A1(n718), .A2(G1348), .ZN(n715) );
  NOR2_X1 U814 ( .A1(G2067), .A2(n739), .ZN(n714) );
  NOR2_X1 U815 ( .A1(n715), .A2(n714), .ZN(n726) );
  NAND2_X1 U816 ( .A1(n726), .A2(n954), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n717), .A2(n716), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n718), .A2(G2072), .ZN(n719) );
  XOR2_X1 U819 ( .A(KEYINPUT27), .B(n719), .Z(n721) );
  NAND2_X1 U820 ( .A1(G1956), .A2(n739), .ZN(n720) );
  NAND2_X1 U821 ( .A1(n721), .A2(n720), .ZN(n729) );
  NOR2_X1 U822 ( .A1(G299), .A2(n729), .ZN(n723) );
  XNOR2_X1 U823 ( .A(n723), .B(n722), .ZN(n724) );
  NAND2_X1 U824 ( .A1(n725), .A2(n724), .ZN(n728) );
  NOR2_X1 U825 ( .A1(n726), .A2(n954), .ZN(n727) );
  NOR2_X1 U826 ( .A1(n728), .A2(n727), .ZN(n732) );
  NAND2_X1 U827 ( .A1(G299), .A2(n729), .ZN(n730) );
  XOR2_X1 U828 ( .A(KEYINPUT28), .B(n730), .Z(n731) );
  NOR2_X1 U829 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U830 ( .A(n733), .B(KEYINPUT29), .ZN(n736) );
  NAND2_X1 U831 ( .A1(G171), .A2(n734), .ZN(n735) );
  NAND2_X1 U832 ( .A1(n736), .A2(n735), .ZN(n737) );
  NAND2_X1 U833 ( .A1(n738), .A2(n737), .ZN(n747) );
  NAND2_X1 U834 ( .A1(G286), .A2(n747), .ZN(n744) );
  NOR2_X1 U835 ( .A1(G1971), .A2(n773), .ZN(n741) );
  NOR2_X1 U836 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U837 ( .A1(n741), .A2(n740), .ZN(n742) );
  NAND2_X1 U838 ( .A1(n742), .A2(G303), .ZN(n743) );
  NAND2_X1 U839 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U840 ( .A1(n745), .A2(G8), .ZN(n746) );
  XNOR2_X1 U841 ( .A(KEYINPUT32), .B(n746), .ZN(n755) );
  INV_X1 U842 ( .A(n747), .ZN(n748) );
  NOR2_X1 U843 ( .A1(n749), .A2(n748), .ZN(n752) );
  NAND2_X1 U844 ( .A1(G8), .A2(n750), .ZN(n751) );
  NAND2_X1 U845 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U846 ( .A1(n755), .A2(n754), .ZN(n767) );
  NOR2_X1 U847 ( .A1(G1976), .A2(G288), .ZN(n961) );
  NOR2_X1 U848 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NOR2_X1 U849 ( .A1(n961), .A2(n960), .ZN(n756) );
  NAND2_X1 U850 ( .A1(n767), .A2(n756), .ZN(n757) );
  NAND2_X1 U851 ( .A1(G1976), .A2(G288), .ZN(n963) );
  NAND2_X1 U852 ( .A1(n757), .A2(n963), .ZN(n758) );
  NOR2_X1 U853 ( .A1(n773), .A2(n758), .ZN(n759) );
  NOR2_X1 U854 ( .A1(KEYINPUT33), .A2(n759), .ZN(n762) );
  NAND2_X1 U855 ( .A1(n961), .A2(KEYINPUT33), .ZN(n760) );
  NOR2_X1 U856 ( .A1(n760), .A2(n773), .ZN(n761) );
  NOR2_X1 U857 ( .A1(n762), .A2(n761), .ZN(n763) );
  XOR2_X1 U858 ( .A(G1981), .B(G305), .Z(n971) );
  NAND2_X1 U859 ( .A1(n763), .A2(n971), .ZN(n770) );
  NOR2_X1 U860 ( .A1(G2090), .A2(G303), .ZN(n764) );
  NAND2_X1 U861 ( .A1(G8), .A2(n764), .ZN(n765) );
  XOR2_X1 U862 ( .A(KEYINPUT101), .B(n765), .Z(n766) );
  NAND2_X1 U863 ( .A1(n767), .A2(n766), .ZN(n768) );
  NAND2_X1 U864 ( .A1(n768), .A2(n773), .ZN(n769) );
  NAND2_X1 U865 ( .A1(n770), .A2(n769), .ZN(n776) );
  NOR2_X1 U866 ( .A1(G1981), .A2(G305), .ZN(n771) );
  XNOR2_X1 U867 ( .A(n771), .B(KEYINPUT24), .ZN(n772) );
  XNOR2_X1 U868 ( .A(n772), .B(KEYINPUT93), .ZN(n774) );
  NOR2_X1 U869 ( .A1(n774), .A2(n773), .ZN(n775) );
  NOR2_X1 U870 ( .A1(n776), .A2(n775), .ZN(n777) );
  NOR2_X1 U871 ( .A1(n778), .A2(n777), .ZN(n791) );
  XNOR2_X1 U872 ( .A(KEYINPUT37), .B(G2067), .ZN(n800) );
  XNOR2_X1 U873 ( .A(KEYINPUT87), .B(KEYINPUT35), .ZN(n782) );
  NAND2_X1 U874 ( .A1(G128), .A2(n869), .ZN(n780) );
  NAND2_X1 U875 ( .A1(G116), .A2(n872), .ZN(n779) );
  NAND2_X1 U876 ( .A1(n780), .A2(n779), .ZN(n781) );
  XNOR2_X1 U877 ( .A(n782), .B(n781), .ZN(n789) );
  XNOR2_X1 U878 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n783) );
  XNOR2_X1 U879 ( .A(n783), .B(KEYINPUT34), .ZN(n787) );
  NAND2_X1 U880 ( .A1(G104), .A2(n864), .ZN(n785) );
  NAND2_X1 U881 ( .A1(G140), .A2(n865), .ZN(n784) );
  NAND2_X1 U882 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U883 ( .A(n787), .B(n786), .Z(n788) );
  NOR2_X1 U884 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U885 ( .A(KEYINPUT36), .B(n790), .ZN(n883) );
  NOR2_X1 U886 ( .A1(n800), .A2(n883), .ZN(n905) );
  NAND2_X1 U887 ( .A1(n804), .A2(n905), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n791), .A2(n798), .ZN(n806) );
  NOR2_X1 U889 ( .A1(G1991), .A2(n863), .ZN(n904) );
  NOR2_X1 U890 ( .A1(G1986), .A2(G290), .ZN(n792) );
  NOR2_X1 U891 ( .A1(n904), .A2(n792), .ZN(n793) );
  NOR2_X1 U892 ( .A1(n794), .A2(n793), .ZN(n796) );
  NOR2_X1 U893 ( .A1(n882), .A2(G1996), .ZN(n795) );
  XNOR2_X1 U894 ( .A(n795), .B(KEYINPUT102), .ZN(n914) );
  NOR2_X1 U895 ( .A1(n796), .A2(n914), .ZN(n797) );
  XNOR2_X1 U896 ( .A(n797), .B(KEYINPUT39), .ZN(n799) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n801) );
  NAND2_X1 U898 ( .A1(n800), .A2(n883), .ZN(n920) );
  NAND2_X1 U899 ( .A1(n801), .A2(n920), .ZN(n802) );
  XOR2_X1 U900 ( .A(KEYINPUT103), .B(n802), .Z(n803) );
  NAND2_X1 U901 ( .A1(n804), .A2(n803), .ZN(n805) );
  NAND2_X1 U902 ( .A1(n806), .A2(n805), .ZN(n807) );
  XNOR2_X1 U903 ( .A(n808), .B(n807), .ZN(G329) );
  XNOR2_X1 U904 ( .A(G2443), .B(G2446), .ZN(n818) );
  XOR2_X1 U905 ( .A(G2430), .B(KEYINPUT106), .Z(n810) );
  XNOR2_X1 U906 ( .A(G2454), .B(G2435), .ZN(n809) );
  XNOR2_X1 U907 ( .A(n810), .B(n809), .ZN(n814) );
  XOR2_X1 U908 ( .A(G2438), .B(G2427), .Z(n812) );
  XNOR2_X1 U909 ( .A(G1348), .B(G1341), .ZN(n811) );
  XNOR2_X1 U910 ( .A(n812), .B(n811), .ZN(n813) );
  XOR2_X1 U911 ( .A(n814), .B(n813), .Z(n816) );
  XNOR2_X1 U912 ( .A(G2451), .B(KEYINPUT105), .ZN(n815) );
  XNOR2_X1 U913 ( .A(n816), .B(n815), .ZN(n817) );
  XNOR2_X1 U914 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n819), .A2(G14), .ZN(n896) );
  XNOR2_X1 U916 ( .A(KEYINPUT107), .B(n896), .ZN(G401) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n820), .ZN(G217) );
  AND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n821) );
  NAND2_X1 U919 ( .A1(G661), .A2(n821), .ZN(G259) );
  NAND2_X1 U920 ( .A1(G3), .A2(G1), .ZN(n822) );
  NAND2_X1 U921 ( .A1(n823), .A2(n822), .ZN(G188) );
  XOR2_X1 U922 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  NOR2_X1 U925 ( .A1(n825), .A2(n824), .ZN(G325) );
  INV_X1 U926 ( .A(G325), .ZN(G261) );
  XOR2_X1 U927 ( .A(G2100), .B(G2096), .Z(n827) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(G2678), .ZN(n826) );
  XNOR2_X1 U929 ( .A(n827), .B(n826), .ZN(n831) );
  XOR2_X1 U930 ( .A(KEYINPUT43), .B(G2090), .Z(n829) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n828) );
  XNOR2_X1 U932 ( .A(n829), .B(n828), .ZN(n830) );
  XOR2_X1 U933 ( .A(n831), .B(n830), .Z(n833) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n832) );
  XNOR2_X1 U935 ( .A(n833), .B(n832), .ZN(G227) );
  XOR2_X1 U936 ( .A(G1976), .B(G1971), .Z(n835) );
  XNOR2_X1 U937 ( .A(G1986), .B(G1956), .ZN(n834) );
  XNOR2_X1 U938 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U939 ( .A(n836), .B(G2474), .Z(n838) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n837) );
  XNOR2_X1 U941 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U942 ( .A(KEYINPUT41), .B(G1981), .Z(n840) );
  XNOR2_X1 U943 ( .A(G1966), .B(G1961), .ZN(n839) );
  XNOR2_X1 U944 ( .A(n840), .B(n839), .ZN(n841) );
  XNOR2_X1 U945 ( .A(n842), .B(n841), .ZN(G229) );
  NAND2_X1 U946 ( .A1(G100), .A2(n864), .ZN(n844) );
  NAND2_X1 U947 ( .A1(G112), .A2(n872), .ZN(n843) );
  NAND2_X1 U948 ( .A1(n844), .A2(n843), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n845), .B(KEYINPUT109), .ZN(n847) );
  NAND2_X1 U950 ( .A1(G136), .A2(n865), .ZN(n846) );
  NAND2_X1 U951 ( .A1(n847), .A2(n846), .ZN(n850) );
  NAND2_X1 U952 ( .A1(n869), .A2(G124), .ZN(n848) );
  XOR2_X1 U953 ( .A(KEYINPUT44), .B(n848), .Z(n849) );
  NOR2_X1 U954 ( .A1(n850), .A2(n849), .ZN(G162) );
  XOR2_X1 U955 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n852) );
  XNOR2_X1 U956 ( .A(G160), .B(KEYINPUT113), .ZN(n851) );
  XNOR2_X1 U957 ( .A(n852), .B(n851), .ZN(n881) );
  NAND2_X1 U958 ( .A1(n864), .A2(G103), .ZN(n853) );
  XNOR2_X1 U959 ( .A(KEYINPUT111), .B(n853), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G127), .A2(n869), .ZN(n855) );
  NAND2_X1 U961 ( .A1(G115), .A2(n872), .ZN(n854) );
  NAND2_X1 U962 ( .A1(n855), .A2(n854), .ZN(n856) );
  XNOR2_X1 U963 ( .A(n856), .B(KEYINPUT47), .ZN(n857) );
  XNOR2_X1 U964 ( .A(n857), .B(KEYINPUT112), .ZN(n859) );
  NAND2_X1 U965 ( .A1(n865), .A2(G139), .ZN(n858) );
  NAND2_X1 U966 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U967 ( .A1(n861), .A2(n860), .ZN(n909) );
  XOR2_X1 U968 ( .A(n909), .B(G162), .Z(n862) );
  XNOR2_X1 U969 ( .A(n863), .B(n862), .ZN(n877) );
  NAND2_X1 U970 ( .A1(G106), .A2(n864), .ZN(n867) );
  NAND2_X1 U971 ( .A1(G142), .A2(n865), .ZN(n866) );
  NAND2_X1 U972 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U973 ( .A(n868), .B(KEYINPUT45), .ZN(n871) );
  NAND2_X1 U974 ( .A1(G130), .A2(n869), .ZN(n870) );
  NAND2_X1 U975 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n872), .A2(G118), .ZN(n873) );
  XOR2_X1 U977 ( .A(KEYINPUT110), .B(n873), .Z(n874) );
  NOR2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U979 ( .A(n877), .B(n876), .Z(n879) );
  XNOR2_X1 U980 ( .A(G164), .B(n903), .ZN(n878) );
  XNOR2_X1 U981 ( .A(n879), .B(n878), .ZN(n880) );
  XNOR2_X1 U982 ( .A(n881), .B(n880), .ZN(n885) );
  XNOR2_X1 U983 ( .A(n883), .B(n882), .ZN(n884) );
  XNOR2_X1 U984 ( .A(n885), .B(n884), .ZN(n886) );
  NOR2_X1 U985 ( .A1(G37), .A2(n886), .ZN(G395) );
  XNOR2_X1 U986 ( .A(n975), .B(G286), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n888), .B(n887), .ZN(n893) );
  XNOR2_X1 U988 ( .A(KEYINPUT115), .B(KEYINPUT114), .ZN(n890) );
  XNOR2_X1 U989 ( .A(n954), .B(KEYINPUT116), .ZN(n889) );
  XNOR2_X1 U990 ( .A(n890), .B(n889), .ZN(n891) );
  XOR2_X1 U991 ( .A(G301), .B(n891), .Z(n892) );
  XNOR2_X1 U992 ( .A(n893), .B(n892), .ZN(n894) );
  NOR2_X1 U993 ( .A1(G37), .A2(n894), .ZN(n895) );
  XOR2_X1 U994 ( .A(KEYINPUT117), .B(n895), .Z(G397) );
  NAND2_X1 U995 ( .A1(G319), .A2(n896), .ZN(n899) );
  NOR2_X1 U996 ( .A1(G227), .A2(G229), .ZN(n897) );
  XNOR2_X1 U997 ( .A(KEYINPUT49), .B(n897), .ZN(n898) );
  NOR2_X1 U998 ( .A1(n899), .A2(n898), .ZN(n901) );
  NOR2_X1 U999 ( .A1(G395), .A2(G397), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(n901), .A2(n900), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  INV_X1 U1002 ( .A(G96), .ZN(G221) );
  INV_X1 U1003 ( .A(G69), .ZN(G235) );
  XOR2_X1 U1004 ( .A(G2084), .B(G160), .Z(n902) );
  NOR2_X1 U1005 ( .A1(n903), .A2(n902), .ZN(n907) );
  NOR2_X1 U1006 ( .A1(n905), .A2(n904), .ZN(n906) );
  NAND2_X1 U1007 ( .A1(n907), .A2(n906), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(KEYINPUT118), .B(n908), .ZN(n919) );
  XOR2_X1 U1009 ( .A(G2072), .B(n909), .Z(n911) );
  XOR2_X1 U1010 ( .A(G164), .B(G2078), .Z(n910) );
  NOR2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT50), .B(n912), .ZN(n917) );
  XOR2_X1 U1013 ( .A(G2090), .B(G162), .Z(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n915) );
  XOR2_X1 U1015 ( .A(KEYINPUT51), .B(n915), .Z(n916) );
  NAND2_X1 U1016 ( .A1(n917), .A2(n916), .ZN(n918) );
  NOR2_X1 U1017 ( .A1(n919), .A2(n918), .ZN(n924) );
  INV_X1 U1018 ( .A(n920), .ZN(n921) );
  NOR2_X1 U1019 ( .A1(n922), .A2(n921), .ZN(n923) );
  NAND2_X1 U1020 ( .A1(n924), .A2(n923), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(KEYINPUT52), .B(n925), .ZN(n926) );
  XNOR2_X1 U1022 ( .A(KEYINPUT119), .B(n926), .ZN(n927) );
  XOR2_X1 U1023 ( .A(KEYINPUT55), .B(KEYINPUT120), .Z(n950) );
  NAND2_X1 U1024 ( .A1(n927), .A2(n950), .ZN(n928) );
  NAND2_X1 U1025 ( .A1(n928), .A2(G29), .ZN(n929) );
  XOR2_X1 U1026 ( .A(KEYINPUT121), .B(n929), .Z(n1010) );
  XNOR2_X1 U1027 ( .A(G1991), .B(G25), .ZN(n931) );
  XNOR2_X1 U1028 ( .A(G33), .B(G2072), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n938) );
  XOR2_X1 U1030 ( .A(G2067), .B(G26), .Z(n932) );
  NAND2_X1 U1031 ( .A1(n932), .A2(G28), .ZN(n936) );
  XOR2_X1 U1032 ( .A(G32), .B(n933), .Z(n934) );
  XNOR2_X1 U1033 ( .A(KEYINPUT122), .B(n934), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n941) );
  XOR2_X1 U1036 ( .A(G27), .B(n939), .Z(n940) );
  NOR2_X1 U1037 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1038 ( .A(n942), .B(KEYINPUT53), .ZN(n943) );
  XNOR2_X1 U1039 ( .A(n943), .B(KEYINPUT123), .ZN(n946) );
  XOR2_X1 U1040 ( .A(G2084), .B(G34), .Z(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT54), .B(n944), .ZN(n945) );
  NAND2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n948) );
  XNOR2_X1 U1043 ( .A(G35), .B(G2090), .ZN(n947) );
  NOR2_X1 U1044 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1045 ( .A(n950), .B(n949), .Z(n952) );
  INV_X1 U1046 ( .A(G29), .ZN(n951) );
  NAND2_X1 U1047 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1048 ( .A1(n953), .A2(G11), .ZN(n1008) );
  XNOR2_X1 U1049 ( .A(G16), .B(KEYINPUT56), .ZN(n981) );
  XNOR2_X1 U1050 ( .A(n954), .B(G1348), .ZN(n956) );
  XNOR2_X1 U1051 ( .A(G299), .B(G1956), .ZN(n955) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(G1971), .A2(G303), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n970) );
  XOR2_X1 U1055 ( .A(G1961), .B(G171), .Z(n959) );
  NOR2_X1 U1056 ( .A1(n960), .A2(n959), .ZN(n968) );
  INV_X1 U1057 ( .A(n961), .ZN(n962) );
  NAND2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1059 ( .A(KEYINPUT125), .B(n964), .Z(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n979) );
  XNOR2_X1 U1063 ( .A(G1966), .B(G168), .ZN(n972) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n973), .B(KEYINPUT57), .ZN(n974) );
  XOR2_X1 U1066 ( .A(KEYINPUT124), .B(n974), .Z(n977) );
  XOR2_X1 U1067 ( .A(n975), .B(G1341), .Z(n976) );
  NOR2_X1 U1068 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1069 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n981), .A2(n980), .ZN(n1006) );
  INV_X1 U1071 ( .A(G16), .ZN(n1004) );
  XOR2_X1 U1072 ( .A(G1348), .B(KEYINPUT59), .Z(n982) );
  XNOR2_X1 U1073 ( .A(G4), .B(n982), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G20), .B(G1956), .ZN(n983) );
  NOR2_X1 U1075 ( .A1(n984), .A2(n983), .ZN(n988) );
  XNOR2_X1 U1076 ( .A(G1341), .B(G19), .ZN(n986) );
  XNOR2_X1 U1077 ( .A(G6), .B(G1981), .ZN(n985) );
  NOR2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1079 ( .A1(n988), .A2(n987), .ZN(n989) );
  XOR2_X1 U1080 ( .A(KEYINPUT126), .B(n989), .Z(n990) );
  XNOR2_X1 U1081 ( .A(KEYINPUT60), .B(n990), .ZN(n994) );
  XNOR2_X1 U1082 ( .A(G1966), .B(G21), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(G5), .B(G1961), .ZN(n991) );
  NOR2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n1001) );
  XNOR2_X1 U1086 ( .A(G1971), .B(G22), .ZN(n996) );
  XNOR2_X1 U1087 ( .A(G23), .B(G1976), .ZN(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n998) );
  XOR2_X1 U1089 ( .A(G1986), .B(G24), .Z(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1091 ( .A(KEYINPUT58), .B(n999), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(KEYINPUT61), .B(n1002), .ZN(n1003) );
  NAND2_X1 U1094 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1095 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1097 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1011), .Z(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

