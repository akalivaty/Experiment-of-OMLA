//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 0 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:26 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n714, new_n715, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021;
  INV_X1    g000(.A(KEYINPUT89), .ZN(new_n187));
  XNOR2_X1  g001(.A(G113), .B(G122), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n188), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G125), .ZN(new_n191));
  NOR3_X1   g005(.A1(new_n191), .A2(KEYINPUT16), .A3(G140), .ZN(new_n192));
  XNOR2_X1  g006(.A(G125), .B(G140), .ZN(new_n193));
  AOI21_X1  g007(.A(new_n192), .B1(new_n193), .B2(KEYINPUT16), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n191), .A2(G140), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT19), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT19), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n193), .A2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n200), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g018(.A1(G237), .A2(G953), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n205), .A2(G143), .A3(G214), .ZN(new_n206));
  INV_X1    g020(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(G143), .B1(new_n205), .B2(G214), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n207), .A2(new_n208), .A3(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n205), .A2(G214), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n210), .B1(new_n213), .B2(new_n206), .ZN(new_n214));
  OAI211_X1 g028(.A(new_n195), .B(new_n204), .C1(new_n209), .C2(new_n214), .ZN(new_n215));
  OAI211_X1 g029(.A(KEYINPUT18), .B(G131), .C1(new_n207), .C2(new_n208), .ZN(new_n216));
  NAND2_X1  g030(.A1(KEYINPUT18), .A2(G131), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n213), .A2(new_n206), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n199), .A2(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n193), .A2(new_n203), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n216), .A2(new_n218), .A3(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n190), .B1(new_n215), .B2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n222), .ZN(new_n224));
  OAI211_X1 g038(.A(KEYINPUT17), .B(G131), .C1(new_n207), .C2(new_n208), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n197), .A2(new_n198), .A3(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n203), .B1(new_n226), .B2(new_n192), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n195), .A2(new_n225), .A3(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n209), .ZN(new_n230));
  INV_X1    g044(.A(new_n214), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n224), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n223), .B1(new_n234), .B2(new_n190), .ZN(new_n235));
  OR2_X1    g049(.A1(G475), .A2(G902), .ZN(new_n236));
  OAI211_X1 g050(.A(KEYINPUT85), .B(KEYINPUT20), .C1(new_n235), .C2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT85), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n215), .A2(new_n222), .ZN(new_n239));
  INV_X1    g053(.A(new_n190), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NOR3_X1   g055(.A1(new_n209), .A2(new_n214), .A3(KEYINPUT17), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n190), .B(new_n222), .C1(new_n242), .C2(new_n228), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n236), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(KEYINPUT20), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n238), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n245), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n237), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n234), .B(new_n240), .ZN(new_n249));
  OAI21_X1  g063(.A(G475), .B1(new_n249), .B2(G902), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XOR2_X1   g065(.A(KEYINPUT9), .B(G234), .Z(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G217), .ZN(new_n254));
  NOR3_X1   g068(.A1(new_n253), .A2(new_n254), .A3(G953), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G128), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT86), .B1(new_n257), .B2(G143), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT86), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(new_n212), .A3(G128), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n212), .A2(G128), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G134), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n262), .B1(new_n258), .B2(new_n260), .ZN(new_n266));
  INV_X1    g080(.A(G134), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G122), .ZN(new_n270));
  OAI21_X1  g084(.A(KEYINPUT14), .B1(new_n270), .B2(G116), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT14), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n272), .A2(new_n273), .A3(G122), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(G116), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n271), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT87), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n276), .A2(new_n277), .A3(G107), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n273), .A2(G122), .ZN(new_n279));
  INV_X1    g093(.A(G107), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n279), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n277), .B1(new_n276), .B2(G107), .ZN(new_n282));
  INV_X1    g096(.A(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n269), .A2(new_n278), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT88), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT13), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n267), .B1(new_n263), .B2(new_n286), .ZN(new_n287));
  OR2_X1    g101(.A1(new_n264), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n279), .A2(new_n275), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G107), .ZN(new_n290));
  AOI22_X1  g104(.A1(new_n264), .A2(new_n287), .B1(new_n290), .B2(new_n281), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n288), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n284), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n285), .B1(new_n284), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n256), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(G902), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n266), .B(G134), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n278), .A2(new_n281), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(new_n282), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n288), .A2(new_n291), .ZN(new_n300));
  OAI21_X1  g114(.A(KEYINPUT88), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n284), .A2(new_n285), .A3(new_n292), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n301), .A2(new_n255), .A3(new_n302), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n295), .A2(new_n296), .A3(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G478), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(KEYINPUT15), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n306), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n295), .A2(new_n303), .A3(new_n296), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(G234), .A2(G237), .ZN(new_n311));
  INV_X1    g125(.A(G953), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(G952), .A3(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  XOR2_X1   g128(.A(KEYINPUT21), .B(G898), .Z(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n311), .A2(G902), .A3(G953), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n314), .B1(new_n316), .B2(new_n318), .ZN(new_n319));
  NOR3_X1   g133(.A1(new_n251), .A2(new_n310), .A3(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT84), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n280), .A3(G104), .ZN(new_n324));
  AND3_X1   g138(.A1(new_n189), .A2(KEYINPUT77), .A3(G107), .ZN(new_n325));
  AOI21_X1  g139(.A(KEYINPUT77), .B1(new_n189), .B2(G107), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n322), .B(new_n324), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G101), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n329), .B1(new_n280), .B2(G104), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n189), .A2(KEYINPUT77), .A3(G107), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G101), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n332), .A2(new_n333), .A3(new_n322), .A4(new_n324), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n328), .A2(KEYINPUT4), .A3(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT4), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n327), .A2(new_n336), .A3(G101), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT2), .B(G113), .ZN(new_n338));
  INV_X1    g152(.A(G119), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT65), .B1(new_n339), .B2(G116), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT65), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n341), .A2(new_n273), .A3(G119), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g157(.A1(new_n273), .A2(G119), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n340), .B2(new_n342), .ZN(new_n346));
  INV_X1    g160(.A(new_n338), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n335), .A2(new_n337), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n280), .A2(G104), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n189), .A2(G107), .ZN(new_n352));
  OAI21_X1  g166(.A(G101), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n334), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n346), .A2(KEYINPUT5), .ZN(new_n356));
  INV_X1    g170(.A(G113), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT5), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n344), .B2(new_n358), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n356), .A2(new_n359), .B1(new_n346), .B2(new_n347), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n355), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(G110), .B(G122), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n350), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  AND2_X1   g177(.A1(KEYINPUT0), .A2(G128), .ZN(new_n364));
  XNOR2_X1  g178(.A(G143), .B(G146), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT64), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n212), .A2(G146), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n203), .A2(G143), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NOR2_X1   g184(.A1(KEYINPUT0), .A2(G128), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n364), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n370), .A2(new_n372), .A3(KEYINPUT64), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G125), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n212), .A2(G146), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n203), .A2(G143), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT1), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G128), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n257), .A2(new_n376), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n381), .A2(new_n368), .A3(new_n369), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n380), .A2(new_n191), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT82), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n380), .A2(KEYINPUT82), .A3(new_n191), .A4(new_n382), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n375), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT7), .ZN(new_n388));
  INV_X1    g202(.A(G224), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n389), .A2(G953), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n387), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI22_X1  g205(.A1(G125), .A2(new_n374), .B1(new_n383), .B2(new_n384), .ZN(new_n392));
  INV_X1    g206(.A(new_n390), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n392), .A2(KEYINPUT7), .A3(new_n393), .A4(new_n386), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n363), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  XOR2_X1   g209(.A(new_n362), .B(KEYINPUT8), .Z(new_n396));
  AOI21_X1  g210(.A(new_n396), .B1(new_n360), .B2(new_n354), .ZN(new_n397));
  INV_X1    g211(.A(new_n359), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT83), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n356), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n346), .A2(KEYINPUT83), .A3(KEYINPUT5), .ZN(new_n401));
  AOI22_X1  g215(.A1(new_n400), .A2(new_n401), .B1(new_n346), .B2(new_n347), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n397), .B1(new_n402), .B2(new_n354), .ZN(new_n403));
  AOI21_X1  g217(.A(G902), .B1(new_n395), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n350), .A2(new_n361), .ZN(new_n405));
  INV_X1    g219(.A(new_n362), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT6), .A3(new_n363), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n387), .B(new_n390), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT6), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n405), .A2(new_n410), .A3(new_n406), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n404), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n404), .A2(new_n412), .A3(new_n414), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(G214), .B1(G237), .B2(G902), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n321), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n404), .A2(new_n412), .A3(new_n414), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n414), .B1(new_n404), .B2(new_n412), .ZN(new_n422));
  OAI211_X1 g236(.A(new_n321), .B(new_n419), .C1(new_n421), .C2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n320), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(new_n374), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n335), .A2(new_n426), .A3(new_n337), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT78), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT79), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n382), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n381), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(new_n432), .A3(new_n380), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n334), .A3(new_n353), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT10), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n377), .A2(new_n379), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n376), .A2(new_n257), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n382), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n439), .A2(new_n435), .ZN(new_n440));
  AOI22_X1  g254(.A1(new_n434), .A2(new_n435), .B1(new_n355), .B2(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n335), .A2(KEYINPUT78), .A3(new_n426), .A4(new_n337), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n429), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT11), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n444), .B1(new_n267), .B2(G137), .ZN(new_n445));
  INV_X1    g259(.A(G137), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT11), .A3(G134), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n267), .A2(G137), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G131), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n445), .A2(new_n447), .A3(new_n210), .A4(new_n448), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n429), .A2(new_n441), .A3(new_n454), .A4(new_n442), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G140), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n312), .A2(G227), .ZN(new_n458));
  XNOR2_X1  g272(.A(new_n457), .B(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n456), .A2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT80), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n354), .A2(new_n439), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n454), .B1(new_n434), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n462), .B1(new_n464), .B2(KEYINPUT12), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT12), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n438), .B1(new_n334), .B2(new_n353), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n355), .B2(new_n433), .ZN(new_n468));
  OAI211_X1 g282(.A(KEYINPUT80), .B(new_n466), .C1(new_n468), .C2(new_n454), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n464), .A2(KEYINPUT12), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n465), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n459), .A3(new_n455), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n461), .A2(KEYINPUT81), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(G469), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT81), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n471), .A2(new_n475), .A3(new_n459), .A4(new_n455), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n473), .A2(new_n474), .A3(new_n296), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n456), .A2(new_n459), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT76), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n471), .B2(new_n455), .ZN(new_n480));
  AOI21_X1  g294(.A(KEYINPUT76), .B1(new_n471), .B2(new_n455), .ZN(new_n481));
  OAI22_X1  g295(.A1(new_n478), .A2(new_n480), .B1(new_n481), .B2(new_n459), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(G469), .ZN(new_n483));
  NAND2_X1  g297(.A1(G469), .A2(G902), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(G221), .B1(new_n253), .B2(G902), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT75), .Z(new_n487));
  NAND2_X1  g301(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n187), .B1(new_n425), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n248), .A2(new_n250), .ZN(new_n490));
  INV_X1    g304(.A(new_n319), .ZN(new_n491));
  NAND4_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n307), .A4(new_n309), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT84), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n492), .B1(new_n494), .B2(new_n423), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n495), .A2(KEYINPUT89), .A3(new_n485), .A4(new_n487), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n452), .A2(new_n367), .A3(new_n373), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n346), .B(new_n338), .ZN(new_n498));
  INV_X1    g312(.A(new_n448), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n267), .A2(G137), .ZN(new_n500));
  OAI21_X1  g314(.A(G131), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n438), .A2(new_n451), .A3(new_n501), .ZN(new_n502));
  AND3_X1   g316(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n498), .B1(new_n497), .B2(new_n502), .ZN(new_n504));
  OAI211_X1 g318(.A(KEYINPUT66), .B(KEYINPUT28), .C1(new_n503), .C2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT28), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n502), .B1(new_n454), .B2(new_n374), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n349), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n497), .A2(new_n498), .A3(new_n502), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT66), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n511), .B1(new_n509), .B2(new_n506), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n505), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n205), .A2(G210), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT30), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n507), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n497), .A2(KEYINPUT30), .A3(new_n502), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n349), .A3(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT31), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n509), .A4(new_n517), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n509), .A3(new_n517), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(KEYINPUT31), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n519), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(G472), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT32), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n529), .ZN(new_n533));
  AOI22_X1  g347(.A1(new_n513), .A2(new_n518), .B1(KEYINPUT31), .B2(new_n526), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n533), .B1(new_n534), .B2(new_n525), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT32), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n523), .A2(new_n509), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n518), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT29), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n538), .B(new_n539), .C1(new_n513), .C2(new_n518), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n508), .A2(KEYINPUT67), .A3(new_n509), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT67), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n504), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(KEYINPUT28), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n509), .A2(new_n506), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n544), .A2(KEYINPUT29), .A3(new_n517), .A4(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n296), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G472), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n532), .A2(new_n536), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT73), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n254), .B1(G234), .B2(new_n296), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n257), .A2(G119), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT23), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n257), .A2(G119), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n553), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(G110), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n257), .A2(KEYINPUT23), .A3(G119), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT69), .ZN(new_n559));
  AND2_X1   g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n558), .A2(new_n559), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n556), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT68), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n339), .B2(G128), .ZN(new_n564));
  NOR3_X1   g378(.A1(new_n257), .A2(KEYINPUT68), .A3(G119), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n555), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g380(.A(KEYINPUT24), .B(G110), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n562), .A2(KEYINPUT70), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g383(.A(KEYINPUT70), .B1(new_n562), .B2(new_n568), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n195), .A2(new_n220), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n195), .A2(new_n227), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G110), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n566), .A2(new_n567), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n312), .A2(G221), .A3(G234), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n579), .B(KEYINPUT71), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT22), .B(G137), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n580), .B(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n572), .A2(new_n578), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n562), .A2(new_n568), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT70), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n562), .A2(KEYINPUT70), .A3(new_n568), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n587), .A2(new_n220), .A3(new_n195), .A4(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n582), .B1(new_n589), .B2(new_n577), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n296), .B1(new_n584), .B2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT25), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n583), .B1(new_n572), .B2(new_n578), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n589), .A2(new_n577), .A3(new_n582), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(KEYINPUT25), .A3(new_n296), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n552), .B1(new_n593), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n551), .A2(G902), .ZN(new_n599));
  XOR2_X1   g413(.A(new_n599), .B(KEYINPUT72), .Z(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n550), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(KEYINPUT25), .B1(new_n596), .B2(new_n296), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n592), .B(G902), .C1(new_n594), .C2(new_n595), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n551), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT73), .A3(new_n602), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n549), .A2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT74), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n531), .B(new_n533), .C1(new_n534), .C2(new_n525), .ZN(new_n613));
  AOI21_X1  g427(.A(KEYINPUT32), .B1(new_n528), .B2(new_n529), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI22_X1  g429(.A1(new_n615), .A2(new_n548), .B1(new_n604), .B2(new_n608), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT74), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n489), .A2(new_n496), .A3(new_n612), .A4(new_n617), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n618), .B(G101), .ZN(G3));
  NAND2_X1  g433(.A1(new_n528), .A2(new_n296), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n535), .B1(new_n620), .B2(G472), .ZN(new_n621));
  AND4_X1   g435(.A1(new_n485), .A2(new_n609), .A3(new_n487), .A4(new_n621), .ZN(new_n622));
  OAI211_X1 g436(.A(new_n491), .B(new_n419), .C1(new_n421), .C2(new_n422), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n305), .A2(G902), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n293), .A2(new_n294), .A3(new_n256), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n255), .B1(new_n301), .B2(new_n302), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n626), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n295), .A2(KEYINPUT33), .A3(new_n303), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n625), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT90), .B(G478), .Z(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n304), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n251), .B1(new_n631), .B2(new_n634), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n623), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n622), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(KEYINPUT91), .ZN(new_n638));
  XNOR2_X1  g452(.A(KEYINPUT34), .B(G104), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  INV_X1    g454(.A(new_n622), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n310), .A2(new_n250), .A3(new_n248), .ZN(new_n642));
  NOR3_X1   g456(.A1(new_n641), .A2(new_n623), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT35), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  NAND2_X1  g459(.A1(new_n620), .A2(G472), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n530), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT36), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n590), .A2(new_n648), .ZN(new_n649));
  OAI211_X1 g463(.A(new_n589), .B(new_n577), .C1(KEYINPUT36), .C2(new_n582), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n651));
  AND3_X1   g465(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n651), .B1(new_n649), .B2(new_n650), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n652), .A2(new_n653), .A3(new_n600), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n598), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n489), .A2(new_n496), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT37), .B(G110), .Z(new_n658));
  XNOR2_X1  g472(.A(new_n657), .B(new_n658), .ZN(G12));
  NOR2_X1   g473(.A1(new_n655), .A2(new_n493), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n660), .A2(new_n549), .A3(new_n485), .A4(new_n487), .ZN(new_n661));
  OR2_X1    g475(.A1(new_n317), .A2(G900), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n314), .B1(new_n662), .B2(KEYINPUT94), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n663), .B1(KEYINPUT94), .B2(new_n662), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n490), .A2(new_n310), .A3(new_n664), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(new_n257), .ZN(G30));
  XOR2_X1   g481(.A(new_n664), .B(KEYINPUT39), .Z(new_n668));
  NOR2_X1   g482(.A1(new_n488), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AND2_X1   g484(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n670), .A2(KEYINPUT40), .ZN(new_n672));
  XOR2_X1   g486(.A(new_n418), .B(KEYINPUT38), .Z(new_n673));
  NAND2_X1  g487(.A1(new_n537), .A2(new_n517), .ZN(new_n674));
  AND2_X1   g488(.A1(new_n541), .A2(new_n543), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n674), .B(new_n296), .C1(new_n675), .C2(new_n517), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n532), .A2(new_n536), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n251), .A2(new_n310), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n655), .A2(new_n419), .ZN(new_n681));
  OR4_X1    g495(.A1(new_n673), .A2(new_n679), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n671), .A2(new_n672), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(new_n212), .ZN(G45));
  OAI211_X1 g498(.A(new_n251), .B(new_n664), .C1(new_n631), .C2(new_n634), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n661), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT95), .B(G146), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G48));
  INV_X1    g502(.A(KEYINPUT96), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n636), .A2(new_n549), .A3(new_n609), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n472), .A2(KEYINPUT81), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n459), .B1(new_n453), .B2(new_n455), .ZN(new_n692));
  OAI211_X1 g506(.A(new_n296), .B(new_n476), .C1(new_n691), .C2(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(G469), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n694), .A2(new_n477), .A3(new_n486), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n689), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n694), .A2(new_n477), .A3(new_n486), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n616), .A2(KEYINPUT96), .A3(new_n636), .A4(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  INV_X1    g515(.A(new_n419), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n702), .B1(new_n416), .B2(new_n417), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n310), .A2(new_n491), .A3(new_n250), .A4(new_n248), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n604), .B2(new_n608), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n697), .A2(new_n703), .A3(new_n549), .A4(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT97), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n694), .A2(new_n703), .A3(new_n477), .A4(new_n486), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n709), .A2(new_n710), .A3(new_n549), .A4(new_n705), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n707), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G116), .ZN(G18));
  INV_X1    g527(.A(new_n549), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n654), .A2(new_n598), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n320), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n714), .A2(new_n708), .A3(new_n716), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n339), .ZN(G21));
  NAND2_X1  g532(.A1(new_n544), .A2(new_n545), .ZN(new_n719));
  AOI22_X1  g533(.A1(new_n719), .A2(new_n518), .B1(KEYINPUT31), .B2(new_n526), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n525), .B1(new_n720), .B2(KEYINPUT98), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n518), .ZN(new_n722));
  AND3_X1   g536(.A1(new_n722), .A2(KEYINPUT98), .A3(new_n527), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n529), .B1(new_n721), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n598), .A2(new_n603), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n724), .A2(new_n725), .A3(new_n646), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(KEYINPUT99), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT99), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n728), .A3(new_n725), .A4(new_n646), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n708), .A2(new_n319), .A3(new_n680), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  INV_X1    g547(.A(new_n685), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n734), .A2(new_n724), .A3(new_n715), .A4(new_n646), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n708), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n191), .ZN(G27));
  XOR2_X1   g551(.A(new_n484), .B(KEYINPUT100), .Z(new_n738));
  NAND3_X1  g552(.A1(new_n477), .A2(new_n483), .A3(new_n738), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n418), .A2(new_n702), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n739), .A2(new_n486), .A3(new_n740), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n549), .A2(new_n725), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n742), .A3(new_n734), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n739), .A2(new_n486), .A3(new_n740), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n744), .A2(new_n610), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n685), .A2(KEYINPUT42), .ZN(new_n746));
  AOI22_X1  g560(.A1(new_n743), .A2(KEYINPUT42), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G131), .ZN(G33));
  XNOR2_X1  g562(.A(new_n665), .B(KEYINPUT101), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n741), .A2(new_n749), .A3(new_n616), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT102), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n745), .A2(KEYINPUT102), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  NAND2_X1  g569(.A1(new_n647), .A2(new_n715), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT106), .Z(new_n757));
  NOR2_X1   g571(.A1(new_n631), .A2(new_n634), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n251), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(KEYINPUT105), .A3(KEYINPUT43), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n767));
  XOR2_X1   g581(.A(new_n767), .B(KEYINPUT107), .Z(new_n768));
  OR2_X1    g582(.A1(new_n482), .A2(KEYINPUT45), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n482), .A2(KEYINPUT45), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(G469), .A3(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT46), .B1(new_n771), .B2(new_n738), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n772), .A2(KEYINPUT104), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(KEYINPUT46), .A3(new_n738), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(KEYINPUT103), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n772), .A2(KEYINPUT104), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n773), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g591(.A(new_n477), .B1(new_n774), .B2(KEYINPUT103), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n668), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n486), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OR2_X1    g596(.A1(new_n766), .A2(KEYINPUT44), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n768), .A2(new_n740), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G137), .ZN(G39));
  INV_X1    g599(.A(KEYINPUT47), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n779), .A2(new_n786), .A3(new_n486), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n486), .B1(new_n777), .B2(new_n778), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(KEYINPUT47), .ZN(new_n789));
  INV_X1    g603(.A(new_n740), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n790), .A2(new_n549), .A3(new_n609), .A4(new_n685), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n787), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NOR2_X1   g607(.A1(G952), .A2(G953), .ZN(new_n794));
  AND2_X1   g608(.A1(new_n712), .A2(new_n657), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n717), .B1(new_n696), .B2(new_n698), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n319), .B1(new_n635), .B2(new_n642), .ZN(new_n797));
  OAI21_X1  g611(.A(new_n797), .B1(new_n420), .B2(new_n424), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  AOI22_X1  g613(.A1(new_n730), .A2(new_n731), .B1(new_n622), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n795), .A2(new_n618), .A3(new_n796), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n735), .A2(new_n744), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n488), .A2(new_n714), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n251), .A2(new_n310), .ZN(new_n804));
  AND4_X1   g618(.A1(new_n804), .A2(new_n740), .A3(new_n715), .A4(new_n664), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n802), .B1(new_n803), .B2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n754), .A2(new_n747), .A3(new_n806), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT108), .B1(new_n801), .B2(new_n807), .ZN(new_n808));
  OAI22_X1  g622(.A1(new_n661), .A2(new_n665), .B1(new_n735), .B2(new_n708), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n686), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n655), .A2(new_n664), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n811), .A2(new_n678), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n739), .A2(new_n486), .ZN(new_n813));
  INV_X1    g627(.A(new_n813), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n493), .A2(new_n680), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n812), .A2(new_n814), .A3(KEYINPUT109), .A4(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(KEYINPUT109), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n811), .A2(new_n678), .A3(new_n815), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n817), .B1(new_n818), .B2(new_n813), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n810), .A2(new_n820), .A3(KEYINPUT52), .ZN(new_n821));
  AOI21_X1  g635(.A(KEYINPUT52), .B1(new_n810), .B2(new_n820), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n807), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n796), .A2(new_n800), .A3(new_n618), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n712), .A2(new_n657), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT108), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n825), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n808), .A2(new_n824), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(KEYINPUT53), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n810), .A2(new_n820), .A3(KEYINPUT52), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n823), .B2(new_n834), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT53), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n808), .A3(new_n837), .A4(new_n830), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n832), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  NOR3_X1   g654(.A1(new_n801), .A2(new_n837), .A3(new_n807), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n836), .A2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n829), .B1(new_n825), .B2(new_n828), .ZN(new_n843));
  NOR4_X1   g657(.A1(new_n807), .A2(new_n826), .A3(KEYINPUT108), .A4(new_n827), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n843), .A2(new_n844), .A3(new_n823), .ZN(new_n845));
  OAI211_X1 g659(.A(new_n840), .B(new_n842), .C1(new_n845), .C2(KEYINPUT53), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n839), .A2(new_n846), .A3(KEYINPUT111), .ZN(new_n847));
  AOI21_X1  g661(.A(KEYINPUT111), .B1(new_n839), .B2(new_n846), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI211_X1 g663(.A(new_n313), .B(new_n765), .C1(new_n729), .C2(new_n727), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n850), .A2(new_n740), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n787), .A2(new_n789), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n694), .A2(new_n477), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(new_n487), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n851), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n697), .A2(new_n314), .A3(new_n740), .ZN(new_n856));
  AOI211_X1 g670(.A(new_n678), .B(new_n856), .C1(new_n604), .C2(new_n608), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(new_n490), .A3(new_n758), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n765), .A2(new_n856), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n646), .A3(new_n715), .A4(new_n724), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT50), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n673), .A2(new_n697), .A3(new_n702), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n850), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT114), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n863), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI211_X1 g681(.A(KEYINPUT114), .B(KEYINPUT50), .C1(new_n850), .C2(new_n864), .ZN(new_n868));
  OAI211_X1 g682(.A(KEYINPUT51), .B(new_n862), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  OR2_X1    g683(.A1(new_n855), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n859), .A2(new_n871), .A3(new_n742), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n871), .B1(new_n859), .B2(new_n742), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n850), .A2(new_n709), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n312), .A2(G952), .ZN(new_n877));
  INV_X1    g691(.A(new_n635), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n857), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n873), .A2(new_n874), .ZN(new_n881));
  OR3_X1    g695(.A1(new_n880), .A2(KEYINPUT116), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g696(.A(KEYINPUT116), .B1(new_n880), .B2(new_n881), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n870), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT51), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n854), .B(KEYINPUT112), .ZN(new_n887));
  INV_X1    g701(.A(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n888), .B1(new_n787), .B2(new_n789), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT113), .ZN(new_n890));
  OR3_X1    g704(.A1(new_n889), .A2(new_n890), .A3(new_n851), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n867), .A2(new_n868), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n889), .B2(new_n851), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n891), .A2(new_n892), .A3(new_n862), .A4(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n885), .B1(new_n886), .B2(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n794), .B1(new_n849), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n725), .A2(new_n487), .A3(new_n419), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n760), .A2(new_n678), .A3(new_n897), .ZN(new_n898));
  OR2_X1    g712(.A1(new_n853), .A2(KEYINPUT49), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n853), .A2(KEYINPUT49), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n898), .A2(new_n673), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(KEYINPUT117), .B1(new_n896), .B2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n839), .A2(new_n846), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT111), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n894), .A2(new_n886), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n839), .A2(new_n846), .A3(KEYINPUT111), .ZN(new_n909));
  INV_X1    g723(.A(new_n885), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n907), .A2(new_n908), .A3(new_n909), .A4(new_n910), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n904), .B(new_n901), .C1(new_n911), .C2(new_n794), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n903), .A2(new_n912), .ZN(G75));
  NOR2_X1   g727(.A1(new_n312), .A2(G952), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT120), .Z(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AOI22_X1  g730(.A1(new_n831), .A2(new_n837), .B1(new_n836), .B2(new_n841), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n296), .ZN(new_n918));
  AOI21_X1  g732(.A(KEYINPUT56), .B1(new_n918), .B2(G210), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n408), .A2(new_n411), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(new_n409), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n921), .B(new_n922), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n916), .B1(new_n919), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n831), .A2(new_n837), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n842), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n928), .A2(KEYINPUT119), .A3(G902), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT119), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n930), .B1(new_n917), .B2(new_n296), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n926), .B1(new_n932), .B2(new_n415), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n924), .A2(new_n933), .ZN(G51));
  AOI21_X1  g748(.A(new_n771), .B1(new_n929), .B2(new_n931), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n473), .A2(new_n476), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n738), .B(KEYINPUT121), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n938), .B(KEYINPUT57), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n927), .A2(new_n840), .A3(new_n842), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n840), .B1(new_n927), .B2(new_n842), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n935), .B1(new_n937), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(KEYINPUT122), .B1(new_n943), .B2(new_n914), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT122), .ZN(new_n945));
  INV_X1    g759(.A(new_n914), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n942), .A2(new_n937), .ZN(new_n947));
  OAI211_X1 g761(.A(new_n945), .B(new_n946), .C1(new_n947), .C2(new_n935), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n944), .A2(new_n948), .ZN(G54));
  AND3_X1   g763(.A1(new_n932), .A2(KEYINPUT58), .A3(G475), .ZN(new_n950));
  INV_X1    g764(.A(new_n235), .ZN(new_n951));
  AND2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n952), .A2(new_n953), .ZN(G60));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n629), .A2(new_n630), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n907), .A2(new_n909), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT59), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n956), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n956), .A2(new_n959), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n940), .B2(new_n941), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(KEYINPUT123), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT123), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n964), .B(new_n961), .C1(new_n940), .C2(new_n941), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n963), .A2(new_n916), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n955), .B1(new_n960), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n959), .B1(new_n847), .B2(new_n848), .ZN(new_n968));
  INV_X1    g782(.A(new_n956), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n915), .B1(new_n962), .B2(KEYINPUT123), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n970), .A2(KEYINPUT124), .A3(new_n965), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n967), .A2(new_n972), .ZN(G63));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n917), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n652), .A2(new_n653), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n915), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n596), .B2(new_n976), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g794(.A(G953), .B1(new_n316), .B2(new_n389), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n981), .B1(new_n828), .B2(G953), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n920), .B1(G898), .B2(new_n312), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n982), .B(new_n983), .ZN(G69));
  AND2_X1   g798(.A1(new_n784), .A2(new_n792), .ZN(new_n985));
  INV_X1    g799(.A(new_n810), .ZN(new_n986));
  NOR2_X1   g800(.A1(new_n683), .A2(new_n986), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT62), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n635), .A2(new_n642), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n989), .A2(KEYINPUT125), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n989), .A2(KEYINPUT125), .ZN(new_n991));
  NOR3_X1   g805(.A1(new_n990), .A2(new_n991), .A3(new_n790), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n992), .A2(new_n612), .A3(new_n617), .A4(new_n669), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n985), .A2(new_n988), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n312), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n521), .A2(new_n522), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n200), .A2(new_n202), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n996), .B(new_n997), .Z(new_n998));
  NAND2_X1  g812(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(G900), .B2(G953), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n754), .A2(new_n747), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT127), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n742), .A2(new_n815), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n986), .B1(new_n782), .B2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n985), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1000), .B1(new_n1005), .B2(G953), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n999), .A2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n312), .B1(G227), .B2(G900), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1008), .B1(new_n1006), .B2(KEYINPUT126), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI211_X1 g824(.A(new_n999), .B(new_n1006), .C1(KEYINPUT126), .C2(new_n1008), .ZN(new_n1011));
  AND2_X1   g825(.A1(new_n1010), .A2(new_n1011), .ZN(G72));
  NAND2_X1  g826(.A1(G472), .A2(G902), .ZN(new_n1013));
  XOR2_X1   g827(.A(new_n1013), .B(KEYINPUT63), .Z(new_n1014));
  OAI21_X1  g828(.A(new_n1014), .B1(new_n994), .B2(new_n801), .ZN(new_n1015));
  INV_X1    g829(.A(new_n674), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n914), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1014), .B1(new_n1005), .B2(new_n801), .ZN(new_n1018));
  NAND4_X1  g832(.A1(new_n1018), .A2(new_n509), .A3(new_n523), .A4(new_n518), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n538), .A2(new_n526), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n832), .A2(new_n838), .A3(new_n1014), .A4(new_n1020), .ZN(new_n1021));
  AND3_X1   g835(.A1(new_n1017), .A2(new_n1019), .A3(new_n1021), .ZN(G57));
endmodule


