//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n702, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n931, new_n932, new_n933, new_n934, new_n935, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  NOR2_X1   g002(.A1(new_n187), .A2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G104), .ZN(new_n192));
  INV_X1    g006(.A(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT78), .B1(new_n195), .B2(G101), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT78), .ZN(new_n197));
  INV_X1    g011(.A(G101), .ZN(new_n198));
  AOI211_X1 g012(.A(new_n197), .B(new_n198), .C1(new_n192), .C2(new_n194), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n193), .B2(G107), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT77), .B1(new_n191), .B2(G104), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT3), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n202), .A2(new_n191), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT77), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(new_n193), .A3(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n205), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n196), .A2(new_n199), .B1(G101), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n209), .A2(new_n211), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  XNOR2_X1  g030(.A(G143), .B(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n211), .A2(KEYINPUT1), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G128), .ZN(new_n220));
  INV_X1    g034(.A(new_n217), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n216), .A2(new_n218), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NOR3_X1   g036(.A1(new_n207), .A2(new_n222), .A3(KEYINPUT79), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n224));
  AND4_X1   g038(.A1(new_n200), .A2(new_n201), .A3(new_n203), .A4(new_n205), .ZN(new_n225));
  XNOR2_X1  g039(.A(G104), .B(G107), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n197), .B1(new_n226), .B2(new_n198), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n195), .A2(KEYINPUT78), .A3(G101), .ZN(new_n228));
  AOI22_X1  g042(.A1(new_n198), .A2(new_n225), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT68), .B1(new_n217), .B2(new_n209), .ZN(new_n230));
  AND4_X1   g044(.A1(KEYINPUT68), .A2(new_n209), .A3(new_n211), .A4(new_n213), .ZN(new_n231));
  AOI21_X1  g045(.A(new_n208), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n232));
  OAI22_X1  g046(.A1(new_n230), .A2(new_n231), .B1(new_n217), .B2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n224), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT64), .B1(new_n210), .B2(G143), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT64), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(new_n212), .A3(G146), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n235), .A2(new_n237), .B1(G143), .B2(new_n210), .ZN(new_n238));
  OAI22_X1  g052(.A1(new_n230), .A2(new_n231), .B1(new_n238), .B2(new_n232), .ZN(new_n239));
  OAI22_X1  g053(.A1(new_n223), .A2(new_n234), .B1(new_n239), .B2(new_n229), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT11), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G137), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(G137), .ZN(new_n244));
  INV_X1    g058(.A(G137), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT11), .A3(G134), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(G131), .ZN(new_n248));
  INV_X1    g062(.A(G131), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n243), .A2(new_n246), .A3(new_n249), .A4(new_n244), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT12), .B1(new_n251), .B2(KEYINPUT80), .ZN(new_n252));
  INV_X1    g066(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n240), .A2(new_n251), .A3(new_n253), .ZN(new_n254));
  OAI21_X1  g068(.A(KEYINPUT79), .B1(new_n207), .B2(new_n222), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n201), .A2(new_n205), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n256), .A2(new_n198), .A3(new_n200), .A4(new_n203), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n227), .A2(new_n228), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n233), .A2(new_n224), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n239), .ZN(new_n260));
  AOI22_X1  g074(.A1(new_n255), .A2(new_n259), .B1(new_n260), .B2(new_n207), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n248), .A2(new_n250), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n252), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n254), .A2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT10), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n265), .B1(new_n223), .B2(new_n234), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n206), .A2(G101), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n257), .A2(KEYINPUT4), .A3(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n236), .B1(new_n212), .B2(G146), .ZN(new_n269));
  NOR3_X1   g083(.A1(new_n210), .A2(KEYINPUT64), .A3(G143), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n211), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  AND2_X1   g085(.A1(KEYINPUT0), .A2(G128), .ZN(new_n272));
  NOR2_X1   g086(.A1(KEYINPUT0), .A2(G128), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n271), .A2(new_n274), .B1(new_n217), .B2(new_n272), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n206), .A2(new_n276), .A3(G101), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n229), .A2(KEYINPUT10), .A3(new_n239), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n266), .A2(new_n280), .A3(new_n262), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n264), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(G110), .B(G140), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT76), .ZN(new_n284));
  INV_X1    g098(.A(G953), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G227), .ZN(new_n286));
  XNOR2_X1  g100(.A(new_n284), .B(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(KEYINPUT10), .B1(new_n255), .B2(new_n259), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n278), .A2(new_n279), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n251), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  NOR3_X1   g104(.A1(new_n288), .A2(new_n289), .A3(new_n251), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n287), .ZN(new_n292));
  AOI22_X1  g106(.A1(new_n282), .A2(new_n287), .B1(new_n290), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G469), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n281), .A2(new_n290), .ZN(new_n295));
  AOI22_X1  g109(.A1(new_n292), .A2(new_n264), .B1(new_n295), .B2(new_n287), .ZN(new_n296));
  NOR4_X1   g110(.A1(new_n296), .A2(KEYINPUT81), .A3(G469), .A4(G902), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n298));
  INV_X1    g112(.A(new_n287), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n253), .B1(new_n240), .B2(new_n251), .ZN(new_n300));
  NOR3_X1   g114(.A1(new_n261), .A2(new_n262), .A3(new_n252), .ZN(new_n301));
  OAI211_X1 g115(.A(new_n281), .B(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n262), .B1(new_n266), .B2(new_n280), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n287), .B1(new_n303), .B2(new_n291), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n298), .B1(new_n305), .B2(new_n187), .ZN(new_n306));
  OAI211_X1 g120(.A(new_n190), .B(new_n294), .C1(new_n297), .C2(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT9), .B(G234), .ZN(new_n308));
  XNOR2_X1  g122(.A(new_n308), .B(KEYINPUT75), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n188), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G221), .ZN(new_n311));
  OAI21_X1  g125(.A(G214), .B1(G237), .B2(G902), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G116), .ZN(new_n315));
  INV_X1    g129(.A(G116), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G119), .ZN(new_n317));
  AND2_X1   g131(.A1(new_n315), .A2(new_n317), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT2), .B(G113), .Z(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n315), .A2(new_n317), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n268), .A2(new_n324), .A3(new_n277), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n318), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G113), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT82), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT82), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT5), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n315), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n327), .A2(new_n335), .B1(new_n318), .B2(new_n319), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n229), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n325), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(G110), .B(G122), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n325), .A2(new_n337), .A3(new_n339), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n341), .A2(KEYINPUT6), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n338), .A2(new_n344), .A3(new_n340), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n216), .A2(new_n218), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n271), .A2(new_n220), .ZN(new_n347));
  INV_X1    g161(.A(G125), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n217), .A2(new_n272), .ZN(new_n350));
  INV_X1    g164(.A(new_n274), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n350), .B1(new_n238), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(G125), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G224), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n355), .A2(G953), .ZN(new_n356));
  XNOR2_X1  g170(.A(new_n354), .B(new_n356), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n343), .A2(new_n345), .A3(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT83), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n343), .A2(KEYINPUT83), .A3(new_n345), .A4(new_n357), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT7), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n349), .A2(new_n353), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n364), .B1(new_n349), .B2(new_n353), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n207), .A2(new_n336), .ZN(new_n368));
  OAI21_X1  g182(.A(G113), .B1(new_n326), .B2(new_n315), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n321), .A2(new_n329), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n320), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n257), .A3(new_n258), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n339), .B(KEYINPUT8), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n368), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT84), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n368), .A2(new_n372), .A3(KEYINPUT84), .A4(new_n373), .ZN(new_n377));
  NAND4_X1  g191(.A1(new_n367), .A2(new_n376), .A3(new_n342), .A4(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n188), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT85), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(KEYINPUT85), .A3(new_n188), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n362), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(G210), .B1(G237), .B2(G902), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n362), .A2(new_n383), .A3(new_n385), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n313), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  AND3_X1   g203(.A1(new_n307), .A2(new_n311), .A3(new_n389), .ZN(new_n390));
  XOR2_X1   g204(.A(KEYINPUT24), .B(G110), .Z(new_n391));
  XNOR2_X1  g205(.A(G119), .B(G128), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  XOR2_X1   g207(.A(new_n393), .B(KEYINPUT71), .Z(new_n394));
  NOR3_X1   g208(.A1(new_n348), .A2(KEYINPUT16), .A3(G140), .ZN(new_n395));
  XNOR2_X1  g209(.A(G125), .B(G140), .ZN(new_n396));
  AOI211_X1 g210(.A(new_n210), .B(new_n395), .C1(KEYINPUT16), .C2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(G140), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n348), .A2(new_n398), .ZN(new_n399));
  NOR2_X1   g213(.A1(G125), .A2(G140), .ZN(new_n400));
  OAI21_X1  g214(.A(KEYINPUT16), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n395), .ZN(new_n402));
  AOI21_X1  g216(.A(G146), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT23), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(G119), .B2(new_n208), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n314), .A2(KEYINPUT23), .A3(G128), .ZN(new_n408));
  OAI22_X1  g222(.A1(new_n407), .A2(new_n408), .B1(G119), .B2(new_n208), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G110), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n394), .A2(new_n405), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n401), .A2(G146), .A3(new_n402), .ZN(new_n412));
  OR2_X1    g226(.A1(new_n412), .A2(KEYINPUT72), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(KEYINPUT72), .ZN(new_n414));
  OAI22_X1  g228(.A1(new_n409), .A2(G110), .B1(new_n392), .B2(new_n391), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n396), .A2(new_n210), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n413), .A2(new_n414), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n411), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n285), .A2(G221), .A3(G234), .ZN(new_n419));
  XNOR2_X1  g233(.A(new_n419), .B(KEYINPUT22), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(G137), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  OR2_X1    g236(.A1(new_n422), .A2(KEYINPUT73), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(KEYINPUT73), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n418), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n411), .A2(KEYINPUT73), .A3(new_n422), .A4(new_n417), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n188), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT25), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n425), .B2(new_n426), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT74), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n430), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G217), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(G234), .B2(new_n188), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n429), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n435), .A2(G902), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n427), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(G101), .ZN(new_n441));
  NOR2_X1   g255(.A1(G237), .A2(G953), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(G210), .ZN(new_n443));
  XNOR2_X1  g257(.A(new_n441), .B(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n444), .B(KEYINPUT70), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n245), .A2(G134), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n249), .B1(new_n244), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT66), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT66), .ZN(new_n449));
  XNOR2_X1  g263(.A(G134), .B(G137), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n449), .B1(new_n450), .B2(new_n249), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n243), .A2(new_n244), .A3(new_n246), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n448), .A2(new_n451), .B1(new_n452), .B2(new_n249), .ZN(new_n453));
  AOI22_X1  g267(.A1(new_n453), .A2(new_n239), .B1(new_n275), .B2(new_n251), .ZN(new_n454));
  INV_X1    g268(.A(new_n324), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n456), .A2(KEYINPUT28), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n454), .B2(new_n455), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(KEYINPUT65), .B1(new_n262), .B2(new_n352), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT65), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n275), .A2(new_n462), .A3(new_n251), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n447), .A2(KEYINPUT66), .ZN(new_n465));
  AOI211_X1 g279(.A(new_n449), .B(new_n249), .C1(new_n244), .C2(new_n446), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n250), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(KEYINPUT67), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT67), .ZN(new_n469));
  OAI211_X1 g283(.A(new_n469), .B(new_n250), .C1(new_n465), .C2(new_n466), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n239), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n455), .B1(new_n464), .B2(new_n471), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n445), .B1(new_n460), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n464), .A2(new_n471), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT30), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n453), .A2(new_n239), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n275), .A2(new_n251), .ZN(new_n478));
  AND3_X1   g292(.A1(new_n477), .A2(KEYINPUT30), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n476), .A2(new_n324), .A3(new_n480), .ZN(new_n481));
  XOR2_X1   g295(.A(KEYINPUT69), .B(KEYINPUT31), .Z(new_n482));
  NAND4_X1  g296(.A1(new_n481), .A2(new_n456), .A3(new_n444), .A4(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n456), .ZN(new_n484));
  INV_X1    g298(.A(new_n444), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n479), .B1(new_n474), .B2(new_n475), .ZN(new_n486));
  AOI211_X1 g300(.A(new_n484), .B(new_n485), .C1(new_n486), .C2(new_n324), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT31), .ZN(new_n488));
  OAI211_X1 g302(.A(new_n473), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(G472), .A2(G902), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(KEYINPUT32), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT32), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n460), .A2(new_n472), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(new_n445), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n484), .B1(new_n486), .B2(new_n324), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n498), .A2(new_n444), .ZN(new_n499));
  NOR3_X1   g313(.A1(new_n497), .A2(new_n499), .A3(KEYINPUT29), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n454), .A2(new_n455), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n457), .B2(new_n459), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT29), .ZN(new_n503));
  NOR3_X1   g317(.A1(new_n502), .A2(new_n503), .A3(new_n485), .ZN(new_n504));
  OR2_X1    g318(.A1(new_n504), .A2(G902), .ZN(new_n505));
  OAI21_X1  g319(.A(G472), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n439), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(G113), .B(G122), .ZN(new_n508));
  XNOR2_X1  g322(.A(new_n508), .B(new_n193), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT86), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G143), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n212), .A2(KEYINPUT86), .ZN(new_n512));
  NAND4_X1  g326(.A1(new_n511), .A2(new_n512), .A3(G214), .A4(new_n442), .ZN(new_n513));
  INV_X1    g327(.A(G237), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n514), .A2(new_n285), .A3(G214), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n212), .A2(KEYINPUT86), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n249), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(G131), .A3(new_n517), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n396), .B(KEYINPUT19), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n210), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n413), .A2(new_n521), .A3(new_n523), .A4(new_n414), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n518), .B1(KEYINPUT18), .B2(G131), .ZN(new_n525));
  NAND2_X1  g339(.A1(KEYINPUT18), .A2(G131), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n526), .B1(new_n513), .B2(new_n517), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n396), .A2(new_n210), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT87), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n416), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n396), .A2(KEYINPUT87), .A3(new_n210), .ZN(new_n531));
  OAI22_X1  g345(.A1(new_n525), .A2(new_n527), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n509), .B1(new_n524), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n519), .A2(new_n534), .A3(new_n520), .ZN(new_n535));
  OR2_X1    g349(.A1(new_n520), .A2(new_n534), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n404), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n509), .A3(new_n532), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT88), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT88), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n537), .A2(new_n532), .A3(new_n540), .A4(new_n509), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n533), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n542), .A2(G475), .A3(G902), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n539), .A2(new_n541), .ZN(new_n544));
  INV_X1    g358(.A(new_n533), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT89), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT20), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(G475), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n546), .A2(new_n550), .A3(new_n188), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT89), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n548), .B1(new_n542), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n537), .A2(new_n532), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n544), .B1(new_n509), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n188), .ZN(new_n557));
  AOI22_X1  g371(.A1(new_n549), .A2(new_n554), .B1(G475), .B2(new_n557), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n285), .A2(G952), .ZN(new_n559));
  NAND2_X1  g373(.A1(G234), .A2(G237), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g375(.A(KEYINPUT21), .B(G898), .Z(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(G902), .A3(G953), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n309), .A2(G217), .A3(new_n285), .ZN(new_n565));
  XNOR2_X1  g379(.A(G128), .B(G143), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT13), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n212), .A2(G128), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n567), .B(G134), .C1(KEYINPUT13), .C2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(G122), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(G116), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n316), .A2(G122), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(G107), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n572), .A3(new_n191), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n574), .A2(new_n575), .B1(new_n242), .B2(new_n566), .ZN(new_n576));
  INV_X1    g390(.A(new_n575), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n570), .A2(G116), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT14), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n571), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT90), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n578), .A2(new_n579), .ZN(new_n583));
  OAI211_X1 g397(.A(KEYINPUT90), .B(new_n571), .C1(new_n578), .C2(new_n579), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n577), .B1(new_n585), .B2(G107), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n566), .B(new_n242), .ZN(new_n587));
  AOI221_X4 g401(.A(new_n565), .B1(new_n569), .B2(new_n576), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(new_n565), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n587), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n576), .A2(new_n569), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n589), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OR2_X1    g406(.A1(new_n588), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n188), .ZN(new_n594));
  INV_X1    g408(.A(G478), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n595), .A2(KEYINPUT15), .ZN(new_n596));
  XOR2_X1   g410(.A(new_n594), .B(new_n596), .Z(new_n597));
  AND3_X1   g411(.A1(new_n558), .A2(new_n564), .A3(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n390), .A2(new_n507), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n489), .A2(new_n188), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT91), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT91), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n489), .A2(new_n603), .A3(new_n188), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(G472), .A3(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT92), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n602), .A2(KEYINPUT92), .A3(G472), .A4(new_n604), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(new_n491), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n311), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n300), .A2(new_n301), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n281), .A2(new_n299), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n304), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n187), .A3(new_n188), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(KEYINPUT81), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n305), .A2(new_n298), .A3(new_n187), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n615), .A2(new_n616), .B1(G469), .B2(new_n293), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n610), .B1(new_n617), .B2(new_n190), .ZN(new_n618));
  INV_X1    g432(.A(new_n439), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n609), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT93), .ZN(new_n622));
  AOI21_X1  g436(.A(G478), .B1(new_n593), .B2(new_n188), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT94), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n624), .B1(new_n588), .B2(new_n592), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(new_n624), .B(KEYINPUT33), .C1(new_n588), .C2(new_n592), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n623), .B1(new_n629), .B2(G478), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n549), .A2(new_n554), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n557), .A2(G475), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  AND3_X1   g448(.A1(new_n362), .A2(new_n383), .A3(new_n385), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n385), .B1(new_n362), .B2(new_n383), .ZN(new_n636));
  OAI211_X1 g450(.A(new_n312), .B(new_n564), .C1(new_n635), .C2(new_n636), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n634), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n622), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n597), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n543), .B(new_n548), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n642), .A2(new_n632), .A3(new_n643), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n637), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n622), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT35), .B(G107), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G9));
  AND2_X1   g462(.A1(new_n607), .A2(new_n608), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n598), .A2(new_n307), .A3(new_n311), .A4(new_n389), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n422), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n418), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n437), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n436), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n650), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n649), .A2(new_n655), .A3(new_n491), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT37), .Z(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G110), .ZN(G12));
  AOI21_X1  g472(.A(new_n654), .B1(new_n495), .B2(new_n506), .ZN(new_n659));
  OR2_X1    g473(.A1(new_n563), .A2(G900), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n561), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n644), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n390), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT95), .B(G128), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G30));
  XNOR2_X1  g480(.A(new_n661), .B(KEYINPUT39), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n618), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n558), .A2(new_n597), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n654), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n501), .A2(new_n456), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n487), .B1(new_n445), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(G472), .B1(new_n675), .B2(G902), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n673), .B1(new_n495), .B2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n313), .B1(new_n668), .B2(KEYINPUT40), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n635), .A2(new_n636), .ZN(new_n679));
  XOR2_X1   g493(.A(new_n679), .B(KEYINPUT38), .Z(new_n680));
  NAND4_X1  g494(.A1(new_n672), .A2(new_n677), .A3(new_n678), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G143), .ZN(G45));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n633), .B2(new_n661), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n558), .A2(new_n630), .A3(KEYINPUT96), .A4(new_n662), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n686), .A2(new_n390), .A3(new_n659), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G146), .ZN(G48));
  INV_X1    g502(.A(KEYINPUT97), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n689), .B1(new_n296), .B2(G902), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n613), .A2(KEYINPUT97), .A3(new_n188), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n691), .A3(G469), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(KEYINPUT98), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n615), .A2(new_n616), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT98), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n690), .A2(new_n691), .A3(new_n695), .A4(G469), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n693), .A2(new_n311), .A3(new_n694), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n698), .A2(new_n507), .A3(new_n638), .ZN(new_n699));
  XNOR2_X1  g513(.A(KEYINPUT41), .B(G113), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n699), .B(new_n700), .ZN(G15));
  NAND3_X1  g515(.A1(new_n698), .A2(new_n507), .A3(new_n645), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G116), .ZN(G18));
  NAND4_X1  g517(.A1(new_n698), .A2(new_n659), .A3(new_n389), .A4(new_n598), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NOR2_X1   g519(.A1(new_n697), .A2(new_n637), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT100), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n601), .B2(G472), .ZN(new_n708));
  INV_X1    g522(.A(G472), .ZN(new_n709));
  AOI211_X1 g523(.A(KEYINPUT100), .B(new_n709), .C1(new_n489), .C2(new_n188), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n502), .A2(KEYINPUT99), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT99), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n712), .B(new_n501), .C1(new_n457), .C2(new_n459), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n711), .A2(new_n445), .A3(new_n713), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n714), .B(new_n483), .C1(new_n487), .C2(new_n488), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n715), .A2(new_n490), .ZN(new_n716));
  NOR4_X1   g530(.A1(new_n708), .A2(new_n710), .A3(new_n439), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n706), .A2(new_n717), .A3(new_n670), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  OAI21_X1  g533(.A(new_n312), .B1(new_n635), .B2(new_n636), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n697), .A2(new_n720), .ZN(new_n721));
  NOR4_X1   g535(.A1(new_n708), .A2(new_n710), .A3(new_n654), .A4(new_n716), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n721), .A2(new_n722), .A3(new_n686), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G125), .ZN(G27));
  INV_X1    g538(.A(KEYINPUT103), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n493), .B1(new_n489), .B2(new_n490), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n489), .A2(new_n493), .A3(new_n490), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n506), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n619), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n189), .B(KEYINPUT101), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n294), .B(new_n730), .C1(new_n297), .C2(new_n306), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n610), .A2(new_n313), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n635), .A2(new_n636), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(KEYINPUT102), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT102), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n731), .A2(new_n734), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n729), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT42), .B1(new_n739), .B2(new_n686), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n731), .A2(new_n734), .A3(new_n737), .ZN(new_n741));
  AOI21_X1  g555(.A(new_n737), .B1(new_n731), .B2(new_n734), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n686), .B(new_n507), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n725), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n739), .A2(KEYINPUT42), .A3(new_n686), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n743), .A2(new_n744), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(KEYINPUT103), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G131), .ZN(G33));
  NAND2_X1  g565(.A1(new_n739), .A2(new_n663), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G134), .ZN(G36));
  OR2_X1    g567(.A1(new_n293), .A2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n293), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT46), .B1(new_n756), .B2(new_n730), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n757), .B1(new_n616), .B2(new_n615), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n730), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n610), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  AND2_X1   g574(.A1(new_n760), .A2(new_n667), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n635), .A2(new_n636), .A3(new_n313), .ZN(new_n762));
  XOR2_X1   g576(.A(new_n762), .B(KEYINPUT105), .Z(new_n763));
  INV_X1    g577(.A(new_n630), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n558), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(KEYINPUT43), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n609), .A2(new_n767), .A3(new_n673), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n763), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT104), .ZN(new_n772));
  AND2_X1   g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  OAI211_X1 g588(.A(new_n761), .B(new_n770), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  XOR2_X1   g590(.A(new_n760), .B(KEYINPUT47), .Z(new_n777));
  NOR3_X1   g591(.A1(new_n777), .A2(new_n685), .A3(new_n684), .ZN(new_n778));
  INV_X1    g592(.A(new_n728), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n779), .A3(new_n439), .A4(new_n762), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G140), .ZN(G42));
  NAND3_X1  g595(.A1(new_n693), .A2(new_n694), .A3(new_n696), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT49), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(KEYINPUT106), .ZN(new_n786));
  INV_X1    g600(.A(new_n680), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n495), .A2(new_n676), .ZN(new_n788));
  OAI211_X1 g602(.A(new_n788), .B(new_n619), .C1(new_n783), .C2(new_n784), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n789), .A2(new_n765), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n786), .A2(new_n787), .A3(new_n732), .A4(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n777), .B1(new_n311), .B2(new_n782), .ZN(new_n792));
  INV_X1    g606(.A(new_n763), .ZN(new_n793));
  INV_X1    g607(.A(new_n561), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n767), .A2(new_n794), .A3(new_n717), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n792), .A2(new_n793), .A3(new_n795), .ZN(new_n796));
  AND3_X1   g610(.A1(new_n783), .A2(new_n794), .A3(new_n734), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n797), .A2(new_n619), .A3(new_n788), .ZN(new_n798));
  INV_X1    g612(.A(new_n558), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n798), .A2(new_n799), .A3(new_n764), .ZN(new_n800));
  XOR2_X1   g614(.A(new_n800), .B(KEYINPUT113), .Z(new_n801));
  NAND3_X1  g615(.A1(new_n797), .A2(new_n722), .A3(new_n767), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n796), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n795), .A2(new_n313), .A3(new_n787), .A4(new_n698), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(KEYINPUT111), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT50), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(KEYINPUT51), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n747), .A2(new_n748), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n718), .A2(new_n704), .A3(new_n699), .A4(new_n702), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n808), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT110), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n618), .A2(new_n389), .A3(new_n598), .A4(new_n673), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n599), .B1(new_n816), .B2(new_n609), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n799), .A2(new_n630), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n558), .A2(new_n597), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n389), .A3(new_n564), .A4(new_n819), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n609), .A2(new_n620), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n817), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n708), .A2(new_n710), .A3(new_n716), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n686), .B(new_n823), .C1(new_n741), .C2(new_n742), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n597), .A2(new_n661), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n825), .B1(new_n495), .B2(new_n506), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n643), .A2(new_n632), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n826), .A2(new_n762), .A3(new_n618), .A4(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n673), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n822), .A2(new_n830), .A3(KEYINPUT53), .A4(new_n752), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n671), .A2(new_n720), .A3(new_n662), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(new_n677), .A3(new_n311), .A4(new_n731), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n723), .A2(new_n833), .A3(new_n664), .A4(new_n687), .ZN(new_n834));
  XNOR2_X1  g648(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n834), .A2(KEYINPUT107), .A3(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n834), .A2(KEYINPUT107), .ZN(new_n837));
  INV_X1    g651(.A(new_n835), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n831), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  OAI211_X1 g654(.A(KEYINPUT110), .B(new_n808), .C1(new_n811), .C2(new_n812), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n815), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  XNOR2_X1  g658(.A(new_n834), .B(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n307), .A2(new_n619), .A3(new_n311), .ZN(new_n846));
  INV_X1    g660(.A(new_n820), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n649), .A2(new_n491), .A3(new_n846), .A4(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n656), .A3(new_n599), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n654), .B1(new_n824), .B2(new_n828), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n849), .A2(new_n850), .A3(new_n809), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n845), .A2(new_n750), .A3(new_n851), .A4(new_n752), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n842), .A2(new_n843), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  AND3_X1   g670(.A1(new_n750), .A2(new_n851), .A3(new_n752), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT53), .B1(new_n839), .B2(new_n836), .ZN(new_n858));
  AOI22_X1  g672(.A1(new_n857), .A2(new_n858), .B1(new_n852), .B2(KEYINPUT53), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(KEYINPUT54), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n795), .A2(new_n721), .ZN(new_n861));
  OAI211_X1 g675(.A(new_n861), .B(new_n559), .C1(new_n634), .C2(new_n798), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT114), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n862), .A2(new_n863), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n797), .A2(new_n507), .A3(new_n767), .ZN(new_n866));
  AOI22_X1  g680(.A1(new_n864), .A2(new_n865), .B1(KEYINPUT48), .B2(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n807), .A2(new_n856), .A3(new_n860), .A4(new_n867), .ZN(new_n868));
  XOR2_X1   g682(.A(new_n806), .B(KEYINPUT112), .Z(new_n869));
  AOI21_X1  g683(.A(KEYINPUT51), .B1(new_n869), .B2(new_n803), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n866), .A2(KEYINPUT48), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n868), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(G952), .A2(G953), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n791), .B1(new_n872), .B2(new_n873), .ZN(G75));
  INV_X1    g688(.A(KEYINPUT116), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT56), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n842), .A2(new_n854), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(G902), .ZN(new_n878));
  INV_X1    g692(.A(G210), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n875), .B(new_n876), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n343), .A2(new_n345), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT115), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n357), .B(KEYINPUT55), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n880), .A2(new_n882), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n885), .B1(new_n884), .B2(new_n886), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n285), .A2(G952), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  INV_X1    g704(.A(KEYINPUT119), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n730), .B(KEYINPUT57), .Z(new_n892));
  AOI21_X1  g706(.A(new_n843), .B1(new_n842), .B2(new_n854), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n892), .B1(new_n855), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT117), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(KEYINPUT117), .B(new_n892), .C1(new_n855), .C2(new_n893), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n296), .B(KEYINPUT118), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AND4_X1   g713(.A1(new_n891), .A2(new_n896), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n898), .B1(new_n894), .B2(new_n895), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n891), .B1(new_n901), .B2(new_n897), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n878), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n756), .B(KEYINPUT120), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n889), .B1(new_n903), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n904), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n542), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n889), .ZN(G60));
  NOR2_X1   g724(.A1(new_n855), .A2(new_n893), .ZN(new_n911));
  INV_X1    g725(.A(new_n627), .ZN(new_n912));
  INV_X1    g726(.A(new_n628), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  NOR3_X1   g730(.A1(new_n911), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n916), .B1(new_n856), .B2(new_n860), .ZN(new_n918));
  INV_X1    g732(.A(new_n914), .ZN(new_n919));
  OR3_X1    g733(.A1(new_n918), .A2(KEYINPUT121), .A3(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT121), .B1(new_n918), .B2(new_n919), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n889), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(G63));
  INV_X1    g736(.A(new_n889), .ZN(new_n923));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n842), .B2(new_n854), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n923), .B1(new_n926), .B2(new_n427), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n652), .B(KEYINPUT122), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n927), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(KEYINPUT61), .ZN(G66));
  INV_X1    g744(.A(new_n562), .ZN(new_n931));
  OAI21_X1  g745(.A(G953), .B1(new_n931), .B2(new_n355), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n849), .A2(new_n809), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n933), .B2(G953), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n882), .B1(G898), .B2(new_n285), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n934), .B(new_n935), .ZN(G69));
  AOI21_X1  g750(.A(new_n285), .B1(G227), .B2(G900), .ZN(new_n937));
  AND3_X1   g751(.A1(new_n723), .A2(new_n664), .A3(new_n687), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n681), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT62), .Z(new_n940));
  NAND2_X1  g754(.A1(new_n818), .A2(new_n819), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n668), .B1(KEYINPUT123), .B2(new_n942), .ZN(new_n943));
  OR2_X1    g757(.A1(new_n942), .A2(KEYINPUT123), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n943), .A2(new_n507), .A3(new_n762), .A4(new_n944), .ZN(new_n945));
  NAND4_X1  g759(.A1(new_n780), .A2(new_n940), .A3(new_n775), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n937), .B1(new_n946), .B2(new_n285), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n486), .B(new_n522), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n780), .A2(new_n775), .ZN(new_n951));
  NAND4_X1  g765(.A1(new_n761), .A2(new_n507), .A3(new_n389), .A4(new_n670), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n750), .A2(new_n752), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT124), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n951), .A2(new_n938), .A3(new_n952), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n948), .B1(new_n955), .B2(new_n285), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n957), .A2(G900), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n957), .A2(G900), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n937), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n950), .B1(new_n956), .B2(new_n960), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n961), .B(KEYINPUT126), .ZN(G72));
  NAND2_X1  g776(.A1(G472), .A2(G902), .ZN(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT63), .Z(new_n964));
  OAI211_X1 g778(.A(new_n859), .B(new_n964), .C1(new_n487), .C2(new_n499), .ZN(new_n965));
  INV_X1    g779(.A(new_n933), .ZN(new_n966));
  OR2_X1    g780(.A1(new_n946), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(KEYINPUT127), .A3(new_n964), .ZN(new_n968));
  INV_X1    g782(.A(new_n498), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n968), .A2(new_n444), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT127), .B1(new_n967), .B2(new_n964), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n923), .B(new_n965), .C1(new_n970), .C2(new_n971), .ZN(new_n972));
  OR2_X1    g786(.A1(new_n955), .A2(new_n966), .ZN(new_n973));
  AOI211_X1 g787(.A(new_n444), .B(new_n969), .C1(new_n973), .C2(new_n964), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n972), .A2(new_n974), .ZN(G57));
endmodule


