//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 0 0 0 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:40 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  INV_X1    g003(.A(G104), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G107), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT3), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G101), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n196), .B1(new_n192), .B2(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n190), .A2(KEYINPUT73), .A3(G107), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n194), .A2(new_n195), .A3(new_n197), .A4(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT74), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n197), .A2(new_n198), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT74), .ZN(new_n202));
  NAND4_X1  g016(.A1(new_n201), .A2(new_n202), .A3(new_n195), .A4(new_n194), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n200), .A2(new_n203), .ZN(new_n204));
  AOI21_X1  g018(.A(KEYINPUT75), .B1(new_n190), .B2(G107), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n190), .A2(G107), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n190), .A2(KEYINPUT75), .A3(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n195), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT5), .ZN(new_n211));
  INV_X1    g025(.A(G119), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G116), .ZN(new_n213));
  XNOR2_X1  g027(.A(new_n213), .B(KEYINPUT76), .ZN(new_n214));
  INV_X1    g028(.A(G113), .ZN(new_n215));
  XNOR2_X1  g029(.A(G116), .B(G119), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n215), .B1(new_n216), .B2(KEYINPUT5), .ZN(new_n217));
  XOR2_X1   g031(.A(KEYINPUT2), .B(G113), .Z(new_n218));
  AOI22_X1  g032(.A1(new_n214), .A2(new_n217), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n204), .A2(new_n210), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT4), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n191), .A2(new_n193), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n197), .A2(new_n198), .ZN(new_n223));
  OAI211_X1 g037(.A(new_n221), .B(G101), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  XOR2_X1   g038(.A(G116), .B(G119), .Z(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT2), .B(G113), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n216), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n195), .B1(new_n201), .B2(new_n194), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n231), .A2(new_n221), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n230), .B1(new_n204), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n188), .B1(new_n220), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n209), .B1(new_n200), .B2(new_n203), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(new_n219), .ZN(new_n236));
  OAI21_X1  g050(.A(G101), .B1(new_n222), .B2(new_n223), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n203), .B2(new_n200), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n236), .B(KEYINPUT77), .C1(new_n239), .C2(new_n230), .ZN(new_n240));
  XNOR2_X1  g054(.A(G110), .B(G122), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT6), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n204), .A2(new_n232), .ZN(new_n245));
  INV_X1    g059(.A(new_n230), .ZN(new_n246));
  AOI22_X1  g060(.A1(new_n245), .A2(new_n246), .B1(new_n235), .B2(new_n219), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n244), .B1(new_n247), .B2(new_n241), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G143), .ZN(new_n251));
  INV_X1    g065(.A(G143), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G146), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT0), .A2(G128), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(new_n253), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G143), .B(G146), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT0), .B(G128), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n255), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(G125), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT68), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G125), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n251), .A2(new_n253), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n251), .A2(KEYINPUT1), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n266), .A2(new_n267), .A3(G128), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n251), .B(new_n253), .C1(KEYINPUT1), .C2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n265), .B1(new_n271), .B2(new_n264), .ZN(new_n272));
  INV_X1    g086(.A(G953), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G224), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT78), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n272), .B(new_n275), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n234), .A2(new_n240), .A3(new_n244), .A4(new_n242), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n249), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n247), .A2(new_n241), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n275), .A2(KEYINPUT7), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n272), .B(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n241), .B(KEYINPUT8), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n235), .A2(new_n219), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n283), .B1(new_n220), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(G902), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n187), .B1(new_n278), .B2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n287), .A2(KEYINPUT79), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT79), .ZN(new_n289));
  AOI211_X1 g103(.A(new_n289), .B(new_n187), .C1(new_n278), .C2(new_n286), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n278), .A2(new_n286), .A3(new_n187), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(G469), .ZN(new_n293));
  INV_X1    g107(.A(G902), .ZN(new_n294));
  INV_X1    g108(.A(new_n271), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n204), .A2(new_n295), .A3(new_n210), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT10), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n258), .B1(new_n231), .B2(new_n221), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n245), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT11), .ZN(new_n301));
  INV_X1    g115(.A(G134), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(G137), .ZN(new_n303));
  INV_X1    g117(.A(G137), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n304), .A2(KEYINPUT11), .A3(G134), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n302), .A2(G137), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G131), .ZN(new_n308));
  INV_X1    g122(.A(G131), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n303), .A2(new_n305), .A3(new_n309), .A4(new_n306), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n235), .A2(KEYINPUT10), .A3(new_n295), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n298), .A2(new_n300), .A3(new_n312), .A4(new_n313), .ZN(new_n314));
  XNOR2_X1  g128(.A(G110), .B(G140), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n273), .A2(G227), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n314), .A2(new_n318), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n235), .A2(new_n295), .ZN(new_n320));
  AOI211_X1 g134(.A(new_n209), .B(new_n271), .C1(new_n200), .C2(new_n203), .ZN(new_n321));
  OAI211_X1 g135(.A(KEYINPUT12), .B(new_n311), .C1(new_n320), .C2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n311), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT12), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n319), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n298), .A2(new_n313), .A3(new_n300), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(new_n311), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n318), .B1(new_n328), .B2(new_n314), .ZN(new_n329));
  OAI211_X1 g143(.A(new_n293), .B(new_n294), .C1(new_n326), .C2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(G469), .A2(G902), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n314), .A2(new_n318), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(new_n328), .ZN(new_n333));
  INV_X1    g147(.A(new_n314), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(new_n322), .B2(new_n325), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n333), .B(G469), .C1(new_n335), .C2(new_n318), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n330), .A2(new_n331), .A3(new_n336), .ZN(new_n337));
  XNOR2_X1  g151(.A(KEYINPUT9), .B(G234), .ZN(new_n338));
  OAI21_X1  g152(.A(G221), .B1(new_n338), .B2(G902), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n339), .B(KEYINPUT72), .ZN(new_n340));
  NOR2_X1   g154(.A1(G475), .A2(G902), .ZN(new_n341));
  NOR2_X1   g155(.A1(G125), .A2(G140), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(G125), .A2(G140), .ZN(new_n344));
  AOI21_X1  g158(.A(G146), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n342), .B1(new_n264), .B2(G140), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n345), .B1(new_n346), .B2(G146), .ZN(new_n347));
  NAND2_X1  g161(.A1(KEYINPUT18), .A2(G131), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  NOR2_X1   g163(.A1(G237), .A2(G953), .ZN(new_n350));
  AND3_X1   g164(.A1(new_n350), .A2(G143), .A3(G214), .ZN(new_n351));
  AOI21_X1  g165(.A(G143), .B1(new_n350), .B2(G214), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n349), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(G237), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n354), .A2(new_n273), .A3(G214), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n252), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n350), .A2(G143), .A3(G214), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n348), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n353), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT80), .B1(new_n347), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n345), .ZN(new_n361));
  XNOR2_X1  g175(.A(KEYINPUT68), .B(G125), .ZN(new_n362));
  INV_X1    g176(.A(G140), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n343), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n361), .B1(new_n364), .B2(new_n250), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT80), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n366), .A3(new_n358), .A4(new_n353), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n360), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n356), .A2(new_n309), .A3(new_n357), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT81), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND4_X1  g185(.A1(new_n356), .A2(KEYINPUT81), .A3(new_n309), .A4(new_n357), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n356), .A2(new_n357), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G131), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n371), .A2(new_n372), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n363), .B1(new_n261), .B2(new_n263), .ZN(new_n376));
  OAI21_X1  g190(.A(KEYINPUT16), .B1(new_n376), .B2(new_n342), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT16), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n264), .A2(KEYINPUT69), .A3(new_n378), .A4(new_n363), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT69), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n363), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n380), .B1(new_n362), .B2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n377), .A2(G146), .A3(new_n379), .A4(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n343), .A2(new_n344), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT19), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n250), .B(new_n386), .C1(new_n364), .C2(new_n385), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n375), .A2(new_n383), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n368), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT82), .ZN(new_n390));
  XNOR2_X1  g204(.A(G113), .B(G122), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n190), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n389), .A2(new_n390), .A3(new_n393), .ZN(new_n394));
  OAI211_X1 g208(.A(new_n379), .B(new_n382), .C1(new_n346), .C2(new_n378), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(new_n250), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT17), .ZN(new_n397));
  NAND4_X1  g211(.A1(new_n371), .A2(new_n374), .A3(new_n397), .A4(new_n372), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n373), .A2(KEYINPUT17), .A3(G131), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n396), .A2(new_n398), .A3(new_n383), .A4(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n368), .A3(new_n392), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n390), .B1(new_n389), .B2(new_n393), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n341), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT20), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n383), .A2(new_n387), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n406), .A2(new_n375), .B1(new_n360), .B2(new_n367), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT82), .B1(new_n407), .B2(new_n392), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n401), .A3(new_n394), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT20), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(new_n341), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n400), .A2(new_n368), .A3(new_n392), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n392), .B1(new_n400), .B2(new_n368), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n294), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT83), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G475), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n400), .A2(new_n368), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n393), .ZN(new_n419));
  AOI21_X1  g233(.A(G902), .B1(new_n419), .B2(new_n401), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n417), .B1(new_n420), .B2(KEYINPUT83), .ZN(new_n421));
  AOI22_X1  g235(.A1(new_n405), .A2(new_n411), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G116), .ZN(new_n423));
  NOR2_X1   g237(.A1(new_n423), .A2(G122), .ZN(new_n424));
  INV_X1    g238(.A(G122), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n425), .A2(G116), .ZN(new_n426));
  OR3_X1    g240(.A1(new_n424), .A2(new_n426), .A3(G107), .ZN(new_n427));
  OAI21_X1  g241(.A(G107), .B1(new_n424), .B2(new_n426), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT84), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n430), .B1(new_n252), .B2(G128), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n269), .A2(KEYINPUT84), .A3(G143), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n252), .A2(G128), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT13), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n252), .A2(KEYINPUT13), .A3(G128), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n433), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G134), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n302), .A3(new_n434), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n429), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(KEYINPUT14), .B1(new_n425), .B2(G116), .ZN(new_n442));
  OAI21_X1  g256(.A(KEYINPUT85), .B1(new_n442), .B2(new_n426), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n423), .A2(G122), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n444), .B(new_n445), .C1(new_n424), .C2(KEYINPUT14), .ZN(new_n446));
  OR2_X1    g260(.A1(new_n445), .A2(KEYINPUT14), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n443), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G107), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n433), .A2(new_n302), .A3(new_n434), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n302), .B1(new_n433), .B2(new_n434), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n427), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n441), .B1(new_n450), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(G217), .ZN(new_n455));
  NOR3_X1   g269(.A1(new_n338), .A2(new_n455), .A3(G953), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n441), .B(new_n456), .C1(new_n450), .C2(new_n453), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(new_n294), .ZN(new_n461));
  INV_X1    g275(.A(G478), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT86), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(KEYINPUT15), .ZN(new_n464));
  INV_X1    g278(.A(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n463), .A2(KEYINPUT15), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n461), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n467), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n469), .B1(new_n460), .B2(new_n294), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n273), .A2(G952), .ZN(new_n471));
  NAND2_X1  g285(.A1(G234), .A2(G237), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XOR2_X1   g287(.A(new_n473), .B(KEYINPUT87), .Z(new_n474));
  AND3_X1   g288(.A1(new_n472), .A2(G902), .A3(G953), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT21), .B(G898), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n478), .B(KEYINPUT88), .Z(new_n479));
  NOR3_X1   g293(.A1(new_n468), .A2(new_n470), .A3(new_n479), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n337), .A2(new_n340), .A3(new_n422), .A4(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G214), .B1(G237), .B2(G902), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NOR3_X1   g297(.A1(new_n292), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n455), .B1(G234), .B2(new_n294), .ZN(new_n485));
  AOI21_X1  g299(.A(KEYINPUT23), .B1(new_n269), .B2(G119), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n269), .A2(G119), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n269), .A2(KEYINPUT23), .A3(G119), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G110), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT24), .B(G110), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT67), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n493), .B1(new_n269), .B2(G119), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n212), .A2(KEYINPUT67), .A3(G128), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n269), .A2(G119), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n491), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n379), .A2(new_n382), .ZN(new_n500));
  AOI21_X1  g314(.A(G146), .B1(new_n500), .B2(new_n377), .ZN(new_n501));
  INV_X1    g315(.A(new_n383), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT70), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n488), .A2(new_n504), .A3(new_n505), .A4(new_n489), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT23), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n507), .B1(new_n212), .B2(G128), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n212), .A2(G128), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(new_n489), .A3(new_n505), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT70), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n497), .A2(new_n492), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n511), .A3(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n383), .A2(new_n513), .A3(new_n361), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n273), .A2(G221), .A3(G234), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT71), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT22), .B(G137), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n516), .B(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n503), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n518), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n498), .B1(new_n396), .B2(new_n383), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n383), .A2(new_n513), .A3(new_n361), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(KEYINPUT25), .B1(new_n524), .B2(new_n294), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT25), .ZN(new_n526));
  AOI211_X1 g340(.A(new_n526), .B(G902), .C1(new_n519), .C2(new_n523), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n485), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n485), .A2(G902), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT32), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n311), .A2(new_n259), .ZN(new_n533));
  INV_X1    g347(.A(new_n229), .ZN(new_n534));
  INV_X1    g348(.A(new_n306), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n302), .A2(G137), .ZN(new_n536));
  OAI21_X1  g350(.A(G131), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND4_X1  g351(.A1(new_n268), .A2(new_n537), .A3(new_n310), .A4(new_n270), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n533), .A2(new_n534), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT64), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n350), .A2(G210), .ZN(new_n541));
  XNOR2_X1  g355(.A(new_n541), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT26), .B(G101), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n542), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT64), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n533), .A2(new_n545), .A3(new_n534), .A4(new_n538), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n540), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n547), .A2(KEYINPUT65), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT65), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n540), .A2(new_n549), .A3(new_n544), .A4(new_n546), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n533), .A2(new_n538), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT30), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT30), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n553), .B1(new_n533), .B2(new_n538), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n229), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g370(.A(KEYINPUT31), .B1(new_n548), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n229), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n540), .A2(new_n546), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n559), .A2(KEYINPUT28), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT28), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n539), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n544), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n557), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n547), .A2(KEYINPUT65), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT31), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n567), .A2(new_n568), .A3(new_n555), .A4(new_n550), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT66), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n550), .A2(new_n555), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT66), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n571), .A2(new_n572), .A3(new_n568), .A4(new_n567), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n566), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(G472), .A2(G902), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n532), .B1(new_n574), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n570), .A2(new_n573), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n571), .A2(new_n567), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n579), .A2(KEYINPUT31), .B1(new_n564), .B2(new_n563), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n576), .A2(new_n532), .ZN(new_n582));
  INV_X1    g396(.A(new_n562), .ZN(new_n583));
  AOI211_X1 g397(.A(new_n564), .B(new_n583), .C1(new_n559), .C2(KEYINPUT28), .ZN(new_n584));
  AOI21_X1  g398(.A(G902), .B1(new_n584), .B2(KEYINPUT29), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n555), .A2(new_n540), .A3(new_n546), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(new_n564), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n560), .A2(new_n544), .A3(new_n562), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n585), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n581), .A2(new_n582), .B1(G472), .B2(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n531), .B1(new_n577), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n484), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n594), .B(G101), .ZN(G3));
  INV_X1    g409(.A(new_n531), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n576), .B1(new_n578), .B2(new_n580), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n574), .A2(G902), .ZN(new_n599));
  INV_X1    g413(.A(G472), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n596), .B(new_n598), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n337), .A2(new_n340), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  INV_X1    g417(.A(new_n479), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n482), .B(new_n604), .C1(new_n291), .C2(new_n287), .ZN(new_n605));
  OAI211_X1 g419(.A(KEYINPUT83), .B(new_n294), .C1(new_n412), .C2(new_n413), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n416), .A2(G475), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n411), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n410), .B1(new_n409), .B2(new_n341), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n607), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT33), .ZN(new_n611));
  INV_X1    g425(.A(new_n459), .ZN(new_n612));
  INV_X1    g426(.A(new_n452), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n613), .A2(new_n440), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n614), .A2(new_n449), .A3(new_n427), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n456), .B1(new_n615), .B2(new_n441), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n611), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT89), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT90), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n458), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n616), .A2(KEYINPUT90), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n459), .A2(KEYINPUT33), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT89), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n460), .A2(new_n624), .A3(new_n611), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n462), .A2(G902), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n618), .A2(new_n623), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n461), .A2(new_n462), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n610), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g445(.A(KEYINPUT91), .B1(new_n605), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n278), .A2(new_n286), .ZN(new_n633));
  INV_X1    g447(.A(new_n187), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n278), .A2(new_n286), .A3(new_n187), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n483), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n405), .A2(new_n411), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n629), .B1(new_n638), .B2(new_n607), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT91), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n637), .A2(new_n639), .A3(new_n640), .A4(new_n604), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n632), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n603), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT34), .B(G104), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G6));
  INV_X1    g459(.A(KEYINPUT92), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n607), .A2(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n421), .A2(KEYINPUT92), .A3(new_n416), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  OR2_X1    g463(.A1(new_n468), .A2(new_n470), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n649), .A2(new_n638), .A3(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n605), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n603), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(new_n192), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  NOR2_X1   g470(.A1(new_n518), .A2(KEYINPUT36), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT94), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n503), .B2(new_n514), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n521), .A2(new_n522), .A3(KEYINPUT94), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n503), .A2(new_n659), .A3(new_n514), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT94), .B1(new_n521), .B2(new_n522), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(new_n664), .A3(new_n657), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n662), .A2(new_n529), .A3(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT95), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n662), .A2(KEYINPUT95), .A3(new_n529), .A4(new_n665), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n528), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n598), .B(new_n670), .C1(new_n599), .C2(new_n600), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT96), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n600), .B1(new_n581), .B2(new_n294), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n528), .A2(new_n668), .A3(new_n669), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n673), .A2(new_n597), .A3(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT96), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n672), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n484), .ZN(new_n679));
  XNOR2_X1  g493(.A(KEYINPUT37), .B(G110), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n680), .B(KEYINPUT97), .Z(new_n681));
  XNOR2_X1  g495(.A(new_n679), .B(new_n681), .ZN(G12));
  NOR2_X1   g496(.A1(new_n602), .A2(new_n674), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n577), .A2(new_n592), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n475), .A2(new_n686), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n474), .A2(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(new_n688), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n649), .A2(new_n638), .A3(new_n650), .A4(new_n689), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n482), .B1(new_n291), .B2(new_n287), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n685), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G128), .ZN(G30));
  NAND2_X1  g508(.A1(new_n635), .A2(new_n289), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n287), .A2(KEYINPUT79), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n636), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n610), .A2(new_n650), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n483), .A3(new_n670), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n688), .B(KEYINPUT39), .Z(new_n702));
  NAND3_X1  g516(.A1(new_n337), .A2(new_n340), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n701), .B1(KEYINPUT40), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n581), .A2(new_n582), .ZN(new_n705));
  AOI22_X1  g519(.A1(new_n571), .A2(new_n567), .B1(new_n564), .B2(new_n559), .ZN(new_n706));
  OAI21_X1  g520(.A(G472), .B1(new_n706), .B2(G902), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n577), .A2(new_n705), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n703), .A2(KEYINPUT40), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OR3_X1    g524(.A1(new_n699), .A2(new_n704), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n610), .A2(new_n630), .A3(new_n689), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n691), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n685), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  NAND2_X1  g530(.A1(new_n325), .A2(new_n322), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n332), .A2(new_n717), .ZN(new_n718));
  AOI22_X1  g532(.A1(new_n296), .A2(new_n297), .B1(new_n245), .B2(new_n299), .ZN(new_n719));
  AOI21_X1  g533(.A(new_n312), .B1(new_n719), .B2(new_n313), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n317), .B1(new_n720), .B2(new_n334), .ZN(new_n721));
  AOI21_X1  g535(.A(G902), .B1(new_n718), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(KEYINPUT99), .B1(new_n722), .B2(new_n293), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n328), .A2(new_n314), .ZN(new_n725));
  AOI22_X1  g539(.A1(new_n725), .A2(new_n317), .B1(new_n332), .B2(new_n717), .ZN(new_n726));
  OAI211_X1 g540(.A(new_n724), .B(G469), .C1(new_n726), .C2(G902), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n723), .A2(new_n727), .ZN(new_n728));
  AND2_X1   g542(.A1(new_n330), .A2(new_n339), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT100), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT100), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n728), .A2(new_n732), .A3(new_n729), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n731), .A2(new_n593), .A3(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n632), .A2(new_n641), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT101), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n733), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n732), .B1(new_n728), .B2(new_n729), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT101), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n739), .A2(new_n740), .A3(new_n593), .A4(new_n642), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT41), .B(G113), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(KEYINPUT102), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n742), .B(new_n744), .ZN(G15));
  NAND4_X1  g559(.A1(new_n731), .A2(new_n593), .A3(new_n652), .A4(new_n733), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G116), .ZN(G18));
  OAI211_X1 g561(.A(new_n607), .B(new_n480), .C1(new_n608), .C2(new_n609), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n674), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n591), .A2(G472), .ZN(new_n750));
  INV_X1    g564(.A(new_n582), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n750), .B1(new_n574), .B2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT32), .B1(new_n581), .B2(new_n575), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n749), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n728), .A2(new_n637), .A3(new_n729), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT103), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n728), .A2(new_n637), .A3(new_n729), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n422), .A2(new_n670), .A3(new_n480), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n577), .B2(new_n592), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT103), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n212), .ZN(G21));
  NOR3_X1   g577(.A1(new_n673), .A2(new_n597), .A3(new_n531), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n605), .A2(new_n700), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n731), .A2(new_n764), .A3(new_n733), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  INV_X1    g581(.A(new_n713), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n757), .A2(new_n675), .A3(new_n768), .ZN(new_n769));
  XOR2_X1   g583(.A(KEYINPUT104), .B(G125), .Z(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G27));
  AND2_X1   g585(.A1(new_n636), .A2(new_n482), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n695), .A2(new_n772), .A3(new_n696), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT105), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n695), .A2(new_n772), .A3(KEYINPUT105), .A4(new_n696), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n337), .A2(new_n339), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n775), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n684), .A2(new_n596), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT106), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT106), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n593), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n778), .A2(new_n780), .A3(new_n768), .A4(new_n782), .ZN(new_n783));
  AND4_X1   g597(.A1(new_n593), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n713), .A2(KEYINPUT42), .ZN(new_n785));
  AOI22_X1  g599(.A1(new_n783), .A2(KEYINPUT42), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G131), .ZN(G33));
  INV_X1    g601(.A(new_n690), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G134), .ZN(G36));
  OAI21_X1  g604(.A(new_n333), .B1(new_n335), .B2(new_n318), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT45), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n293), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n792), .B2(new_n791), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT46), .B1(new_n794), .B2(new_n331), .ZN(new_n795));
  INV_X1    g609(.A(new_n330), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n794), .A2(KEYINPUT46), .A3(new_n331), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(new_n339), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n702), .ZN(new_n801));
  XNOR2_X1  g615(.A(KEYINPUT107), .B(KEYINPUT108), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n801), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n800), .A2(new_n702), .A3(new_n802), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n775), .A2(new_n776), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT109), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT43), .B1(new_n422), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n422), .A2(new_n630), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n810), .B(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n670), .C1(new_n597), .C2(new_n673), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  XOR2_X1   g631(.A(KEYINPUT110), .B(G137), .Z(new_n818));
  XNOR2_X1  g632(.A(new_n817), .B(new_n818), .ZN(G39));
  NAND2_X1  g633(.A1(new_n799), .A2(new_n339), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT47), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n684), .A2(new_n596), .A3(new_n713), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n807), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G140), .ZN(G42));
  NAND2_X1  g639(.A1(new_n766), .A2(new_n746), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n762), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n780), .A2(new_n782), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n775), .A2(new_n768), .A3(new_n776), .A4(new_n777), .ZN(new_n829));
  OAI21_X1  g643(.A(KEYINPUT42), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n784), .A2(new_n785), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n827), .A2(new_n742), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT113), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n684), .B(new_n683), .C1(new_n692), .C2(new_n714), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n691), .A2(new_n700), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n670), .A2(new_n688), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n708), .A2(new_n777), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n834), .A2(new_n769), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n834), .A2(KEYINPUT52), .A3(new_n837), .A4(new_n769), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n671), .A2(new_n713), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n784), .A2(new_n788), .B1(new_n778), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n649), .A2(new_n638), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n845), .A2(new_n650), .A3(new_n688), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n775), .A3(new_n776), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT112), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT112), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n846), .A2(new_n775), .A3(new_n849), .A4(new_n776), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n848), .A2(new_n685), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n844), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n422), .A2(new_n650), .ZN(new_n853));
  NOR4_X1   g667(.A1(new_n292), .A2(new_n483), .A3(new_n479), .A4(new_n853), .ZN(new_n854));
  AOI22_X1  g668(.A1(new_n854), .A2(new_n603), .B1(new_n484), .B2(new_n593), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n288), .A2(new_n290), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n483), .B1(new_n856), .B2(new_n636), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n857), .A2(KEYINPUT111), .A3(new_n604), .A4(new_n639), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n697), .A2(new_n482), .A3(new_n604), .A4(new_n639), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT111), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n861), .A3(new_n603), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n679), .A2(new_n855), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT53), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n852), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n786), .A2(new_n866), .A3(new_n742), .A4(new_n827), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n833), .A2(new_n842), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n844), .A2(new_n851), .ZN(new_n871));
  INV_X1    g685(.A(new_n863), .ZN(new_n872));
  AND4_X1   g686(.A1(KEYINPUT53), .A2(new_n871), .A3(new_n872), .A4(new_n842), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT114), .A3(new_n833), .A4(new_n867), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n832), .A2(new_n863), .A3(new_n852), .ZN(new_n876));
  AOI21_X1  g690(.A(KEYINPUT53), .B1(new_n876), .B2(new_n842), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n880));
  INV_X1    g694(.A(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n827), .A2(new_n742), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n873), .A2(new_n786), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(new_n474), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n812), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n889), .A2(new_n601), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n730), .A2(new_n482), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n699), .A3(new_n891), .ZN(new_n892));
  XOR2_X1   g706(.A(new_n892), .B(KEYINPUT50), .Z(new_n893));
  NAND2_X1  g707(.A1(new_n728), .A2(new_n330), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n340), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n807), .B(new_n890), .C1(new_n822), .C2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n730), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n807), .A2(new_n897), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n898), .B(KEYINPUT116), .ZN(new_n899));
  INV_X1    g713(.A(new_n889), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n899), .A2(new_n675), .A3(new_n900), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n893), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n708), .A2(new_n531), .A3(new_n474), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n899), .A2(new_n903), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT117), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n904), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n422), .A2(new_n629), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n902), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n890), .A2(new_n757), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n910), .A2(new_n471), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n906), .B2(new_n631), .ZN(new_n912));
  AOI22_X1  g726(.A1(new_n908), .A2(new_n909), .B1(new_n912), .B2(KEYINPUT118), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n914), .B(new_n911), .C1(new_n906), .C2(new_n631), .ZN(new_n915));
  INV_X1    g729(.A(new_n828), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n899), .A2(new_n916), .A3(new_n900), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT48), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n915), .A2(new_n918), .ZN(new_n919));
  OAI211_X1 g733(.A(new_n913), .B(new_n919), .C1(new_n909), .C2(new_n908), .ZN(new_n920));
  OAI22_X1  g734(.A1(new_n887), .A2(new_n920), .B1(G952), .B2(G953), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n894), .B(KEYINPUT49), .Z(new_n922));
  NAND3_X1  g736(.A1(new_n596), .A2(new_n482), .A3(new_n340), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n708), .A2(new_n923), .A3(new_n811), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n699), .A3(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n921), .A2(new_n925), .ZN(G75));
  NOR2_X1   g740(.A1(new_n273), .A2(G952), .ZN(new_n927));
  INV_X1    g741(.A(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT56), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n879), .A2(G902), .ZN(new_n930));
  INV_X1    g744(.A(G210), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n249), .A2(new_n277), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(new_n276), .Z(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n928), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT119), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n877), .B1(new_n870), .B2(new_n874), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n294), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT56), .B1(new_n939), .B2(G210), .ZN(new_n940));
  INV_X1    g754(.A(new_n935), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n932), .A2(KEYINPUT119), .A3(new_n935), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n936), .B1(new_n942), .B2(new_n943), .ZN(G51));
  NAND2_X1  g758(.A1(new_n879), .A2(new_n881), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT120), .B1(new_n938), .B2(new_n880), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n879), .A2(KEYINPUT120), .A3(new_n881), .ZN(new_n948));
  XOR2_X1   g762(.A(new_n331), .B(KEYINPUT57), .Z(new_n949));
  NAND3_X1  g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(new_n726), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  OR2_X1    g766(.A1(new_n930), .A2(new_n794), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n927), .B1(new_n952), .B2(new_n953), .ZN(G54));
  AND2_X1   g768(.A1(KEYINPUT58), .A2(G475), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n939), .A2(new_n409), .A3(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n409), .B1(new_n939), .B2(new_n955), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n956), .A2(new_n957), .A3(new_n927), .ZN(G60));
  NAND2_X1  g772(.A1(G478), .A2(G902), .ZN(new_n959));
  XOR2_X1   g773(.A(new_n959), .B(KEYINPUT59), .Z(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n882), .B2(new_n886), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n618), .A2(new_n625), .A3(new_n623), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n927), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n963), .A2(new_n960), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n947), .A2(new_n948), .A3(new_n965), .ZN(new_n966));
  AND2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(G63));
  NAND2_X1  g781(.A1(G217), .A2(G902), .ZN(new_n968));
  XNOR2_X1  g782(.A(new_n968), .B(KEYINPUT121), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n969), .B(KEYINPUT60), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n879), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n524), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n927), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n662), .A2(new_n665), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n973), .B1(new_n974), .B2(new_n971), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI211_X1 g791(.A(new_n973), .B(KEYINPUT61), .C1(new_n974), .C2(new_n971), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(G66));
  INV_X1    g793(.A(G224), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n476), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n883), .A2(new_n872), .ZN(new_n982));
  XOR2_X1   g796(.A(new_n982), .B(KEYINPUT122), .Z(new_n983));
  OAI21_X1  g797(.A(new_n981), .B1(new_n983), .B2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n933), .B1(G898), .B2(new_n273), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT123), .Z(new_n986));
  XNOR2_X1  g800(.A(new_n984), .B(new_n986), .ZN(G69));
  NAND2_X1  g801(.A1(new_n631), .A2(new_n853), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(KEYINPUT124), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n703), .B1(new_n988), .B2(KEYINPUT124), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n807), .A2(new_n593), .A3(new_n989), .A4(new_n990), .ZN(new_n991));
  AND2_X1   g805(.A1(new_n834), .A2(new_n769), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n711), .A2(new_n992), .ZN(new_n993));
  XOR2_X1   g807(.A(new_n993), .B(KEYINPUT62), .Z(new_n994));
  NAND4_X1  g808(.A1(new_n817), .A2(new_n824), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n273), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n552), .A2(new_n554), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n386), .B1(new_n364), .B2(new_n385), .ZN(new_n998));
  XOR2_X1   g812(.A(new_n997), .B(new_n998), .Z(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n686), .A2(G953), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1001), .B(KEYINPUT125), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n824), .A2(new_n789), .A3(new_n992), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n916), .A2(new_n835), .ZN(new_n1005));
  AND2_X1   g819(.A1(new_n816), .A2(new_n1005), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1004), .B(new_n786), .C1(new_n806), .C2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n1003), .B1(new_n1007), .B2(new_n273), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1000), .B1(new_n1008), .B2(new_n999), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n273), .B1(G227), .B2(G900), .ZN(new_n1010));
  XNOR2_X1  g824(.A(new_n1009), .B(new_n1010), .ZN(G72));
  NAND2_X1  g825(.A1(G472), .A2(G902), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT63), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1013), .B(KEYINPUT126), .ZN(new_n1014));
  INV_X1    g828(.A(new_n983), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n1015), .B2(new_n995), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1016), .A2(new_n544), .A3(new_n586), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1013), .B1(new_n579), .B2(new_n587), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n927), .B1(new_n885), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1014), .B1(new_n1015), .B2(new_n1007), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n586), .A2(new_n544), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G57));
endmodule


