

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758;

  BUF_X1 U376 ( .A(n702), .Z(n355) );
  XNOR2_X1 U377 ( .A(n371), .B(KEYINPUT1), .ZN(n702) );
  XNOR2_X1 U378 ( .A(n478), .B(n363), .ZN(n479) );
  XNOR2_X1 U379 ( .A(n362), .B(n640), .ZN(n442) );
  XNOR2_X1 U380 ( .A(n365), .B(n429), .ZN(n747) );
  XOR2_X1 U381 ( .A(G104), .B(G107), .Z(n365) );
  XNOR2_X1 U382 ( .A(G128), .B(G143), .ZN(n468) );
  INV_X1 U383 ( .A(KEYINPUT64), .ZN(n406) );
  AND2_X4 U384 ( .A1(n378), .A2(n377), .ZN(n736) );
  OR2_X2 U385 ( .A1(n660), .A2(G902), .ZN(n436) );
  XNOR2_X1 U386 ( .A(n356), .B(KEYINPUT124), .ZN(G66) );
  NOR2_X2 U387 ( .A1(n740), .A2(n739), .ZN(n356) );
  NOR2_X2 U388 ( .A1(n734), .A2(n739), .ZN(n735) );
  AND2_X2 U389 ( .A1(n384), .A2(n755), .ZN(n383) );
  XNOR2_X2 U390 ( .A(n602), .B(KEYINPUT105), .ZN(n608) );
  NOR2_X2 U391 ( .A1(n629), .A2(n739), .ZN(n631) );
  XNOR2_X1 U392 ( .A(n506), .B(KEYINPUT19), .ZN(n544) );
  NAND2_X1 U393 ( .A1(n551), .A2(n550), .ZN(n554) );
  AND2_X1 U394 ( .A1(n502), .A2(n501), .ZN(n388) );
  NOR2_X1 U395 ( .A1(n514), .A2(n490), .ZN(n481) );
  XNOR2_X1 U396 ( .A(n498), .B(n497), .ZN(n555) );
  OR2_X1 U397 ( .A1(n738), .A2(G902), .ZN(n421) );
  XNOR2_X1 U398 ( .A(n468), .B(G134), .ZN(n428) );
  XNOR2_X1 U399 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n464) );
  INV_X1 U400 ( .A(n628), .ZN(n357) );
  BUF_X1 U401 ( .A(n730), .Z(n358) );
  INV_X1 U402 ( .A(n373), .ZN(n359) );
  XNOR2_X1 U403 ( .A(n566), .B(n368), .ZN(n568) );
  NOR2_X1 U404 ( .A1(n461), .A2(n483), .ZN(n462) );
  XNOR2_X1 U405 ( .A(n493), .B(n492), .ZN(n693) );
  NAND2_X1 U406 ( .A1(n375), .A2(n374), .ZN(n377) );
  AND2_X1 U407 ( .A1(n622), .A2(KEYINPUT2), .ZN(n374) );
  NAND2_X1 U408 ( .A1(n383), .A2(n382), .ZN(n381) );
  NOR2_X1 U409 ( .A1(n522), .A2(n360), .ZN(n380) );
  XOR2_X1 U410 ( .A(KEYINPUT96), .B(KEYINPUT77), .Z(n440) );
  XNOR2_X1 U411 ( .A(G140), .B(G113), .ZN(n393) );
  XNOR2_X1 U412 ( .A(G143), .B(G104), .ZN(n389) );
  XNOR2_X1 U413 ( .A(n428), .B(n427), .ZN(n638) );
  NAND2_X1 U414 ( .A1(n479), .A2(n690), .ZN(n506) );
  XNOR2_X1 U415 ( .A(n400), .B(n399), .ZN(n516) );
  XNOR2_X1 U416 ( .A(G119), .B(G116), .ZN(n446) );
  INV_X1 U417 ( .A(G953), .ZN(n742) );
  XNOR2_X1 U418 ( .A(G110), .B(G128), .ZN(n413) );
  XOR2_X1 U419 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n403) );
  XNOR2_X1 U420 ( .A(G107), .B(G116), .ZN(n401) );
  XNOR2_X1 U421 ( .A(n408), .B(n407), .ZN(n416) );
  XNOR2_X1 U422 ( .A(G140), .B(G137), .ZN(n431) );
  XNOR2_X1 U423 ( .A(G146), .B(G125), .ZN(n467) );
  XNOR2_X1 U424 ( .A(n386), .B(n369), .ZN(n562) );
  XNOR2_X1 U425 ( .A(n412), .B(G478), .ZN(n518) );
  AND2_X1 U426 ( .A1(n513), .A2(n512), .ZN(n360) );
  OR2_X1 U427 ( .A1(n617), .A2(n616), .ZN(n361) );
  XOR2_X1 U428 ( .A(KEYINPUT70), .B(G101), .Z(n362) );
  XOR2_X1 U429 ( .A(n477), .B(KEYINPUT90), .Z(n363) );
  XOR2_X1 U430 ( .A(KEYINPUT23), .B(G119), .Z(n364) );
  AND2_X1 U431 ( .A1(G217), .A2(n424), .ZN(n366) );
  NOR2_X1 U432 ( .A1(n700), .A2(n373), .ZN(n367) );
  XOR2_X1 U433 ( .A(KEYINPUT107), .B(KEYINPUT33), .Z(n368) );
  XOR2_X1 U434 ( .A(n559), .B(KEYINPUT32), .Z(n369) );
  NAND2_X1 U435 ( .A1(n620), .A2(KEYINPUT67), .ZN(n370) );
  AND2_X1 U436 ( .A1(n371), .A2(n563), .ZN(n437) );
  XNOR2_X1 U437 ( .A(n371), .B(n487), .ZN(n488) );
  XNOR2_X2 U438 ( .A(n436), .B(G469), .ZN(n371) );
  NAND2_X1 U439 ( .A1(n359), .A2(n372), .ZN(n723) );
  INV_X1 U440 ( .A(n722), .ZN(n372) );
  INV_X1 U441 ( .A(n568), .ZN(n373) );
  NAND2_X1 U442 ( .A1(n361), .A2(n619), .ZN(n376) );
  INV_X1 U443 ( .A(n686), .ZN(n375) );
  NAND2_X1 U444 ( .A1(n376), .A2(n370), .ZN(n378) );
  INV_X1 U445 ( .A(n377), .ZN(n685) );
  NAND2_X1 U446 ( .A1(n379), .A2(KEYINPUT72), .ZN(n385) );
  NAND2_X1 U447 ( .A1(n380), .A2(n755), .ZN(n379) );
  XNOR2_X2 U448 ( .A(n504), .B(KEYINPUT114), .ZN(n755) );
  NAND2_X1 U449 ( .A1(n385), .A2(n381), .ZN(n523) );
  INV_X1 U450 ( .A(n522), .ZN(n382) );
  NOR2_X1 U451 ( .A1(n360), .A2(KEYINPUT72), .ZN(n384) );
  INV_X1 U452 ( .A(n562), .ZN(n633) );
  NAND2_X1 U453 ( .A1(n584), .A2(n558), .ZN(n386) );
  XNOR2_X2 U454 ( .A(n554), .B(n553), .ZN(n584) );
  BUF_X1 U455 ( .A(n623), .Z(n686) );
  OR2_X1 U456 ( .A1(G902), .A2(G237), .ZN(n387) );
  INV_X1 U457 ( .A(n586), .ZN(n556) );
  XNOR2_X1 U458 ( .A(n525), .B(KEYINPUT86), .ZN(n526) );
  INV_X1 U459 ( .A(KEYINPUT8), .ZN(n407) );
  INV_X1 U460 ( .A(KEYINPUT103), .ZN(n492) );
  XNOR2_X1 U461 ( .A(n415), .B(n414), .ZN(n418) );
  BUF_X1 U462 ( .A(n498), .Z(n708) );
  AND2_X1 U463 ( .A1(n583), .A2(n557), .ZN(n558) );
  NOR2_X1 U464 ( .A1(n514), .A2(n535), .ZN(n515) );
  INV_X1 U465 ( .A(KEYINPUT63), .ZN(n630) );
  XNOR2_X1 U466 ( .A(n467), .B(KEYINPUT10), .ZN(n419) );
  XNOR2_X1 U467 ( .A(KEYINPUT71), .B(G131), .ZN(n427) );
  XNOR2_X1 U468 ( .A(n427), .B(n389), .ZN(n390) );
  XNOR2_X1 U469 ( .A(n419), .B(n390), .ZN(n398) );
  XOR2_X1 U470 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n392) );
  NOR2_X1 U471 ( .A1(G953), .A2(G237), .ZN(n443) );
  NAND2_X1 U472 ( .A1(n443), .A2(G214), .ZN(n391) );
  XNOR2_X1 U473 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U474 ( .A(KEYINPUT97), .B(G122), .Z(n394) );
  XNOR2_X1 U475 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U476 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U477 ( .A(n398), .B(n397), .ZN(n651) );
  INV_X1 U478 ( .A(G902), .ZN(n457) );
  NAND2_X1 U479 ( .A1(n651), .A2(n457), .ZN(n400) );
  XNOR2_X1 U480 ( .A(KEYINPUT13), .B(G475), .ZN(n399) );
  XNOR2_X1 U481 ( .A(KEYINPUT98), .B(n516), .ZN(n509) );
  XNOR2_X1 U482 ( .A(n401), .B(KEYINPUT7), .ZN(n405) );
  XNOR2_X1 U483 ( .A(G122), .B(KEYINPUT9), .ZN(n402) );
  XNOR2_X1 U484 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U485 ( .A(n405), .B(n404), .Z(n410) );
  XNOR2_X2 U486 ( .A(n406), .B(G953), .ZN(n463) );
  NAND2_X1 U487 ( .A1(n463), .A2(G234), .ZN(n408) );
  NAND2_X1 U488 ( .A1(G217), .A2(n416), .ZN(n409) );
  XNOR2_X1 U489 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U490 ( .A(n428), .B(n411), .ZN(n649) );
  NAND2_X1 U491 ( .A1(n649), .A2(n457), .ZN(n412) );
  NOR2_X1 U492 ( .A1(n509), .A2(n518), .ZN(n676) );
  INV_X1 U493 ( .A(n676), .ZN(n679) );
  XNOR2_X1 U494 ( .A(n364), .B(n413), .ZN(n415) );
  XOR2_X1 U495 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n414) );
  NAND2_X1 U496 ( .A1(n416), .A2(G221), .ZN(n417) );
  XNOR2_X1 U497 ( .A(n418), .B(n417), .ZN(n420) );
  XNOR2_X1 U498 ( .A(n419), .B(n431), .ZN(n636) );
  XNOR2_X1 U499 ( .A(n420), .B(n636), .ZN(n738) );
  XNOR2_X2 U500 ( .A(n421), .B(KEYINPUT25), .ZN(n423) );
  XNOR2_X1 U501 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  NAND2_X1 U502 ( .A1(n618), .A2(G234), .ZN(n422) );
  XNOR2_X1 U503 ( .A(n422), .B(KEYINPUT20), .ZN(n424) );
  XNOR2_X2 U504 ( .A(n423), .B(n366), .ZN(n586) );
  NAND2_X1 U505 ( .A1(G221), .A2(n424), .ZN(n425) );
  XNOR2_X1 U506 ( .A(KEYINPUT21), .B(n425), .ZN(n705) );
  INV_X1 U507 ( .A(KEYINPUT94), .ZN(n426) );
  XNOR2_X1 U508 ( .A(n705), .B(n426), .ZN(n563) );
  XNOR2_X1 U509 ( .A(n638), .B(G146), .ZN(n450) );
  XNOR2_X2 U510 ( .A(KEYINPUT4), .B(KEYINPUT66), .ZN(n640) );
  XNOR2_X1 U511 ( .A(G110), .B(KEYINPUT78), .ZN(n429) );
  XNOR2_X1 U512 ( .A(n442), .B(n747), .ZN(n471) );
  XNOR2_X1 U513 ( .A(KEYINPUT79), .B(KEYINPUT93), .ZN(n430) );
  XNOR2_X1 U514 ( .A(n431), .B(n430), .ZN(n433) );
  NAND2_X1 U515 ( .A1(n463), .A2(G227), .ZN(n432) );
  XNOR2_X1 U516 ( .A(n433), .B(n432), .ZN(n434) );
  XNOR2_X1 U517 ( .A(n471), .B(n434), .ZN(n435) );
  XNOR2_X1 U518 ( .A(n450), .B(n435), .ZN(n660) );
  NAND2_X1 U519 ( .A1(n586), .A2(n437), .ZN(n438) );
  XNOR2_X1 U520 ( .A(n438), .B(KEYINPUT95), .ZN(n596) );
  XOR2_X1 U521 ( .A(KEYINPUT30), .B(KEYINPUT109), .Z(n455) );
  XOR2_X1 U522 ( .A(G137), .B(KEYINPUT5), .Z(n439) );
  XNOR2_X1 U523 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U524 ( .A(n442), .B(n441), .ZN(n445) );
  NAND2_X1 U525 ( .A1(n443), .A2(G210), .ZN(n444) );
  XNOR2_X1 U526 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U527 ( .A(KEYINPUT89), .B(G113), .Z(n447) );
  XNOR2_X1 U528 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U529 ( .A(n448), .B(KEYINPUT3), .ZN(n474) );
  XNOR2_X1 U530 ( .A(n449), .B(n474), .ZN(n451) );
  XNOR2_X1 U531 ( .A(n451), .B(n450), .ZN(n624) );
  NAND2_X1 U532 ( .A1(n624), .A2(n457), .ZN(n453) );
  XOR2_X1 U533 ( .A(KEYINPUT73), .B(G472), .Z(n452) );
  XNOR2_X2 U534 ( .A(n453), .B(n452), .ZN(n498) );
  XNOR2_X1 U535 ( .A(KEYINPUT76), .B(n387), .ZN(n476) );
  NAND2_X1 U536 ( .A1(n476), .A2(G214), .ZN(n690) );
  NAND2_X1 U537 ( .A1(n498), .A2(n690), .ZN(n454) );
  XNOR2_X1 U538 ( .A(n455), .B(n454), .ZN(n461) );
  NAND2_X1 U539 ( .A1(G234), .A2(G237), .ZN(n456) );
  XNOR2_X1 U540 ( .A(n456), .B(KEYINPUT14), .ZN(n718) );
  INV_X1 U541 ( .A(n463), .ZN(n628) );
  NOR2_X1 U542 ( .A1(n457), .A2(G900), .ZN(n458) );
  NAND2_X1 U543 ( .A1(n628), .A2(n458), .ZN(n459) );
  NAND2_X1 U544 ( .A1(n742), .A2(G952), .ZN(n540) );
  NAND2_X1 U545 ( .A1(n459), .A2(n540), .ZN(n460) );
  NAND2_X1 U546 ( .A1(n718), .A2(n460), .ZN(n483) );
  NAND2_X1 U547 ( .A1(n596), .A2(n462), .ZN(n514) );
  NAND2_X1 U548 ( .A1(n463), .A2(G224), .ZN(n466) );
  XNOR2_X1 U549 ( .A(n464), .B(KEYINPUT80), .ZN(n465) );
  XNOR2_X1 U550 ( .A(n466), .B(n465), .ZN(n470) );
  XNOR2_X1 U551 ( .A(n468), .B(n467), .ZN(n469) );
  XNOR2_X1 U552 ( .A(n470), .B(n469), .ZN(n472) );
  XNOR2_X1 U553 ( .A(n472), .B(n471), .ZN(n475) );
  XNOR2_X1 U554 ( .A(KEYINPUT16), .B(G122), .ZN(n473) );
  XNOR2_X1 U555 ( .A(n474), .B(n473), .ZN(n749) );
  XNOR2_X1 U556 ( .A(n475), .B(n749), .ZN(n730) );
  INV_X1 U557 ( .A(n618), .ZN(n619) );
  OR2_X2 U558 ( .A1(n730), .A2(n619), .ZN(n478) );
  NAND2_X1 U559 ( .A1(n476), .A2(G210), .ZN(n477) );
  INV_X1 U560 ( .A(n479), .ZN(n535) );
  XNOR2_X1 U561 ( .A(KEYINPUT38), .B(KEYINPUT75), .ZN(n480) );
  XNOR2_X1 U562 ( .A(n535), .B(n480), .ZN(n490) );
  XNOR2_X1 U563 ( .A(n481), .B(KEYINPUT39), .ZN(n528) );
  NOR2_X1 U564 ( .A1(n679), .A2(n528), .ZN(n482) );
  XNOR2_X1 U565 ( .A(n482), .B(KEYINPUT40), .ZN(n758) );
  XOR2_X1 U566 ( .A(KEYINPUT28), .B(KEYINPUT112), .Z(n486) );
  NOR2_X1 U567 ( .A1(n705), .A2(n483), .ZN(n484) );
  AND2_X1 U568 ( .A1(n556), .A2(n484), .ZN(n499) );
  NAND2_X1 U569 ( .A1(n499), .A2(n708), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n486), .B(n485), .ZN(n489) );
  INV_X1 U571 ( .A(KEYINPUT111), .ZN(n487) );
  NAND2_X1 U572 ( .A1(n489), .A2(n488), .ZN(n505) );
  INV_X1 U573 ( .A(n490), .ZN(n691) );
  NAND2_X1 U574 ( .A1(n691), .A2(n690), .ZN(n694) );
  INV_X1 U575 ( .A(n518), .ZN(n491) );
  NAND2_X1 U576 ( .A1(n491), .A2(n516), .ZN(n493) );
  NOR2_X1 U577 ( .A1(n694), .A2(n693), .ZN(n494) );
  XNOR2_X1 U578 ( .A(n494), .B(KEYINPUT41), .ZN(n722) );
  NOR2_X1 U579 ( .A1(n505), .A2(n722), .ZN(n495) );
  XNOR2_X1 U580 ( .A(KEYINPUT42), .B(n495), .ZN(n757) );
  NOR2_X1 U581 ( .A1(n758), .A2(n757), .ZN(n496) );
  XOR2_X1 U582 ( .A(KEYINPUT46), .B(n496), .Z(n524) );
  INV_X1 U583 ( .A(KEYINPUT6), .ZN(n497) );
  AND2_X1 U584 ( .A1(n555), .A2(n676), .ZN(n500) );
  NAND2_X1 U585 ( .A1(n500), .A2(n499), .ZN(n531) );
  XNOR2_X1 U586 ( .A(n531), .B(KEYINPUT113), .ZN(n502) );
  INV_X1 U587 ( .A(n690), .ZN(n530) );
  INV_X1 U588 ( .A(n506), .ZN(n501) );
  XNOR2_X1 U589 ( .A(n388), .B(KEYINPUT36), .ZN(n503) );
  NAND2_X1 U590 ( .A1(n503), .A2(n355), .ZN(n504) );
  INV_X1 U591 ( .A(n505), .ZN(n507) );
  NAND2_X1 U592 ( .A1(n507), .A2(n544), .ZN(n508) );
  XNOR2_X1 U593 ( .A(n508), .B(KEYINPUT47), .ZN(n513) );
  INV_X1 U594 ( .A(n508), .ZN(n677) );
  NAND2_X1 U595 ( .A1(n518), .A2(n509), .ZN(n510) );
  XNOR2_X1 U596 ( .A(n510), .B(KEYINPUT101), .ZN(n670) );
  NOR2_X1 U597 ( .A1(n670), .A2(n676), .ZN(n511) );
  XNOR2_X1 U598 ( .A(KEYINPUT102), .B(n511), .ZN(n695) );
  NAND2_X1 U599 ( .A1(n677), .A2(n695), .ZN(n512) );
  XNOR2_X1 U600 ( .A(n515), .B(KEYINPUT110), .ZN(n519) );
  INV_X1 U601 ( .A(n516), .ZN(n517) );
  AND2_X1 U602 ( .A1(n518), .A2(n517), .ZN(n571) );
  NAND2_X1 U603 ( .A1(n519), .A2(n571), .ZN(n675) );
  NAND2_X1 U604 ( .A1(n695), .A2(KEYINPUT47), .ZN(n520) );
  NAND2_X1 U605 ( .A1(n675), .A2(n520), .ZN(n521) );
  XNOR2_X1 U606 ( .A(n521), .B(KEYINPUT82), .ZN(n522) );
  NOR2_X1 U607 ( .A1(n524), .A2(n523), .ZN(n527) );
  INV_X1 U608 ( .A(KEYINPUT48), .ZN(n525) );
  XNOR2_X1 U609 ( .A(n527), .B(n526), .ZN(n538) );
  INV_X1 U610 ( .A(n670), .ZN(n682) );
  NOR2_X1 U611 ( .A1(n682), .A2(n528), .ZN(n529) );
  XNOR2_X1 U612 ( .A(n529), .B(KEYINPUT115), .ZN(n754) );
  NOR2_X1 U613 ( .A1(n531), .A2(n530), .ZN(n532) );
  INV_X1 U614 ( .A(n355), .ZN(n587) );
  NAND2_X1 U615 ( .A1(n532), .A2(n587), .ZN(n534) );
  XNOR2_X1 U616 ( .A(KEYINPUT108), .B(KEYINPUT43), .ZN(n533) );
  XNOR2_X1 U617 ( .A(n534), .B(n533), .ZN(n536) );
  NAND2_X1 U618 ( .A1(n536), .A2(n535), .ZN(n632) );
  NAND2_X1 U619 ( .A1(n754), .A2(n632), .ZN(n537) );
  OR2_X2 U620 ( .A1(n538), .A2(n537), .ZN(n621) );
  NOR2_X1 U621 ( .A1(G898), .A2(n742), .ZN(n539) );
  XOR2_X1 U622 ( .A(KEYINPUT91), .B(n539), .Z(n751) );
  NAND2_X1 U623 ( .A1(n751), .A2(G902), .ZN(n541) );
  NAND2_X1 U624 ( .A1(n541), .A2(n540), .ZN(n542) );
  AND2_X1 U625 ( .A1(n542), .A2(n718), .ZN(n543) );
  NAND2_X1 U626 ( .A1(n544), .A2(n543), .ZN(n547) );
  INV_X1 U627 ( .A(KEYINPUT69), .ZN(n545) );
  XNOR2_X1 U628 ( .A(n545), .B(KEYINPUT0), .ZN(n546) );
  XNOR2_X2 U629 ( .A(n547), .B(n546), .ZN(n592) );
  INV_X1 U630 ( .A(n592), .ZN(n551) );
  INV_X1 U631 ( .A(n563), .ZN(n548) );
  NOR2_X1 U632 ( .A1(n693), .A2(n548), .ZN(n549) );
  XNOR2_X1 U633 ( .A(n549), .B(KEYINPUT104), .ZN(n550) );
  INV_X1 U634 ( .A(KEYINPUT74), .ZN(n552) );
  XNOR2_X1 U635 ( .A(n552), .B(KEYINPUT22), .ZN(n553) );
  AND2_X1 U636 ( .A1(n556), .A2(n355), .ZN(n557) );
  INV_X1 U637 ( .A(KEYINPUT81), .ZN(n559) );
  OR2_X1 U638 ( .A1(n708), .A2(n586), .ZN(n560) );
  NOR2_X1 U639 ( .A1(n355), .A2(n560), .ZN(n561) );
  AND2_X1 U640 ( .A1(n584), .A2(n561), .ZN(n669) );
  OR2_X1 U641 ( .A1(n562), .A2(n669), .ZN(n574) );
  AND2_X1 U642 ( .A1(n586), .A2(n563), .ZN(n701) );
  NAND2_X1 U643 ( .A1(n701), .A2(n702), .ZN(n590) );
  INV_X1 U644 ( .A(KEYINPUT106), .ZN(n564) );
  XNOR2_X1 U645 ( .A(n590), .B(n564), .ZN(n565) );
  NAND2_X1 U646 ( .A1(n565), .A2(n555), .ZN(n566) );
  XNOR2_X1 U647 ( .A(n592), .B(KEYINPUT92), .ZN(n598) );
  INV_X1 U648 ( .A(n598), .ZN(n567) );
  NAND2_X1 U649 ( .A1(n568), .A2(n567), .ZN(n570) );
  INV_X1 U650 ( .A(KEYINPUT34), .ZN(n569) );
  XNOR2_X1 U651 ( .A(n570), .B(n569), .ZN(n572) );
  NAND2_X1 U652 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X2 U653 ( .A(n573), .B(KEYINPUT35), .ZN(n605) );
  NOR2_X1 U654 ( .A1(n574), .A2(n605), .ZN(n575) );
  NOR2_X1 U655 ( .A1(n575), .A2(KEYINPUT44), .ZN(n576) );
  INV_X1 U656 ( .A(n576), .ZN(n582) );
  NAND2_X1 U657 ( .A1(n605), .A2(KEYINPUT88), .ZN(n580) );
  INV_X1 U658 ( .A(KEYINPUT44), .ZN(n577) );
  NOR2_X1 U659 ( .A1(n669), .A2(n577), .ZN(n578) );
  AND2_X1 U660 ( .A1(n633), .A2(n578), .ZN(n579) );
  NAND2_X1 U661 ( .A1(n580), .A2(n579), .ZN(n581) );
  NAND2_X1 U662 ( .A1(n582), .A2(n581), .ZN(n612) );
  INV_X1 U663 ( .A(n555), .ZN(n583) );
  NAND2_X1 U664 ( .A1(n584), .A2(n583), .ZN(n585) );
  XNOR2_X1 U665 ( .A(n585), .B(KEYINPUT87), .ZN(n589) );
  AND2_X1 U666 ( .A1(n587), .A2(n586), .ZN(n588) );
  NAND2_X1 U667 ( .A1(n589), .A2(n588), .ZN(n634) );
  INV_X1 U668 ( .A(n590), .ZN(n591) );
  NAND2_X1 U669 ( .A1(n591), .A2(n708), .ZN(n712) );
  OR2_X1 U670 ( .A1(n592), .A2(n712), .ZN(n594) );
  INV_X1 U671 ( .A(KEYINPUT31), .ZN(n593) );
  XNOR2_X1 U672 ( .A(n594), .B(n593), .ZN(n681) );
  INV_X1 U673 ( .A(n708), .ZN(n595) );
  NAND2_X1 U674 ( .A1(n596), .A2(n595), .ZN(n597) );
  OR2_X1 U675 ( .A1(n598), .A2(n597), .ZN(n665) );
  NAND2_X1 U676 ( .A1(n681), .A2(n665), .ZN(n600) );
  INV_X1 U677 ( .A(n695), .ZN(n599) );
  NAND2_X1 U678 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U679 ( .A1(n634), .A2(n601), .ZN(n602) );
  INV_X1 U680 ( .A(n608), .ZN(n604) );
  INV_X1 U681 ( .A(KEYINPUT88), .ZN(n603) );
  NAND2_X1 U682 ( .A1(n604), .A2(n603), .ZN(n610) );
  NAND2_X1 U683 ( .A1(n605), .A2(KEYINPUT44), .ZN(n606) );
  NAND2_X1 U684 ( .A1(n606), .A2(n603), .ZN(n607) );
  NAND2_X1 U685 ( .A1(n608), .A2(n607), .ZN(n609) );
  NAND2_X1 U686 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(n614) );
  XNOR2_X1 U688 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n613) );
  XNOR2_X1 U689 ( .A(n614), .B(n613), .ZN(n623) );
  NOR2_X1 U690 ( .A1(n621), .A2(n623), .ZN(n617) );
  INV_X1 U691 ( .A(KEYINPUT2), .ZN(n615) );
  NOR2_X1 U692 ( .A1(n615), .A2(KEYINPUT67), .ZN(n616) );
  NAND2_X1 U693 ( .A1(n619), .A2(KEYINPUT2), .ZN(n620) );
  INV_X1 U694 ( .A(n621), .ZN(n622) );
  NAND2_X1 U695 ( .A1(n736), .A2(G472), .ZN(n626) );
  XOR2_X1 U696 ( .A(KEYINPUT62), .B(n624), .Z(n625) );
  XNOR2_X1 U697 ( .A(n626), .B(n625), .ZN(n629) );
  INV_X1 U698 ( .A(G952), .ZN(n627) );
  NAND2_X1 U699 ( .A1(n628), .A2(n627), .ZN(n654) );
  INV_X1 U700 ( .A(n654), .ZN(n739) );
  XNOR2_X1 U701 ( .A(n631), .B(n630), .ZN(G57) );
  XNOR2_X1 U702 ( .A(n632), .B(G140), .ZN(G42) );
  XNOR2_X1 U703 ( .A(n633), .B(G119), .ZN(G21) );
  XNOR2_X1 U704 ( .A(n634), .B(G101), .ZN(G3) );
  XOR2_X1 U705 ( .A(n605), .B(G122), .Z(G24) );
  XOR2_X1 U706 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n635) );
  XNOR2_X1 U707 ( .A(n636), .B(n635), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n642) );
  XOR2_X1 U710 ( .A(n642), .B(n622), .Z(n641) );
  NAND2_X1 U711 ( .A1(n641), .A2(n357), .ZN(n647) );
  XNOR2_X1 U712 ( .A(G227), .B(n642), .ZN(n643) );
  NAND2_X1 U713 ( .A1(n643), .A2(G900), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n644), .A2(G953), .ZN(n645) );
  XOR2_X1 U715 ( .A(KEYINPUT127), .B(n645), .Z(n646) );
  NAND2_X1 U716 ( .A1(n647), .A2(n646), .ZN(G72) );
  NAND2_X1 U717 ( .A1(n736), .A2(G478), .ZN(n648) );
  XOR2_X1 U718 ( .A(n649), .B(n648), .Z(n650) );
  NOR2_X1 U719 ( .A1(n650), .A2(n739), .ZN(G63) );
  NAND2_X1 U720 ( .A1(n736), .A2(G475), .ZN(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT59), .B(n651), .Z(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n655) );
  NAND2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n657) );
  XOR2_X1 U724 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n656) );
  XNOR2_X1 U725 ( .A(n657), .B(n656), .ZN(G60) );
  NAND2_X1 U726 ( .A1(n736), .A2(G469), .ZN(n662) );
  XNOR2_X1 U727 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n658) );
  XNOR2_X1 U728 ( .A(n658), .B(KEYINPUT57), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n662), .B(n661), .ZN(n663) );
  NOR2_X1 U731 ( .A1(n663), .A2(n739), .ZN(G54) );
  NOR2_X1 U732 ( .A1(n679), .A2(n665), .ZN(n664) );
  XOR2_X1 U733 ( .A(G104), .B(n664), .Z(G6) );
  NOR2_X1 U734 ( .A1(n682), .A2(n665), .ZN(n667) );
  XNOR2_X1 U735 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n666) );
  XNOR2_X1 U736 ( .A(n667), .B(n666), .ZN(n668) );
  XNOR2_X1 U737 ( .A(G107), .B(n668), .ZN(G9) );
  XOR2_X1 U738 ( .A(G110), .B(n669), .Z(G12) );
  XOR2_X1 U739 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n672) );
  NAND2_X1 U740 ( .A1(n677), .A2(n670), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n672), .B(n671), .ZN(n673) );
  XNOR2_X1 U742 ( .A(G128), .B(n673), .ZN(G30) );
  XOR2_X1 U743 ( .A(G143), .B(KEYINPUT117), .Z(n674) );
  XNOR2_X1 U744 ( .A(n675), .B(n674), .ZN(G45) );
  NAND2_X1 U745 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(n678), .B(G146), .ZN(G48) );
  NOR2_X1 U747 ( .A1(n679), .A2(n681), .ZN(n680) );
  XOR2_X1 U748 ( .A(G113), .B(n680), .Z(G15) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n683) );
  XOR2_X1 U750 ( .A(G116), .B(n683), .Z(G18) );
  NOR2_X1 U751 ( .A1(n622), .A2(KEYINPUT2), .ZN(n684) );
  NOR2_X1 U752 ( .A1(n685), .A2(n684), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n375), .A2(KEYINPUT2), .ZN(n687) );
  XNOR2_X1 U754 ( .A(n687), .B(KEYINPUT85), .ZN(n688) );
  AND2_X1 U755 ( .A1(n689), .A2(n688), .ZN(n726) );
  NOR2_X1 U756 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n698) );
  NOR2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U759 ( .A(n696), .B(KEYINPUT120), .ZN(n697) );
  NOR2_X1 U760 ( .A1(n698), .A2(n697), .ZN(n699) );
  XOR2_X1 U761 ( .A(KEYINPUT121), .B(n699), .Z(n700) );
  XOR2_X1 U762 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n704) );
  NOR2_X1 U763 ( .A1(n355), .A2(n701), .ZN(n703) );
  XOR2_X1 U764 ( .A(n704), .B(n703), .Z(n711) );
  NAND2_X1 U765 ( .A1(n556), .A2(n705), .ZN(n706) );
  XNOR2_X1 U766 ( .A(KEYINPUT49), .B(n706), .ZN(n707) );
  NOR2_X1 U767 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U768 ( .A(n709), .B(KEYINPUT118), .ZN(n710) );
  NAND2_X1 U769 ( .A1(n711), .A2(n710), .ZN(n713) );
  NAND2_X1 U770 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U771 ( .A(KEYINPUT51), .B(n714), .ZN(n715) );
  NOR2_X1 U772 ( .A1(n722), .A2(n715), .ZN(n716) );
  NOR2_X1 U773 ( .A1(n367), .A2(n716), .ZN(n717) );
  XNOR2_X1 U774 ( .A(KEYINPUT52), .B(n717), .ZN(n720) );
  NAND2_X1 U775 ( .A1(G952), .A2(n718), .ZN(n719) );
  NOR2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U777 ( .A1(G953), .A2(n721), .ZN(n724) );
  NAND2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U779 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U780 ( .A(KEYINPUT53), .B(n727), .ZN(G75) );
  NAND2_X1 U781 ( .A1(n736), .A2(G210), .ZN(n733) );
  XOR2_X1 U782 ( .A(KEYINPUT55), .B(KEYINPUT83), .Z(n729) );
  XNOR2_X1 U783 ( .A(KEYINPUT54), .B(KEYINPUT122), .ZN(n728) );
  XNOR2_X1 U784 ( .A(n729), .B(n728), .ZN(n731) );
  XOR2_X1 U785 ( .A(n731), .B(n358), .Z(n732) );
  XNOR2_X1 U786 ( .A(n733), .B(n732), .ZN(n734) );
  XNOR2_X1 U787 ( .A(n735), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U788 ( .A1(n736), .A2(G217), .ZN(n737) );
  XNOR2_X1 U789 ( .A(n738), .B(n737), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n375), .A2(n742), .ZN(n746) );
  NAND2_X1 U791 ( .A1(G953), .A2(G224), .ZN(n743) );
  XNOR2_X1 U792 ( .A(KEYINPUT61), .B(n743), .ZN(n744) );
  NAND2_X1 U793 ( .A1(n744), .A2(G898), .ZN(n745) );
  NAND2_X1 U794 ( .A1(n746), .A2(n745), .ZN(n753) );
  XOR2_X1 U795 ( .A(G101), .B(n747), .Z(n748) );
  XNOR2_X1 U796 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X1 U797 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U798 ( .A(n753), .B(n752), .ZN(G69) );
  XNOR2_X1 U799 ( .A(G134), .B(n754), .ZN(G36) );
  XOR2_X1 U800 ( .A(G125), .B(n755), .Z(n756) );
  XNOR2_X1 U801 ( .A(KEYINPUT37), .B(n756), .ZN(G27) );
  XOR2_X1 U802 ( .A(G137), .B(n757), .Z(G39) );
  XOR2_X1 U803 ( .A(n758), .B(G131), .Z(G33) );
endmodule

