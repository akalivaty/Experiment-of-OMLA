//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 1 1 1 1 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:39 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n529, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n558, new_n559,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n610, new_n611, new_n612, new_n615, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1241, new_n1242;
  XNOR2_X1  g000(.A(KEYINPUT64), .B(G452), .ZN(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XOR2_X1   g013(.A(KEYINPUT66), .B(G120), .Z(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  NAND2_X1  g032(.A1(new_n455), .A2(G567), .ZN(new_n458));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OAI21_X1  g034(.A(new_n458), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  OR2_X1    g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n472), .A2(G2104), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n471), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n468), .A2(new_n474), .ZN(G160));
  OR2_X1    g050(.A1(G100), .A2(G2105), .ZN(new_n476));
  OAI211_X1 g051(.A(new_n476), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n477));
  XNOR2_X1  g052(.A(KEYINPUT3), .B(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(G124), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n481), .B1(G136), .B2(new_n471), .ZN(G162));
  INV_X1    g057(.A(KEYINPUT4), .ZN(new_n483));
  INV_X1    g058(.A(KEYINPUT70), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(new_n472), .A3(G138), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n483), .B1(new_n465), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n487));
  INV_X1    g062(.A(G138), .ZN(new_n488));
  NOR3_X1   g063(.A1(new_n488), .A2(KEYINPUT70), .A3(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n478), .A2(KEYINPUT4), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT69), .B1(new_n472), .B2(G114), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  INV_X1    g067(.A(G114), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n492), .A2(new_n493), .A3(G2105), .ZN(new_n494));
  OR2_X1    g069(.A1(G102), .A2(G2105), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n491), .A2(new_n494), .A3(G2104), .A4(new_n495), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n486), .A2(new_n487), .A3(new_n490), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT71), .ZN(new_n499));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n499), .B1(new_n500), .B2(KEYINPUT72), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT71), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT6), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(new_n499), .B(KEYINPUT6), .C1(new_n500), .C2(KEYINPUT72), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n504), .A2(G543), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AOI22_X1  g088(.A1(new_n513), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n514), .A2(new_n500), .ZN(new_n515));
  AND3_X1   g090(.A1(new_n504), .A2(new_n505), .A3(new_n513), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G88), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n508), .A2(new_n515), .A3(new_n517), .ZN(G303));
  INV_X1    g093(.A(G303), .ZN(G166));
  NAND2_X1  g094(.A1(new_n507), .A2(G51), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(G89), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  OR2_X1    g097(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n522), .A2(KEYINPUT7), .ZN(new_n524));
  AND2_X1   g099(.A1(G63), .A2(G651), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n523), .A2(new_n524), .B1(new_n513), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n520), .A2(new_n521), .A3(new_n526), .ZN(G286));
  INV_X1    g102(.A(G286), .ZN(G168));
  NAND4_X1  g103(.A1(new_n504), .A2(G52), .A3(G543), .A4(new_n505), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n504), .A2(G90), .A3(new_n505), .A4(new_n513), .ZN(new_n530));
  AOI21_X1  g105(.A(KEYINPUT73), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT73), .ZN(new_n533));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  AND2_X1   g109(.A1(KEYINPUT5), .A2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(G64), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n534), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n532), .A2(new_n533), .B1(G651), .B2(new_n539), .ZN(G171));
  NAND4_X1  g115(.A1(new_n504), .A2(G43), .A3(G543), .A4(new_n505), .ZN(new_n541));
  NAND4_X1  g116(.A1(new_n504), .A2(G81), .A3(new_n505), .A4(new_n513), .ZN(new_n542));
  AND2_X1   g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n541), .A2(new_n542), .A3(KEYINPUT75), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n513), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT74), .B1(new_n546), .B2(new_n500), .ZN(new_n547));
  NAND2_X1  g122(.A1(G68), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(G56), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n537), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n550), .A2(new_n551), .A3(G651), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n544), .A2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  NAND4_X1  g131(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND4_X1  g134(.A1(G319), .A2(G483), .A3(G661), .A4(new_n559), .ZN(G188));
  AND4_X1   g135(.A1(G91), .A2(new_n504), .A3(new_n505), .A4(new_n513), .ZN(new_n561));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  INV_X1    g137(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n563), .B1(new_n513), .B2(G65), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT76), .B1(new_n564), .B2(new_n500), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n562), .B1(new_n537), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT76), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n567), .A2(new_n568), .A3(G651), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n561), .B1(new_n565), .B2(new_n569), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n504), .A2(G53), .A3(G543), .A4(new_n505), .ZN(new_n571));
  XNOR2_X1  g146(.A(new_n571), .B(KEYINPUT9), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n570), .A2(new_n572), .ZN(G299));
  NAND2_X1  g148(.A1(new_n539), .A2(G651), .ZN(new_n574));
  INV_X1    g149(.A(new_n533), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n531), .ZN(G301));
  NAND2_X1  g151(.A1(new_n507), .A2(G49), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n516), .A2(G87), .ZN(new_n578));
  OAI21_X1  g153(.A(G651), .B1(new_n513), .B2(G74), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G288));
  INV_X1    g155(.A(G61), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n511), .B2(new_n512), .ZN(new_n582));
  NAND2_X1  g157(.A1(G73), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT77), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n504), .A2(G48), .A3(G543), .A4(new_n505), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT77), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n588), .B(G651), .C1(new_n582), .C2(new_n584), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n504), .A2(G86), .A3(new_n505), .A4(new_n513), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(G305));
  NAND2_X1  g166(.A1(new_n507), .A2(G47), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n516), .A2(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n513), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n592), .B(new_n593), .C1(new_n500), .C2(new_n594), .ZN(G290));
  NAND2_X1  g170(.A1(G301), .A2(G868), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n504), .A2(G92), .A3(new_n505), .A4(new_n513), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  INV_X1    g173(.A(G66), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n599), .B1(new_n511), .B2(new_n512), .ZN(new_n600));
  AND2_X1   g175(.A1(G79), .A2(G543), .ZN(new_n601));
  OAI21_X1  g176(.A(G651), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND4_X1  g177(.A1(new_n504), .A2(G54), .A3(G543), .A4(new_n505), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n602), .A2(new_n603), .A3(KEYINPUT78), .ZN(new_n604));
  AOI21_X1  g179(.A(KEYINPUT78), .B1(new_n602), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n598), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G284));
  OAI21_X1  g183(.A(new_n596), .B1(new_n607), .B2(G868), .ZN(G321));
  INV_X1    g184(.A(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(G286), .A2(new_n610), .ZN(new_n611));
  XOR2_X1   g186(.A(G299), .B(KEYINPUT79), .Z(new_n612));
  AOI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(G297));
  AOI21_X1  g188(.A(new_n611), .B1(new_n612), .B2(new_n610), .ZN(G280));
  INV_X1    g189(.A(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n607), .B1(new_n615), .B2(G860), .ZN(G148));
  NAND2_X1  g191(.A1(new_n554), .A2(new_n610), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n606), .A2(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n610), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n478), .A2(new_n473), .ZN(new_n621));
  XOR2_X1   g196(.A(KEYINPUT80), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n621), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n471), .A2(G135), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n472), .A2(G111), .ZN(new_n629));
  OAI21_X1  g204(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n630));
  INV_X1    g205(.A(G123), .ZN(new_n631));
  OAI221_X1 g206(.A(new_n628), .B1(new_n629), .B2(new_n630), .C1(new_n631), .C2(new_n479), .ZN(new_n632));
  INV_X1    g207(.A(G2096), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n626), .A2(new_n627), .A3(new_n634), .ZN(G156));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2427), .B(G2430), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  AND2_X1   g215(.A1(new_n640), .A2(KEYINPUT82), .ZN(new_n641));
  NOR2_X1   g216(.A1(new_n640), .A2(KEYINPUT82), .ZN(new_n642));
  OAI22_X1  g217(.A1(new_n641), .A2(new_n642), .B1(new_n637), .B2(new_n638), .ZN(new_n643));
  XNOR2_X1  g218(.A(G1341), .B(G1348), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2451), .B(G2454), .Z(new_n646));
  XNOR2_X1  g221(.A(G2443), .B(G2446), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n645), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT81), .B(KEYINPUT16), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n652), .A2(G14), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT83), .Z(G401));
  INV_X1    g230(.A(KEYINPUT18), .ZN(new_n656));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n659), .A2(KEYINPUT17), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n656), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(new_n625), .ZN(new_n663));
  XOR2_X1   g238(.A(G2072), .B(G2078), .Z(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n659), .B2(KEYINPUT18), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(new_n633), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n663), .B(new_n666), .ZN(G227));
  XOR2_X1   g242(.A(G1971), .B(G1976), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  AND2_X1   g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n670), .A2(new_n671), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n669), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  AOI21_X1  g251(.A(new_n676), .B1(new_n669), .B2(new_n675), .ZN(new_n677));
  NAND2_X1  g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  XOR2_X1   g255(.A(G1991), .B(G1996), .Z(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1981), .B(G1986), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n680), .A2(new_n681), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n680), .A2(new_n681), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n685), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(G229));
  INV_X1    g265(.A(G16), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT86), .ZN(new_n694));
  INV_X1    g269(.A(G1971), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR2_X1   g271(.A1(G16), .A2(G23), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT85), .Z(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G288), .B2(new_n691), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT33), .ZN(new_n700));
  INV_X1    g275(.A(G1976), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n691), .A2(G6), .ZN(new_n703));
  OAI21_X1  g278(.A(G61), .B1(new_n535), .B2(new_n536), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n500), .B1(new_n704), .B2(new_n583), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n587), .B1(new_n705), .B2(new_n588), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n589), .A2(new_n590), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n703), .B1(new_n708), .B2(new_n691), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n694), .A2(new_n695), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n696), .A2(new_n702), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT84), .B(KEYINPUT34), .Z(new_n714));
  OR2_X1    g289(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n714), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n471), .A2(G131), .ZN(new_n717));
  NOR2_X1   g292(.A1(new_n472), .A2(G107), .ZN(new_n718));
  OAI21_X1  g293(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n719));
  INV_X1    g294(.A(G119), .ZN(new_n720));
  OAI221_X1 g295(.A(new_n717), .B1(new_n718), .B2(new_n719), .C1(new_n720), .C2(new_n479), .ZN(new_n721));
  MUX2_X1   g296(.A(G25), .B(new_n721), .S(G29), .Z(new_n722));
  XOR2_X1   g297(.A(KEYINPUT35), .B(G1991), .Z(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(G1986), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n691), .A2(G24), .ZN(new_n726));
  AOI21_X1  g301(.A(new_n726), .B1(G290), .B2(G16), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n724), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n725), .B2(new_n727), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n715), .A2(new_n716), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT36), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n691), .A2(G21), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G168), .B2(new_n691), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n691), .A2(G19), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n735), .B1(new_n555), .B2(new_n691), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(G1341), .ZN(new_n737));
  NOR2_X1   g312(.A1(G29), .A2(G35), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n738), .B1(G162), .B2(G29), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT92), .B(KEYINPUT29), .Z(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  AOI211_X1 g317(.A(new_n734), .B(new_n737), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n691), .A2(G20), .ZN(new_n744));
  XOR2_X1   g319(.A(new_n744), .B(KEYINPUT23), .Z(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G299), .B2(G16), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(G1956), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n607), .A2(new_n691), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(G4), .B2(new_n691), .ZN(new_n749));
  XOR2_X1   g324(.A(KEYINPUT87), .B(G1348), .Z(new_n750));
  NAND2_X1  g325(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g326(.A1(new_n743), .A2(new_n747), .A3(new_n751), .ZN(new_n752));
  INV_X1    g327(.A(G1961), .ZN(new_n753));
  NOR2_X1   g328(.A1(G171), .A2(new_n691), .ZN(new_n754));
  AOI21_X1  g329(.A(new_n754), .B1(G5), .B2(new_n691), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n753), .A2(new_n755), .B1(new_n736), .B2(G1341), .ZN(new_n756));
  OAI221_X1 g331(.A(new_n756), .B1(new_n753), .B2(new_n755), .C1(new_n749), .C2(new_n750), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n741), .A2(new_n742), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT25), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n471), .A2(G139), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(G115), .A2(G2104), .ZN(new_n764));
  INV_X1    g339(.A(G127), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n764), .B1(new_n465), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(G2105), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT88), .ZN(new_n768));
  INV_X1    g343(.A(G29), .ZN(new_n769));
  NOR2_X1   g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(new_n769), .B2(G33), .ZN(new_n771));
  INV_X1    g346(.A(G2072), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n758), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n769), .A2(G32), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n473), .A2(G105), .ZN(new_n775));
  NAND3_X1  g350(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT26), .ZN(new_n777));
  INV_X1    g352(.A(new_n479), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n775), .B(new_n777), .C1(new_n778), .C2(G129), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n471), .A2(G141), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT90), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n774), .B1(new_n783), .B2(new_n769), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT27), .B(G1996), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OAI211_X1 g361(.A(new_n773), .B(new_n786), .C1(new_n772), .C2(new_n771), .ZN(new_n787));
  XNOR2_X1  g362(.A(KEYINPUT31), .B(G11), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(KEYINPUT91), .ZN(new_n789));
  INV_X1    g364(.A(KEYINPUT30), .ZN(new_n790));
  AND2_X1   g365(.A1(new_n790), .A2(G28), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n769), .B1(new_n790), .B2(G28), .ZN(new_n792));
  OAI221_X1 g367(.A(new_n789), .B1(new_n791), .B2(new_n792), .C1(new_n632), .C2(new_n769), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n471), .A2(G140), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n472), .A2(G116), .ZN(new_n795));
  OAI21_X1  g370(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n796));
  INV_X1    g371(.A(G128), .ZN(new_n797));
  OAI221_X1 g372(.A(new_n794), .B1(new_n795), .B2(new_n796), .C1(new_n797), .C2(new_n479), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n798), .A2(G29), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n769), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2067), .ZN(new_n803));
  INV_X1    g378(.A(G2078), .ZN(new_n804));
  NAND2_X1  g379(.A1(G164), .A2(G29), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G27), .B2(G29), .ZN(new_n806));
  AOI211_X1 g381(.A(new_n793), .B(new_n803), .C1(new_n804), .C2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n808));
  INV_X1    g383(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g384(.A(G29), .B1(new_n809), .B2(G34), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G34), .B2(new_n809), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(G160), .B2(new_n769), .ZN(new_n812));
  INV_X1    g387(.A(G2084), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n807), .B(new_n814), .C1(new_n804), .C2(new_n806), .ZN(new_n815));
  NOR4_X1   g390(.A1(new_n752), .A2(new_n757), .A3(new_n787), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n731), .A2(new_n816), .ZN(G150));
  INV_X1    g392(.A(G150), .ZN(G311));
  NOR2_X1   g393(.A1(new_n606), .A2(new_n615), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT94), .ZN(new_n820));
  XOR2_X1   g395(.A(new_n820), .B(KEYINPUT38), .Z(new_n821));
  OR2_X1    g396(.A1(new_n543), .A2(KEYINPUT75), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n504), .A2(G93), .A3(new_n505), .A4(new_n513), .ZN(new_n823));
  INV_X1    g398(.A(G55), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n823), .B1(new_n506), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g400(.A1(G80), .A2(G543), .ZN(new_n826));
  INV_X1    g401(.A(G67), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n537), .B2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n500), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  OAI211_X1 g405(.A(KEYINPUT93), .B(new_n826), .C1(new_n537), .C2(new_n827), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n825), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND2_X1   g407(.A1(new_n547), .A2(new_n552), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n822), .A2(new_n832), .A3(new_n545), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n831), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n507), .A2(G55), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n835), .A2(new_n836), .A3(new_n823), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n544), .B2(new_n553), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n834), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n821), .B(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT39), .ZN(new_n841));
  AOI21_X1  g416(.A(G860), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n837), .A2(G860), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT37), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(G145));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  XNOR2_X1  g422(.A(G160), .B(new_n632), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(G162), .Z(new_n849));
  XOR2_X1   g424(.A(new_n721), .B(new_n623), .Z(new_n850));
  NAND2_X1  g425(.A1(new_n778), .A2(G130), .ZN(new_n851));
  OAI21_X1  g426(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n852));
  INV_X1    g427(.A(G118), .ZN(new_n853));
  AOI22_X1  g428(.A1(new_n852), .A2(KEYINPUT95), .B1(new_n853), .B2(G2105), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n854), .B1(KEYINPUT95), .B2(new_n852), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n471), .A2(G142), .ZN(new_n856));
  AND3_X1   g431(.A1(new_n851), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n850), .B(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n767), .B(KEYINPUT88), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n798), .B(G164), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n768), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n783), .A3(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n783), .B1(new_n862), .B2(new_n864), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n859), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT96), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n862), .A2(new_n864), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n782), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n865), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT96), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n859), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n869), .A2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n866), .A2(new_n867), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n876), .A2(new_n858), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n849), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(G37), .ZN(new_n879));
  NAND4_X1  g454(.A1(new_n871), .A2(KEYINPUT97), .A3(new_n858), .A4(new_n865), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n868), .A2(new_n880), .A3(new_n849), .ZN(new_n881));
  AOI21_X1  g456(.A(KEYINPUT97), .B1(new_n876), .B2(new_n858), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n847), .B1(new_n878), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n883), .ZN(new_n885));
  AOI21_X1  g460(.A(new_n873), .B1(new_n872), .B2(new_n859), .ZN(new_n886));
  AOI211_X1 g461(.A(KEYINPUT96), .B(new_n858), .C1(new_n871), .C2(new_n865), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n877), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n849), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n885), .A2(new_n890), .A3(KEYINPUT98), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n884), .A2(new_n891), .A3(KEYINPUT40), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT40), .B1(new_n884), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G395));
  XOR2_X1   g469(.A(G303), .B(G288), .Z(new_n895));
  XNOR2_X1  g470(.A(G290), .B(G305), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n895), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n834), .A2(new_n838), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n898), .B1(new_n834), .B2(new_n838), .ZN(new_n901));
  OAI22_X1  g476(.A1(new_n900), .A2(new_n901), .B1(G559), .B2(new_n606), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n618), .A3(new_n899), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n606), .A2(G299), .ZN(new_n906));
  OR2_X1    g481(.A1(new_n604), .A2(new_n605), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n907), .A2(new_n572), .A3(new_n570), .A4(new_n598), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT41), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT41), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n906), .A2(new_n911), .A3(new_n908), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n905), .A2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT100), .ZN(new_n915));
  XNOR2_X1  g490(.A(new_n909), .B(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n916), .A2(new_n902), .A3(new_n904), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT42), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n914), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n897), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  INV_X1    g498(.A(new_n897), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n922), .A2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n926), .A2(G868), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n832), .A2(G868), .ZN(new_n928));
  INV_X1    g503(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(G295));
  INV_X1    g505(.A(KEYINPUT101), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n931), .A3(new_n929), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n610), .B1(new_n922), .B2(new_n925), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT101), .B1(new_n933), .B2(new_n928), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(G331));
  INV_X1    g510(.A(KEYINPUT102), .ZN(new_n936));
  NOR2_X1   g511(.A1(G171), .A2(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(G286), .B1(G171), .B2(new_n936), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n839), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g514(.A(G168), .B1(G301), .B2(KEYINPUT102), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n940), .A2(new_n838), .A3(new_n834), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n939), .A2(new_n937), .A3(new_n941), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n943), .A2(new_n944), .B1(new_n912), .B2(new_n910), .ZN(new_n945));
  AND3_X1   g520(.A1(new_n939), .A2(new_n937), .A3(new_n941), .ZN(new_n946));
  NOR3_X1   g521(.A1(new_n946), .A2(new_n942), .A3(new_n909), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n897), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(new_n906), .A3(new_n908), .A4(new_n944), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n913), .B1(new_n946), .B2(new_n942), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(new_n924), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n948), .A2(new_n879), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n946), .A2(new_n942), .ZN(new_n955));
  INV_X1    g530(.A(new_n916), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n912), .B(KEYINPUT104), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT105), .B1(new_n909), .B2(KEYINPUT41), .ZN(new_n959));
  AND3_X1   g534(.A1(new_n909), .A2(KEYINPUT105), .A3(KEYINPUT41), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n958), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n957), .B(new_n897), .C1(new_n961), .C2(new_n955), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n962), .A2(new_n879), .A3(new_n951), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n954), .B1(new_n953), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(KEYINPUT44), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT103), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n951), .A2(new_n879), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n924), .B1(new_n949), .B2(new_n950), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n966), .B(KEYINPUT43), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n952), .B2(KEYINPUT43), .ZN(new_n971));
  AND4_X1   g546(.A1(new_n953), .A2(new_n962), .A3(new_n879), .A4(new_n951), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n970), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n965), .B1(new_n973), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT63), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT109), .ZN(new_n976));
  NOR3_X1   g551(.A1(new_n465), .A2(new_n483), .A3(new_n485), .ZN(new_n977));
  AOI21_X1  g552(.A(KEYINPUT4), .B1(new_n478), .B2(new_n489), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n496), .A2(new_n487), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT50), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n976), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n497), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n985), .A2(KEYINPUT109), .A3(KEYINPUT50), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n983), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(KEYINPUT108), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT108), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n497), .A2(new_n990), .A3(new_n984), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n982), .A3(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n987), .A2(new_n742), .A3(new_n988), .A4(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n468), .A2(G40), .A3(new_n474), .ZN(new_n994));
  XOR2_X1   g569(.A(KEYINPUT106), .B(KEYINPUT45), .Z(new_n995));
  AOI21_X1  g570(.A(new_n994), .B1(new_n985), .B2(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n984), .ZN(new_n997));
  AOI21_X1  g572(.A(G1971), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n993), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(G303), .A2(G8), .ZN(new_n1001));
  XNOR2_X1  g576(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1002));
  INV_X1    g577(.A(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(G303), .A2(G8), .A3(new_n1002), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1000), .A2(G8), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n988), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n989), .A2(new_n991), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(KEYINPUT50), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n998), .B1(new_n1011), .B2(new_n742), .ZN(new_n1012));
  INV_X1    g587(.A(G8), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n585), .A2(new_n587), .A3(new_n590), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(G1981), .ZN(new_n1016));
  INV_X1    g591(.A(G1981), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT111), .B1(new_n708), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n1019));
  NOR4_X1   g594(.A1(new_n706), .A2(new_n707), .A3(new_n1019), .A4(G1981), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n497), .A2(new_n990), .A3(new_n984), .ZN(new_n1024));
  AOI21_X1  g599(.A(new_n990), .B1(new_n497), .B2(new_n984), .ZN(new_n1025));
  NOR2_X1   g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1013), .B1(new_n1026), .B2(new_n988), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1019), .B1(G305), .B2(G1981), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n708), .A2(KEYINPUT111), .A3(new_n1017), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1030), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1023), .A2(new_n1027), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n989), .A2(new_n988), .A3(new_n991), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n577), .A2(new_n578), .A3(G1976), .A4(new_n579), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(G8), .A3(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1035), .A2(KEYINPUT52), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT52), .B1(G288), .B2(new_n701), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1033), .A2(new_n1037), .A3(G8), .A4(new_n1034), .ZN(new_n1038));
  AND2_X1   g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1008), .A2(new_n1014), .A3(new_n1032), .A4(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G286), .A2(new_n1013), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n987), .A2(new_n813), .A3(new_n988), .A4(new_n992), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT45), .B1(new_n989), .B2(new_n991), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n988), .B1(new_n985), .B2(new_n995), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1044), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1042), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n975), .B1(new_n1040), .B2(new_n1049), .ZN(new_n1050));
  AOI211_X1 g625(.A(new_n1013), .B(new_n1006), .C1(new_n993), .C2(new_n999), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1052), .A2(KEYINPUT63), .A3(new_n1041), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1039), .A2(new_n1032), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1013), .B1(new_n993), .B2(new_n999), .ZN(new_n1057));
  OR2_X1    g632(.A1(new_n1057), .A2(new_n1007), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1054), .A2(new_n1055), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1008), .A2(KEYINPUT63), .A3(new_n1048), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1039), .B(new_n1032), .C1(new_n1057), .C2(new_n1007), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT113), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1050), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(G288), .A2(G1976), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n1023), .B2(new_n1031), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1030), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1027), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1039), .A2(new_n1032), .A3(new_n1057), .A4(new_n1007), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1069), .A2(KEYINPUT112), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT112), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1067), .A2(new_n1068), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1070), .A2(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1063), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT114), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT50), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n994), .B1(new_n981), .B2(new_n982), .ZN(new_n1078));
  AOI21_X1  g653(.A(G1956), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(KEYINPUT56), .B(G2072), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n996), .A2(new_n997), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT57), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT9), .ZN(new_n1084));
  XNOR2_X1  g659(.A(new_n571), .B(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n1086));
  OAI21_X1  g661(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT116), .ZN(new_n1088));
  AND3_X1   g663(.A1(new_n570), .A2(new_n572), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1088), .B1(new_n570), .B2(new_n572), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1087), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n565), .A2(new_n569), .ZN(new_n1092));
  INV_X1    g667(.A(new_n561), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(KEYINPUT116), .B1(new_n1094), .B2(new_n1085), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT57), .B1(new_n572), .B2(KEYINPUT115), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n570), .A2(new_n572), .A3(new_n1088), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1096), .A3(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1091), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1082), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1082), .A2(new_n1099), .A3(KEYINPUT117), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1091), .B(new_n1098), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n992), .A2(new_n988), .ZN(new_n1106));
  AOI21_X1  g681(.A(KEYINPUT109), .B1(new_n985), .B2(KEYINPUT50), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n976), .B(new_n982), .C1(new_n497), .C2(new_n984), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n750), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1033), .A2(G2067), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n606), .B1(new_n1110), .B2(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1105), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n994), .B1(new_n1026), .B2(new_n982), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n987), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1111), .B1(new_n1117), .B2(new_n750), .ZN(new_n1118));
  NOR3_X1   g693(.A1(new_n1118), .A2(KEYINPUT118), .A3(new_n606), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1104), .B1(new_n1115), .B2(new_n1119), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n996), .A2(new_n997), .ZN(new_n1122));
  XOR2_X1   g697(.A(KEYINPUT119), .B(G1996), .Z(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT58), .B(G1341), .Z(new_n1125));
  NAND2_X1  g700(.A1(new_n1033), .A2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1125), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1124), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n555), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AND3_X1   g707(.A1(new_n1033), .A2(KEYINPUT120), .A3(new_n1125), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT120), .B1(new_n1033), .B2(new_n1125), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1133), .A2(new_n1134), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1135), .A2(KEYINPUT121), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1121), .B1(new_n1132), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT60), .ZN(new_n1138));
  NAND3_X1  g713(.A1(new_n1118), .A2(new_n1138), .A3(new_n607), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1110), .A2(new_n606), .A3(new_n1112), .ZN(new_n1140));
  OAI21_X1  g715(.A(KEYINPUT60), .B1(new_n1140), .B2(new_n1113), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1137), .A2(new_n1139), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n554), .B1(new_n1135), .B2(KEYINPUT121), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT59), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1145), .A2(KEYINPUT122), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1143), .A2(new_n1144), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT123), .ZN(new_n1148));
  AND4_X1   g723(.A1(new_n1148), .A2(new_n1100), .A3(KEYINPUT61), .A4(new_n1105), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1150), .B1(new_n1082), .B2(new_n1099), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1151), .B2(new_n1105), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1147), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1120), .B1(new_n1142), .B2(new_n1153), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n753), .B1(new_n1106), .B2(new_n1109), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT125), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI211_X1 g732(.A(KEYINPUT125), .B(new_n753), .C1(new_n1106), .C2(new_n1109), .ZN(new_n1158));
  INV_X1    g733(.A(new_n1122), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n804), .A2(KEYINPUT53), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n996), .A2(new_n804), .A3(new_n997), .ZN(new_n1161));
  XNOR2_X1  g736(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1159), .A2(new_n1160), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1157), .A2(G301), .A3(new_n1158), .A4(new_n1163), .ZN(new_n1164));
  AOI21_X1  g739(.A(G1961), .B1(new_n1116), .B2(new_n987), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT45), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1166), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n985), .A2(new_n995), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n988), .A3(new_n1160), .A4(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  OAI21_X1  g746(.A(G171), .B1(new_n1165), .B2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(KEYINPUT54), .B1(new_n1164), .B2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT126), .ZN(new_n1174));
  XNOR2_X1  g749(.A(new_n1173), .B(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1043), .A2(G168), .A3(new_n1047), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1176), .A2(G8), .ZN(new_n1177));
  AOI21_X1  g752(.A(G168), .B1(new_n1043), .B2(new_n1047), .ZN(new_n1178));
  OAI21_X1  g753(.A(KEYINPUT51), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT51), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1176), .A2(new_n1180), .A3(G8), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1179), .A2(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1157), .A2(new_n1158), .A3(new_n1163), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1183), .A2(G171), .ZN(new_n1184));
  INV_X1    g759(.A(KEYINPUT54), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1165), .A2(new_n1171), .ZN(new_n1186));
  AOI21_X1  g761(.A(new_n1185), .B1(new_n1186), .B2(G301), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g763(.A(new_n1040), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1102), .A2(new_n1150), .A3(new_n1103), .ZN(new_n1190));
  AND4_X1   g765(.A1(new_n1182), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND3_X1  g766(.A1(new_n1154), .A2(new_n1175), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g767(.A(KEYINPUT127), .ZN(new_n1193));
  INV_X1    g768(.A(new_n1181), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1178), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1195), .A2(G8), .A3(new_n1176), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1194), .B1(new_n1196), .B2(KEYINPUT51), .ZN(new_n1197));
  INV_X1    g772(.A(KEYINPUT62), .ZN(new_n1198));
  OAI21_X1  g773(.A(new_n1193), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1182), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n1040), .A2(new_n1172), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1063), .A2(new_n1073), .A3(KEYINPUT114), .ZN(new_n1204));
  NAND4_X1  g779(.A1(new_n1076), .A2(new_n1192), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n985), .A2(new_n995), .ZN(new_n1206));
  NOR2_X1   g781(.A1(new_n1206), .A2(new_n994), .ZN(new_n1207));
  XNOR2_X1  g782(.A(new_n798), .B(G2067), .ZN(new_n1208));
  XNOR2_X1  g783(.A(new_n1208), .B(KEYINPUT107), .ZN(new_n1209));
  INV_X1    g784(.A(G1996), .ZN(new_n1210));
  XNOR2_X1  g785(.A(new_n782), .B(new_n1210), .ZN(new_n1211));
  INV_X1    g786(.A(new_n723), .ZN(new_n1212));
  OR2_X1    g787(.A1(new_n721), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n721), .A2(new_n1212), .ZN(new_n1214));
  AND4_X1   g789(.A1(new_n1209), .A2(new_n1211), .A3(new_n1213), .A4(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g791(.A(G290), .B(G1986), .ZN(new_n1217));
  OAI21_X1  g792(.A(new_n1207), .B1(new_n1216), .B2(new_n1217), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1205), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g794(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1220));
  XOR2_X1   g795(.A(new_n1220), .B(KEYINPUT46), .Z(new_n1221));
  NAND2_X1  g796(.A1(new_n1209), .A2(new_n783), .ZN(new_n1222));
  AOI21_X1  g797(.A(new_n1221), .B1(new_n1222), .B2(new_n1207), .ZN(new_n1223));
  XOR2_X1   g798(.A(new_n1223), .B(KEYINPUT47), .Z(new_n1224));
  NAND2_X1  g799(.A1(new_n1216), .A2(new_n1207), .ZN(new_n1225));
  NOR2_X1   g800(.A1(G290), .A2(G1986), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1226), .A2(new_n1207), .ZN(new_n1227));
  XNOR2_X1  g802(.A(new_n1227), .B(KEYINPUT48), .ZN(new_n1228));
  NAND2_X1  g803(.A1(new_n1209), .A2(new_n1211), .ZN(new_n1229));
  OAI22_X1  g804(.A1(new_n1229), .A2(new_n1213), .B1(G2067), .B2(new_n798), .ZN(new_n1230));
  AOI22_X1  g805(.A1(new_n1225), .A2(new_n1228), .B1(new_n1207), .B2(new_n1230), .ZN(new_n1231));
  AND2_X1   g806(.A1(new_n1224), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g807(.A1(new_n1219), .A2(new_n1232), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g808(.A1(G227), .A2(new_n460), .ZN(new_n1235));
  AND3_X1   g809(.A1(new_n654), .A2(new_n689), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g810(.A(KEYINPUT98), .B1(new_n885), .B2(new_n890), .ZN(new_n1237));
  NOR3_X1   g811(.A1(new_n878), .A2(new_n847), .A3(new_n883), .ZN(new_n1238));
  OAI21_X1  g812(.A(new_n1236), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1239), .A2(new_n973), .ZN(G308));
  NAND2_X1  g814(.A1(new_n884), .A2(new_n891), .ZN(new_n1241));
  OR2_X1    g815(.A1(new_n971), .A2(new_n972), .ZN(new_n1242));
  OAI211_X1 g816(.A(new_n1241), .B(new_n1236), .C1(new_n1242), .C2(new_n970), .ZN(G225));
endmodule


