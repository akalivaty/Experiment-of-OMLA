//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0 1 0 1 1 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:03 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G952), .ZN(new_n189));
  NAND2_X1  g003(.A1(G234), .A2(G237), .ZN(new_n190));
  AND2_X1   g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  AND3_X1   g006(.A1(new_n190), .A2(G902), .A3(G953), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT21), .B(G898), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT2), .B(G113), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  OR2_X1    g012(.A1(KEYINPUT68), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(KEYINPUT68), .A2(G119), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(G116), .A3(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G116), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G119), .ZN(new_n203));
  AND2_X1   g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT67), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n198), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n201), .A2(new_n203), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT67), .A3(new_n197), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT4), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT78), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G104), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n211), .A2(KEYINPUT3), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n213), .A2(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT3), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n213), .A3(KEYINPUT78), .A4(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n210), .B(G101), .C1(new_n217), .C2(new_n221), .ZN(new_n222));
  OAI21_X1  g036(.A(G101), .B1(new_n217), .B2(new_n221), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n219), .A2(KEYINPUT78), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n219), .A2(KEYINPUT78), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(new_n214), .ZN(new_n226));
  INV_X1    g040(.A(G101), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n226), .A2(new_n227), .A3(new_n218), .A4(new_n220), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n209), .A2(new_n222), .A3(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(G110), .B(G122), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT84), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n201), .A2(KEYINPUT5), .A3(new_n203), .ZN(new_n233));
  INV_X1    g047(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(G113), .B1(new_n201), .B2(KEYINPUT5), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n232), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OR2_X1    g050(.A1(new_n201), .A2(KEYINPUT5), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n237), .A2(KEYINPUT84), .A3(G113), .A4(new_n233), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n204), .A2(new_n198), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n236), .A2(new_n238), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT79), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n218), .A2(new_n214), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n228), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n241), .B1(new_n228), .B2(new_n243), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n230), .B(new_n231), .C1(new_n240), .C2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G143), .ZN(new_n248));
  OAI21_X1  g062(.A(KEYINPUT1), .B1(new_n248), .B2(G146), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G128), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(KEYINPUT65), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G143), .ZN(new_n253));
  AOI21_X1  g067(.A(G146), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(G146), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n255), .A2(G143), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n250), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n251), .A2(new_n253), .A3(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT66), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n248), .B2(G146), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n255), .A2(KEYINPUT66), .A3(G143), .ZN(new_n261));
  INV_X1    g075(.A(G128), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT1), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n257), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G125), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT0), .A2(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n271), .B1(new_n254), .B2(new_n256), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n269), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(G125), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT86), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT7), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n268), .A2(new_n275), .A3(new_n277), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT85), .B(G224), .Z(new_n279));
  OAI21_X1  g093(.A(KEYINPUT7), .B1(new_n279), .B2(G953), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(new_n280), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n268), .A2(new_n275), .A3(new_n282), .A4(new_n277), .ZN(new_n283));
  AND3_X1   g097(.A1(new_n247), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n228), .A2(new_n243), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n240), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n239), .B1(new_n234), .B2(new_n235), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n286), .B1(new_n246), .B2(new_n287), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n231), .B(KEYINPUT8), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n284), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n230), .B1(new_n240), .B2(new_n246), .ZN(new_n292));
  INV_X1    g106(.A(new_n231), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(KEYINPUT6), .A3(new_n247), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n296), .A3(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n268), .A2(new_n275), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n279), .A2(G953), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n295), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n291), .A2(new_n301), .A3(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n302), .B1(new_n291), .B2(new_n301), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n187), .B(new_n196), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G475), .ZN(new_n306));
  INV_X1    g120(.A(G902), .ZN(new_n307));
  INV_X1    g121(.A(G237), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(new_n188), .A3(G214), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n251), .A2(new_n253), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n309), .B1(new_n310), .B2(KEYINPUT87), .ZN(new_n311));
  AOI21_X1  g125(.A(G143), .B1(new_n252), .B2(KEYINPUT87), .ZN(new_n312));
  NAND4_X1  g126(.A1(new_n312), .A2(G214), .A3(new_n308), .A4(new_n188), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G131), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT17), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n311), .A2(G131), .A3(new_n313), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(new_n321), .A3(G125), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(G125), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n267), .A2(G140), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n322), .B1(new_n325), .B2(new_n320), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(new_n255), .ZN(new_n327));
  XNOR2_X1  g141(.A(G125), .B(G140), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(KEYINPUT16), .ZN(new_n329));
  AOI21_X1  g143(.A(G146), .B1(new_n329), .B2(new_n322), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT17), .A4(G131), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n319), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n328), .B(G146), .ZN(new_n334));
  NAND2_X1  g148(.A1(KEYINPUT18), .A2(G131), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n314), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT18), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(new_n318), .ZN(new_n338));
  XNOR2_X1  g152(.A(G113), .B(G122), .ZN(new_n339));
  OR2_X1    g153(.A1(new_n339), .A2(KEYINPUT90), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(KEYINPUT90), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT89), .B(G104), .ZN(new_n343));
  XNOR2_X1  g157(.A(new_n342), .B(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n333), .A2(new_n338), .A3(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n344), .B1(new_n333), .B2(new_n338), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n307), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n306), .B1(new_n347), .B2(KEYINPUT91), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT91), .ZN(new_n349));
  OAI211_X1 g163(.A(new_n349), .B(new_n307), .C1(new_n345), .C2(new_n346), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(G475), .A2(G902), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT88), .ZN(new_n353));
  INV_X1    g167(.A(new_n318), .ZN(new_n354));
  AOI21_X1  g168(.A(G131), .B1(new_n311), .B2(new_n313), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n353), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n316), .A2(KEYINPUT88), .A3(new_n318), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n328), .B(KEYINPUT19), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n327), .B1(new_n255), .B2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n344), .B1(new_n360), .B2(new_n338), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n352), .B1(new_n345), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(KEYINPUT20), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT20), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n364), .B(new_n352), .C1(new_n345), .C2(new_n361), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n351), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G478), .ZN(new_n368));
  NOR2_X1   g182(.A1(new_n368), .A2(KEYINPUT15), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT92), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n310), .A2(new_n262), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(KEYINPUT13), .ZN(new_n372));
  XNOR2_X1  g186(.A(KEYINPUT65), .B(G143), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G128), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT13), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(KEYINPUT92), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n262), .A2(G143), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n371), .A2(KEYINPUT13), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n372), .A2(new_n376), .A3(new_n377), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G134), .ZN(new_n380));
  INV_X1    g194(.A(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G116), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n202), .A2(G122), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n384), .B(G107), .ZN(new_n385));
  INV_X1    g199(.A(G134), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n374), .A2(new_n386), .A3(new_n377), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n380), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n213), .B1(new_n382), .B2(KEYINPUT14), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n391), .A2(new_n384), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n384), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n374), .A2(new_n377), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G134), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n394), .B1(new_n387), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  XNOR2_X1  g212(.A(KEYINPUT9), .B(G234), .ZN(new_n399));
  INV_X1    g213(.A(G217), .ZN(new_n400));
  NOR3_X1   g214(.A1(new_n399), .A2(new_n400), .A3(G953), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(new_n401), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n388), .B1(new_n379), .B2(G134), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n403), .B1(new_n404), .B2(new_n397), .ZN(new_n405));
  AOI21_X1  g219(.A(G902), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT93), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI211_X1 g222(.A(KEYINPUT93), .B(G902), .C1(new_n402), .C2(new_n405), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n369), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  OAI22_X1  g224(.A1(new_n406), .A2(new_n407), .B1(KEYINPUT15), .B2(new_n368), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n305), .A2(new_n367), .A3(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G221), .B1(new_n399), .B2(G902), .ZN(new_n414));
  XOR2_X1   g228(.A(new_n414), .B(KEYINPUT77), .Z(new_n415));
  INV_X1    g229(.A(G469), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT10), .ZN(new_n417));
  AND4_X1   g231(.A1(new_n258), .A2(new_n260), .A3(new_n261), .A4(new_n263), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n258), .A2(new_n260), .A3(new_n261), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT1), .ZN(new_n420));
  OAI21_X1  g234(.A(G128), .B1(new_n254), .B2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(new_n418), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n417), .B1(new_n422), .B2(new_n285), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n417), .B1(new_n257), .B2(new_n264), .ZN(new_n424));
  OAI21_X1  g238(.A(new_n424), .B1(new_n244), .B2(new_n245), .ZN(new_n425));
  AND2_X1   g239(.A1(new_n272), .A2(new_n273), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n229), .A2(new_n426), .A3(new_n222), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n423), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT11), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n429), .B1(new_n386), .B2(G137), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n386), .A2(G137), .ZN(new_n431));
  INV_X1    g245(.A(G137), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n432), .A2(KEYINPUT11), .A3(G134), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n431), .A3(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(G131), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n430), .A2(new_n433), .A3(new_n315), .A4(new_n431), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n437), .B(KEYINPUT80), .Z(new_n438));
  OR2_X1    g252(.A1(new_n428), .A2(new_n438), .ZN(new_n439));
  AND3_X1   g253(.A1(new_n428), .A2(KEYINPUT82), .A3(new_n437), .ZN(new_n440));
  AOI21_X1  g254(.A(KEYINPUT82), .B1(new_n428), .B2(new_n437), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n439), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G110), .B(G140), .ZN(new_n443));
  AND2_X1   g257(.A1(new_n188), .A2(G227), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n442), .A2(KEYINPUT83), .A3(new_n445), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n428), .A2(new_n438), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(new_n445), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n246), .A2(new_n266), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n449), .B1(new_n285), .B2(new_n422), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT12), .ZN(new_n451));
  NAND4_X1  g265(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n451), .A4(new_n437), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(KEYINPUT81), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n422), .A2(new_n285), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n246), .B2(new_n266), .ZN(new_n456));
  INV_X1    g270(.A(new_n437), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n453), .B(new_n454), .C1(new_n456), .C2(new_n457), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n448), .A2(new_n452), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n446), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT83), .B1(new_n442), .B2(new_n445), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n416), .B(new_n307), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n416), .A2(new_n307), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n452), .A2(new_n458), .A3(new_n439), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n428), .A2(new_n437), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT82), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n428), .A2(KEYINPUT82), .A3(new_n437), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n464), .A2(new_n445), .B1(new_n469), .B2(new_n448), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n463), .B1(new_n470), .B2(G469), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n415), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n413), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT94), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n400), .B1(G234), .B2(new_n307), .ZN(new_n476));
  XNOR2_X1  g290(.A(KEYINPUT22), .B(G137), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT24), .B(G110), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n199), .A2(G128), .A3(new_n200), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n262), .A2(G119), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n485), .B1(new_n327), .B2(new_n330), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n262), .A2(KEYINPUT23), .A3(G119), .ZN(new_n487));
  XOR2_X1   g301(.A(new_n487), .B(KEYINPUT72), .Z(new_n488));
  NAND2_X1  g302(.A1(new_n483), .A2(KEYINPUT23), .ZN(new_n489));
  INV_X1    g303(.A(new_n200), .ZN(new_n490));
  NOR2_X1   g304(.A1(KEYINPUT68), .A2(G119), .ZN(new_n491));
  OAI211_X1 g305(.A(KEYINPUT73), .B(new_n262), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(G128), .B1(new_n199), .B2(new_n200), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n488), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n486), .B1(G110), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n329), .A2(G146), .A3(new_n322), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(G146), .B2(new_n325), .ZN(new_n499));
  INV_X1    g313(.A(G110), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n500), .B(new_n488), .C1(new_n493), .C2(new_n495), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n483), .A2(new_n484), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n502), .A2(new_n481), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT74), .ZN(new_n505));
  NOR3_X1   g319(.A1(new_n497), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n501), .A2(new_n503), .ZN(new_n507));
  INV_X1    g321(.A(new_n499), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n496), .A2(G110), .ZN(new_n510));
  INV_X1    g324(.A(new_n485), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n326), .A2(new_n255), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n511), .B1(new_n512), .B2(new_n498), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(KEYINPUT74), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n480), .B1(new_n506), .B2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n480), .B1(new_n509), .B2(new_n514), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT25), .B1(new_n519), .B2(new_n307), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n505), .B1(new_n497), .B2(new_n504), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n509), .A2(KEYINPUT74), .A3(new_n514), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n479), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  OAI211_X1 g337(.A(KEYINPUT25), .B(new_n307), .C1(new_n523), .C2(new_n517), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n476), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT75), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n527), .B1(new_n516), .B2(new_n518), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n523), .A2(KEYINPUT75), .A3(new_n517), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n476), .A2(G902), .ZN(new_n531));
  XOR2_X1   g345(.A(new_n531), .B(KEYINPUT76), .Z(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n526), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g349(.A1(G472), .A2(G902), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n308), .A2(new_n188), .A3(G210), .ZN(new_n538));
  XNOR2_X1  g352(.A(new_n538), .B(KEYINPUT27), .ZN(new_n539));
  XNOR2_X1  g353(.A(KEYINPUT26), .B(G101), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n539), .B(new_n540), .Z(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n431), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n386), .A2(G137), .ZN(new_n544));
  OAI21_X1  g358(.A(G131), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n545), .A2(new_n436), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n265), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n437), .A2(new_n272), .A3(new_n273), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n549), .A2(new_n209), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n547), .A2(new_n548), .B1(new_n206), .B2(new_n208), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT28), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n426), .A2(new_n437), .B1(new_n265), .B2(new_n546), .ZN(new_n553));
  INV_X1    g367(.A(new_n209), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT28), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n542), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n547), .A2(new_n548), .A3(KEYINPUT30), .ZN(new_n559));
  XOR2_X1   g373(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n560));
  OAI211_X1 g374(.A(new_n559), .B(new_n209), .C1(new_n553), .C2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT31), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n541), .B1(new_n553), .B2(new_n554), .ZN(new_n563));
  AND3_X1   g377(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n558), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(new_n563), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT69), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT69), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n561), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n567), .A2(KEYINPUT31), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n537), .B1(new_n565), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g385(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT32), .ZN(new_n574));
  AOI211_X1 g388(.A(new_n574), .B(new_n537), .C1(new_n565), .C2(new_n570), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n552), .A2(new_n542), .A3(new_n557), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n561), .A2(new_n555), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n581), .B2(new_n541), .ZN(new_n582));
  AOI211_X1 g396(.A(KEYINPUT71), .B(new_n542), .C1(new_n561), .C2(new_n555), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n579), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n307), .B1(new_n577), .B2(new_n578), .ZN(new_n585));
  OAI21_X1  g399(.A(G472), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n535), .B1(new_n576), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n413), .A2(new_n472), .A3(KEYINPUT94), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n475), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(G101), .ZN(G3));
  INV_X1    g404(.A(KEYINPUT25), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n521), .A2(new_n522), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n517), .B1(new_n592), .B2(new_n480), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n591), .B1(new_n593), .B2(G902), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(new_n524), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n595), .A2(new_n476), .B1(new_n530), .B2(new_n533), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n565), .A2(new_n570), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n307), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n571), .B1(new_n598), .B2(G472), .ZN(new_n599));
  AND3_X1   g413(.A1(new_n472), .A2(new_n596), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n403), .B2(KEYINPUT95), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n401), .B1(new_n390), .B2(new_n398), .ZN(new_n604));
  NOR3_X1   g418(.A1(new_n404), .A2(new_n397), .A3(new_n403), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n603), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n402), .A2(new_n405), .A3(new_n602), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n368), .A2(G902), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT96), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n606), .A2(KEYINPUT96), .A3(new_n607), .A4(new_n608), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT97), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n613), .B1(new_n406), .B2(G478), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n307), .B1(new_n604), .B2(new_n605), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n615), .A2(KEYINPUT97), .A3(new_n368), .ZN(new_n616));
  AOI22_X1  g430(.A1(new_n611), .A2(new_n612), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n367), .ZN(new_n619));
  OAI21_X1  g433(.A(KEYINPUT98), .B1(new_n619), .B2(new_n305), .ZN(new_n620));
  INV_X1    g434(.A(new_n305), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n348), .A2(new_n350), .B1(new_n363), .B2(new_n365), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n617), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n600), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT34), .B(G104), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(KEYINPUT100), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n365), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n630), .B1(new_n365), .B2(KEYINPUT99), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n363), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n365), .A2(KEYINPUT99), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(KEYINPUT100), .ZN(new_n635));
  INV_X1    g449(.A(new_n363), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n365), .A2(KEYINPUT99), .A3(new_n630), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n635), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  AND2_X1   g452(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n621), .A2(new_n639), .A3(new_n351), .A4(new_n412), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n600), .A2(new_n641), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NOR2_X1   g458(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n592), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n592), .A2(new_n645), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n646), .A2(new_n647), .A3(new_n532), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n526), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n599), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT101), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n475), .A2(new_n652), .A3(new_n588), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(KEYINPUT102), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n653), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(new_n476), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n594), .B2(new_n524), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n658), .A2(new_n648), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n659), .B1(new_n576), .B2(new_n586), .ZN(new_n660));
  INV_X1    g474(.A(new_n187), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n291), .A2(new_n301), .ZN(new_n662));
  INV_X1    g476(.A(new_n302), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n291), .A2(new_n301), .A3(new_n302), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n661), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(G900), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n193), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n192), .A2(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g484(.A(new_n670), .B1(new_n348), .B2(new_n350), .ZN(new_n671));
  AND4_X1   g485(.A1(new_n412), .A2(new_n633), .A3(new_n638), .A4(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n660), .A2(new_n472), .A3(new_n666), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  AOI22_X1  g488(.A1(new_n366), .A2(new_n351), .B1(new_n410), .B2(new_n411), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n659), .A2(new_n187), .A3(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(KEYINPUT104), .ZN(new_n678));
  INV_X1    g492(.A(new_n569), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n568), .B1(new_n561), .B2(new_n563), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n550), .A2(new_n551), .ZN(new_n682));
  OAI211_X1 g496(.A(new_n681), .B(G472), .C1(new_n542), .C2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(G472), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n307), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n683), .A2(KEYINPUT103), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n691), .A2(new_n576), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n664), .A2(new_n665), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT38), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n677), .A2(new_n678), .A3(new_n692), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(KEYINPUT105), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n669), .B(KEYINPUT39), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n472), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT40), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(new_n373), .ZN(G45));
  NOR3_X1   g515(.A1(new_n617), .A2(new_n623), .A3(new_n670), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n660), .A2(new_n472), .A3(new_n666), .A4(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G146), .ZN(G48));
  INV_X1    g518(.A(new_n626), .ZN(new_n705));
  INV_X1    g519(.A(new_n415), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n462), .A2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n307), .B1(new_n460), .B2(new_n461), .ZN(new_n708));
  AOI21_X1  g522(.A(KEYINPUT106), .B1(new_n708), .B2(G469), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT106), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT83), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n447), .B1(new_n467), .B2(new_n468), .ZN(new_n712));
  INV_X1    g526(.A(new_n445), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n711), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n714), .A2(new_n459), .A3(new_n446), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n710), .B(new_n416), .C1(new_n715), .C2(new_n307), .ZN(new_n716));
  OAI211_X1 g530(.A(new_n587), .B(new_n707), .C1(new_n709), .C2(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n705), .A2(new_n717), .ZN(new_n718));
  XOR2_X1   g532(.A(KEYINPUT41), .B(G113), .Z(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NOR2_X1   g534(.A1(new_n717), .A2(new_n640), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(new_n202), .ZN(G18));
  INV_X1    g536(.A(KEYINPUT107), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n707), .B1(new_n716), .B2(new_n709), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n660), .A2(new_n413), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n723), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n462), .A2(new_n706), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n708), .A2(G469), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(new_n710), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n708), .A2(KEYINPUT106), .A3(G469), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n571), .A2(KEYINPUT32), .ZN(new_n732));
  OAI211_X1 g546(.A(new_n586), .B(new_n732), .C1(new_n571), .C2(new_n572), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n367), .A2(new_n412), .ZN(new_n734));
  AND4_X1   g548(.A1(new_n733), .A2(new_n621), .A3(new_n734), .A4(new_n650), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n731), .A2(KEYINPUT107), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n726), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G119), .ZN(G21));
  NAND2_X1  g552(.A1(new_n367), .A2(new_n412), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n305), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT108), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n598), .A2(new_n741), .A3(G472), .ZN(new_n742));
  AOI21_X1  g556(.A(G902), .B1(new_n565), .B2(new_n570), .ZN(new_n743));
  OAI21_X1  g557(.A(KEYINPUT108), .B1(new_n743), .B2(new_n684), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n597), .A2(new_n536), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n740), .A2(new_n596), .A3(new_n742), .A4(new_n746), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT109), .B1(new_n724), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n729), .A2(new_n730), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n596), .A2(new_n745), .A3(new_n742), .A4(new_n744), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n666), .A2(new_n196), .A3(new_n675), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT109), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n749), .A2(new_n752), .A3(new_n753), .A4(new_n707), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  OAI211_X1 g570(.A(new_n707), .B(new_n666), .C1(new_n716), .C2(new_n709), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n746), .A2(new_n702), .A3(new_n650), .A4(new_n742), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n267), .ZN(G27));
  INV_X1    g574(.A(KEYINPUT42), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n664), .A2(new_n187), .A3(new_n665), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n415), .B(new_n762), .C1(new_n462), .C2(new_n471), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n745), .A2(new_n574), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n764), .A2(new_n586), .A3(new_n732), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n702), .A2(new_n765), .A3(new_n596), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n761), .B1(new_n763), .B2(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(new_n762), .ZN(new_n768));
  NOR4_X1   g582(.A1(new_n617), .A2(new_n623), .A3(KEYINPUT42), .A4(new_n670), .ZN(new_n769));
  AND4_X1   g583(.A1(new_n587), .A2(new_n472), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n767), .A2(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(G131), .ZN(G33));
  AND3_X1   g586(.A1(new_n587), .A2(new_n472), .A3(new_n768), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n672), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  XNOR2_X1  g589(.A(new_n623), .B(KEYINPUT111), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT43), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n617), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(KEYINPUT112), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n776), .A2(new_n781), .A3(new_n778), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n777), .B1(new_n617), .B2(new_n367), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT113), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n783), .A2(KEYINPUT113), .A3(new_n784), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n659), .A2(new_n599), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT44), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n787), .A2(KEYINPUT44), .A3(new_n788), .A4(new_n789), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n792), .A2(new_n768), .A3(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n463), .ZN(new_n795));
  AND2_X1   g609(.A1(new_n470), .A2(KEYINPUT45), .ZN(new_n796));
  OAI21_X1  g610(.A(G469), .B1(new_n470), .B2(KEYINPUT45), .ZN(new_n797));
  OAI211_X1 g611(.A(KEYINPUT46), .B(new_n795), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n462), .ZN(new_n799));
  OR2_X1    g613(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n799), .A2(KEYINPUT110), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n796), .A2(new_n797), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n463), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n800), .B(new_n801), .C1(new_n803), .C2(KEYINPUT46), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n706), .A3(new_n697), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n794), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G137), .ZN(G39));
  NAND3_X1  g621(.A1(new_n618), .A2(new_n367), .A3(new_n669), .ZN(new_n808));
  NOR4_X1   g622(.A1(new_n808), .A2(new_n733), .A3(new_n596), .A4(new_n762), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n804), .A2(new_n706), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT47), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n804), .A2(KEYINPUT47), .A3(new_n706), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n810), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(new_n321), .ZN(G42));
  NAND2_X1  g630(.A1(new_n749), .A2(new_n462), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n817), .B(KEYINPUT115), .Z(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(new_n415), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n813), .A3(new_n814), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n750), .A2(new_n192), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n820), .A2(new_n768), .A3(new_n785), .A4(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n785), .A2(new_n821), .ZN(new_n823));
  OR3_X1    g637(.A1(new_n724), .A2(new_n187), .A3(new_n694), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OR2_X1    g639(.A1(new_n825), .A2(KEYINPUT50), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(KEYINPUT50), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n742), .A2(new_n745), .A3(new_n744), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n828), .A2(new_n659), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n724), .A2(new_n192), .A3(new_n762), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n785), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n826), .A2(new_n827), .B1(new_n829), .B2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(new_n830), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n691), .A2(new_n576), .A3(new_n596), .ZN(new_n834));
  OR3_X1    g648(.A1(new_n833), .A2(KEYINPUT119), .A3(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(KEYINPUT119), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n835), .A2(new_n623), .A3(new_n617), .A4(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n822), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n822), .A2(new_n832), .A3(KEYINPUT51), .A4(new_n837), .ZN(new_n841));
  INV_X1    g655(.A(new_n189), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT120), .ZN(new_n843));
  OR3_X1    g657(.A1(new_n823), .A2(new_n843), .A3(new_n757), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n843), .B1(new_n823), .B2(new_n757), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n842), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n765), .A2(new_n596), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n831), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT48), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT48), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n831), .A2(new_n850), .A3(new_n847), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n835), .A2(new_n624), .A3(new_n836), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n846), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT121), .ZN(new_n855));
  AND2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n855), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n840), .B(new_n841), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n587), .B(new_n731), .C1(new_n626), .C2(new_n641), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n737), .A2(new_n755), .A3(new_n771), .A4(new_n859), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n671), .A2(new_n410), .A3(new_n411), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n733), .A2(new_n639), .A3(new_n650), .A4(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n758), .A2(new_n862), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n773), .A2(new_n672), .B1(new_n863), .B2(new_n763), .ZN(new_n864));
  INV_X1    g678(.A(new_n412), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n619), .B1(new_n865), .B2(new_n367), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n600), .A2(new_n621), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n864), .A2(new_n589), .A3(new_n653), .A4(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n860), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT52), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n462), .A2(new_n471), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n187), .B1(new_n303), .B2(new_n304), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n739), .ZN(new_n873));
  NOR4_X1   g687(.A1(new_n658), .A2(new_n415), .A3(new_n648), .A4(new_n670), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n692), .A2(new_n871), .A3(new_n873), .A4(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n673), .A2(new_n703), .A3(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n870), .B1(new_n876), .B2(new_n759), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n808), .A2(new_n828), .A3(new_n659), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n731), .A2(new_n666), .A3(new_n878), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n733), .A2(new_n666), .A3(new_n650), .ZN(new_n880));
  OAI211_X1 g694(.A(new_n880), .B(new_n472), .C1(new_n672), .C2(new_n702), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n879), .A2(KEYINPUT52), .A3(new_n881), .A4(new_n875), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n877), .A2(KEYINPUT117), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT117), .B1(new_n877), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n869), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT53), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT116), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n877), .A2(new_n887), .A3(new_n882), .ZN(new_n888));
  OAI211_X1 g702(.A(KEYINPUT116), .B(new_n870), .C1(new_n876), .C2(new_n759), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n890), .A2(new_n891), .A3(new_n869), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n886), .A2(KEYINPUT54), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n885), .A2(new_n891), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n868), .A2(new_n891), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n860), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n717), .B1(new_n705), .B2(new_n640), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n726), .B2(new_n736), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n899), .A2(KEYINPUT118), .A3(new_n755), .A4(new_n771), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n890), .A2(new_n895), .A3(new_n897), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT54), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n894), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n893), .A2(new_n903), .ZN(new_n904));
  OAI22_X1  g718(.A1(new_n858), .A2(new_n904), .B1(G952), .B2(G953), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT49), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n818), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n818), .A2(new_n906), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n776), .A2(new_n706), .A3(new_n187), .A4(new_n618), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n909), .A2(new_n535), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(KEYINPUT114), .ZN(new_n912));
  AOI211_X1 g726(.A(new_n692), .B(new_n694), .C1(new_n911), .C2(KEYINPUT114), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n907), .A2(new_n908), .A3(new_n912), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n905), .A2(new_n914), .ZN(G75));
  INV_X1    g729(.A(KEYINPUT56), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n295), .A2(new_n297), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n300), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT55), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n900), .A2(new_n897), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n895), .A2(new_n889), .A3(new_n888), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n877), .A2(new_n882), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT117), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n877), .A2(KEYINPUT117), .A3(new_n882), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT53), .B1(new_n928), .B2(new_n869), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n923), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(G210), .A2(G902), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n916), .B(new_n920), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n894), .B2(new_n901), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n919), .B1(new_n933), .B2(KEYINPUT56), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n188), .A2(G952), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT122), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n932), .A2(new_n934), .A3(KEYINPUT122), .A4(new_n936), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n940), .ZN(G51));
  NAND2_X1  g755(.A1(new_n894), .A2(new_n901), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n942), .A2(KEYINPUT54), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(new_n903), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n463), .B(KEYINPUT57), .Z(new_n945));
  OAI21_X1  g759(.A(new_n715), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n930), .A2(new_n307), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n802), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n935), .B1(new_n946), .B2(new_n948), .ZN(G54));
  NAND3_X1  g763(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .ZN(new_n950));
  OR2_X1    g764(.A1(new_n345), .A2(new_n361), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .A4(new_n951), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n953), .A2(new_n954), .A3(new_n936), .ZN(G60));
  NAND2_X1  g769(.A1(G478), .A2(G902), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n956), .B(KEYINPUT59), .Z(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n904), .A2(new_n958), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT123), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n606), .A2(new_n607), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n959), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n943), .A2(new_n903), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n957), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n935), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n957), .B1(new_n893), .B2(new_n903), .ZN(new_n966));
  INV_X1    g780(.A(new_n961), .ZN(new_n967));
  OAI21_X1  g781(.A(KEYINPUT123), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AND3_X1   g782(.A1(new_n962), .A2(new_n965), .A3(new_n968), .ZN(G63));
  NAND2_X1  g783(.A1(G217), .A2(G902), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n970), .B(KEYINPUT60), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g786(.A(new_n972), .B1(new_n923), .B2(new_n929), .ZN(new_n973));
  INV_X1    g787(.A(new_n530), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n935), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT124), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n646), .A2(new_n647), .ZN(new_n977));
  AND4_X1   g791(.A1(new_n976), .A2(new_n942), .A3(new_n977), .A4(new_n972), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n971), .B1(new_n894), .B2(new_n901), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n976), .B1(new_n979), .B2(new_n977), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n975), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT61), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  OAI211_X1 g797(.A(KEYINPUT61), .B(new_n975), .C1(new_n978), .C2(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G66));
  AND2_X1   g799(.A1(new_n589), .A2(new_n867), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n899), .A2(new_n653), .A3(new_n755), .A4(new_n986), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n987), .A2(new_n188), .ZN(new_n988));
  OAI21_X1  g802(.A(G953), .B1(new_n279), .B2(new_n194), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n917), .B1(G898), .B2(new_n188), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT125), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n990), .B(new_n992), .ZN(G69));
  OAI21_X1  g807(.A(new_n559), .B1(new_n553), .B2(new_n560), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n994), .B(KEYINPUT126), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(KEYINPUT127), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(new_n358), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT62), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n879), .A2(new_n881), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n700), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(new_n999), .ZN(new_n1001));
  OAI211_X1 g815(.A(KEYINPUT62), .B(new_n1001), .C1(new_n696), .C2(new_n699), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n815), .B1(new_n1000), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n698), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n1004), .A2(new_n587), .A3(new_n768), .A4(new_n866), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1003), .A2(new_n806), .A3(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n997), .B1(new_n1006), .B2(new_n188), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n997), .B1(new_n667), .B2(new_n188), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n847), .A2(new_n873), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n805), .B1(new_n794), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1001), .A2(new_n771), .A3(new_n774), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n815), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1008), .B1(new_n1013), .B2(new_n188), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1015));
  OR3_X1    g829(.A1(new_n1007), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1015), .B1(new_n1007), .B2(new_n1014), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1016), .A2(new_n1017), .ZN(G72));
  XNOR2_X1  g832(.A(new_n685), .B(KEYINPUT63), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1019), .B1(new_n1006), .B2(new_n987), .ZN(new_n1020));
  INV_X1    g834(.A(new_n581), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n541), .ZN(new_n1022));
  NAND2_X1  g836(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1019), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n582), .A2(new_n583), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(new_n681), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n886), .A2(new_n892), .A3(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n1010), .A2(new_n1012), .A3(new_n987), .ZN(new_n1028));
  OAI211_X1 g842(.A(new_n541), .B(new_n1021), .C1(new_n1028), .C2(new_n1024), .ZN(new_n1029));
  AND4_X1   g843(.A1(new_n936), .A2(new_n1023), .A3(new_n1027), .A4(new_n1029), .ZN(G57));
endmodule


