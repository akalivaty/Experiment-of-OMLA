//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 0 1 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n578, new_n579, new_n580, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT65), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NAND2_X1  g046(.A1(G101), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n472), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  AND2_X1   g052(.A1(new_n465), .A2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(new_n475), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  OR3_X1    g055(.A1(new_n479), .A2(KEYINPUT66), .A3(new_n480), .ZN(new_n481));
  OAI21_X1  g056(.A(KEYINPUT66), .B1(new_n479), .B2(new_n480), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n468), .A2(new_n475), .ZN(new_n483));
  AOI22_X1  g058(.A1(new_n481), .A2(new_n482), .B1(G124), .B2(new_n483), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n486));
  AND2_X1   g061(.A1(new_n484), .A2(new_n486), .ZN(G162));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  INV_X1    g063(.A(G126), .ZN(new_n489));
  OAI21_X1  g064(.A(new_n488), .B1(new_n468), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n464), .A2(G2105), .ZN(new_n491));
  AOI22_X1  g066(.A1(new_n490), .A2(G2105), .B1(G102), .B2(new_n491), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n475), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(G164));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT5), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n502), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NOR2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n498), .B(new_n500), .C1(new_n506), .C2(new_n507), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n505), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  INV_X1    g091(.A(G51), .ZN(new_n517));
  INV_X1    g092(.A(G89), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n509), .A2(new_n517), .B1(new_n518), .B2(new_n512), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n499), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n497), .A2(KEYINPUT5), .ZN(new_n522));
  OAI21_X1  g097(.A(KEYINPUT67), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n498), .A2(new_n500), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n526), .A2(G63), .A3(G651), .ZN(new_n527));
  AND2_X1   g102(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n529));
  OAI211_X1 g104(.A(new_n516), .B(new_n520), .C1(new_n528), .C2(new_n529), .ZN(G286));
  INV_X1    g105(.A(G286), .ZN(G168));
  NAND2_X1  g106(.A1(G77), .A2(G543), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n533), .B1(new_n526), .B2(G64), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT69), .B1(new_n534), .B2(new_n504), .ZN(new_n535));
  INV_X1    g110(.A(G52), .ZN(new_n536));
  INV_X1    g111(.A(G90), .ZN(new_n537));
  OAI22_X1  g112(.A1(new_n509), .A2(new_n536), .B1(new_n537), .B2(new_n512), .ZN(new_n538));
  INV_X1    g113(.A(new_n538), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n498), .A2(new_n500), .A3(new_n524), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n524), .B1(new_n498), .B2(new_n500), .ZN(new_n541));
  OAI21_X1  g116(.A(G64), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(new_n532), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT69), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(new_n544), .A3(G651), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n535), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(G171));
  INV_X1    g122(.A(G43), .ZN(new_n548));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n509), .A2(new_n548), .B1(new_n549), .B2(new_n512), .ZN(new_n550));
  INV_X1    g125(.A(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n526), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n551), .B1(new_n504), .B2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT70), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n556), .A2(new_n560), .ZN(G188));
  NAND2_X1  g136(.A1(G78), .A2(G543), .ZN(new_n562));
  XOR2_X1   g137(.A(new_n562), .B(KEYINPUT71), .Z(new_n563));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n501), .B(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n563), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n512), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n567), .A2(G651), .B1(G91), .B2(new_n568), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n508), .A2(G53), .A3(G543), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT9), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(G299));
  NAND2_X1  g147(.A1(new_n546), .A2(KEYINPUT73), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT73), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n535), .A2(new_n545), .A3(new_n574), .A4(new_n539), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n573), .A2(new_n575), .ZN(G301));
  INV_X1    g151(.A(G166), .ZN(G303));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n509), .A2(new_n578), .B1(new_n579), .B2(new_n512), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n526), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  NAND2_X1  g158(.A1(G73), .A2(G543), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT74), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n498), .A2(new_n500), .A3(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n504), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI211_X1 g162(.A(G48), .B(G543), .C1(new_n506), .C2(new_n507), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n512), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n526), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n504), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n509), .A2(new_n595), .B1(new_n596), .B2(new_n512), .ZN(new_n597));
  OR3_X1    g172(.A1(new_n594), .A2(KEYINPUT75), .A3(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT75), .B1(new_n594), .B2(new_n597), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G290));
  NAND2_X1  g175(.A1(G301), .A2(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(G79), .A2(G543), .ZN(new_n602));
  INV_X1    g177(.A(G66), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n565), .B2(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(new_n509), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n604), .A2(G651), .B1(G54), .B2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(G92), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n512), .A2(new_n607), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(KEYINPUT76), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G284));
  OAI21_X1  g187(.A(new_n601), .B1(new_n611), .B2(G868), .ZN(G321));
  NAND2_X1  g188(.A1(G286), .A2(G868), .ZN(new_n614));
  INV_X1    g189(.A(G299), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G297));
  OAI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(G868), .ZN(G280));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n611), .B1(new_n618), .B2(G860), .ZN(G148));
  INV_X1    g194(.A(G868), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n553), .A2(new_n620), .ZN(new_n621));
  AND2_X1   g196(.A1(new_n611), .A2(new_n618), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(new_n620), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g199(.A1(new_n475), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT12), .Z(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT13), .Z(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n483), .A2(G123), .ZN(new_n629));
  NOR2_X1   g204(.A1(new_n468), .A2(G2105), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(G135), .ZN(new_n631));
  NOR2_X1   g206(.A1(G99), .A2(G2105), .ZN(new_n632));
  OAI21_X1  g207(.A(G2104), .B1(new_n475), .B2(G111), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n629), .B(new_n631), .C1(new_n632), .C2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2096), .Z(new_n635));
  NAND2_X1  g210(.A1(new_n628), .A2(new_n635), .ZN(G156));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XOR2_X1   g213(.A(G2443), .B(G2446), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(G2427), .B(G2438), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2430), .ZN(new_n644));
  XOR2_X1   g219(.A(KEYINPUT15), .B(G2435), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(KEYINPUT14), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n642), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n648), .A2(G14), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(KEYINPUT77), .ZN(G401));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT17), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT78), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  NAND3_X1  g230(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT79), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n654), .A2(new_n651), .ZN(new_n658));
  INV_X1    g233(.A(new_n655), .ZN(new_n659));
  OAI211_X1 g234(.A(new_n658), .B(new_n659), .C1(new_n652), .C2(new_n654), .ZN(new_n660));
  INV_X1    g235(.A(new_n651), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n661), .A2(new_n655), .A3(new_n653), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(KEYINPUT18), .Z(new_n663));
  NAND3_X1  g238(.A1(new_n657), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2096), .B(G2100), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT80), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n664), .B(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(G227));
  XNOR2_X1  g243(.A(G1971), .B(G1976), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT19), .ZN(new_n670));
  XOR2_X1   g245(.A(G1956), .B(G2474), .Z(new_n671));
  XOR2_X1   g246(.A(G1961), .B(G1966), .Z(new_n672));
  NAND2_X1  g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(new_n670), .ZN(new_n675));
  NOR2_X1   g250(.A1(new_n671), .A2(new_n672), .ZN(new_n676));
  AOI22_X1  g251(.A1(new_n674), .A2(KEYINPUT20), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n676), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n678), .A2(new_n670), .A3(new_n673), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n677), .B(new_n679), .C1(KEYINPUT20), .C2(new_n674), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1986), .B(G1996), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(G1981), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1991), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n682), .B(new_n685), .ZN(G229));
  AND2_X1   g261(.A1(KEYINPUT81), .A2(G16), .ZN(new_n687));
  NOR2_X1   g262(.A1(KEYINPUT81), .A2(G16), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G24), .ZN(new_n691));
  INV_X1    g266(.A(G290), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n691), .B1(new_n692), .B2(new_n690), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(G1986), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(G1986), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G119), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n630), .A2(G131), .ZN(new_n697));
  OR2_X1    g272(.A1(G95), .A2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n698), .B(G2104), .C1(G107), .C2(new_n475), .ZN(new_n699));
  NAND3_X1  g274(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  MUX2_X1   g275(.A(G25), .B(new_n700), .S(G29), .Z(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT35), .B(G1991), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n695), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G6), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n591), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT82), .ZN(new_n708));
  XOR2_X1   g283(.A(KEYINPUT32), .B(G1981), .Z(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n708), .A2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n690), .A2(G22), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(G166), .B2(new_n690), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n710), .B(new_n711), .C1(G1971), .C2(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n705), .A2(G23), .ZN(new_n715));
  AND2_X1   g290(.A1(new_n581), .A2(new_n582), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n705), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT33), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1976), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n714), .B(new_n719), .C1(G1971), .C2(new_n713), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n694), .B(new_n704), .C1(new_n720), .C2(KEYINPUT34), .ZN(new_n721));
  OAI221_X1 g296(.A(new_n721), .B1(KEYINPUT34), .B2(new_n720), .C1(new_n702), .C2(new_n701), .ZN(new_n722));
  NAND2_X1  g297(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n723));
  OR2_X1    g298(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n705), .A2(G5), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n725), .B1(G171), .B2(new_n705), .ZN(new_n726));
  INV_X1    g301(.A(G1961), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(KEYINPUT83), .A2(KEYINPUT36), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n722), .A2(new_n723), .A3(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n554), .A2(new_n690), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G19), .B2(new_n690), .ZN(new_n732));
  INV_X1    g307(.A(G1341), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G1966), .ZN(new_n735));
  NAND2_X1  g310(.A1(G168), .A2(G16), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(G16), .B2(G21), .ZN(new_n737));
  INV_X1    g312(.A(G29), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G33), .ZN(new_n739));
  AOI22_X1  g314(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n740));
  NOR2_X1   g315(.A1(new_n740), .A2(new_n475), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n630), .A2(G139), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n491), .A2(G103), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT25), .ZN(new_n744));
  NOR3_X1   g319(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT87), .Z(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n739), .B1(new_n747), .B2(new_n738), .ZN(new_n748));
  OAI221_X1 g323(.A(new_n734), .B1(new_n735), .B2(new_n737), .C1(new_n748), .C2(G2072), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n735), .B2(new_n737), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n738), .A2(G27), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(G164), .B2(new_n738), .ZN(new_n752));
  INV_X1    g327(.A(G2078), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND4_X1  g329(.A1(new_n465), .A2(new_n467), .A3(G129), .A4(G2105), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT88), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XOR2_X1   g332(.A(new_n757), .B(KEYINPUT26), .Z(new_n758));
  AOI22_X1  g333(.A1(new_n630), .A2(G141), .B1(G105), .B2(new_n491), .ZN(new_n759));
  AND3_X1   g334(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(G29), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(KEYINPUT89), .C1(G29), .C2(G32), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(KEYINPUT89), .B2(new_n761), .ZN(new_n763));
  XNOR2_X1  g338(.A(KEYINPUT27), .B(G1996), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(KEYINPUT24), .A2(G34), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  NOR2_X1   g342(.A1(KEYINPUT24), .A2(G34), .ZN(new_n768));
  NOR3_X1   g343(.A1(new_n767), .A2(new_n768), .A3(G29), .ZN(new_n769));
  INV_X1    g344(.A(G160), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n769), .B1(new_n770), .B2(G29), .ZN(new_n771));
  INV_X1    g346(.A(G2084), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT30), .B(G28), .Z(new_n774));
  MUX2_X1   g349(.A(new_n774), .B(new_n634), .S(G29), .Z(new_n775));
  XNOR2_X1  g350(.A(KEYINPUT31), .B(G11), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n771), .A2(new_n772), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n773), .A2(new_n775), .A3(new_n776), .A4(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n732), .A2(new_n733), .ZN(new_n779));
  AOI211_X1 g354(.A(new_n778), .B(new_n779), .C1(G2072), .C2(new_n748), .ZN(new_n780));
  NAND4_X1  g355(.A1(new_n750), .A2(new_n754), .A3(new_n765), .A4(new_n780), .ZN(new_n781));
  NOR2_X1   g356(.A1(G4), .A2(G16), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(new_n611), .B2(G16), .ZN(new_n783));
  INV_X1    g358(.A(G1348), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n690), .A2(KEYINPUT23), .A3(G20), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n787));
  INV_X1    g362(.A(G20), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n689), .B2(new_n788), .ZN(new_n789));
  OAI211_X1 g364(.A(new_n786), .B(new_n789), .C1(new_n615), .C2(new_n705), .ZN(new_n790));
  INV_X1    g365(.A(G1956), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n738), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n738), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT29), .B(G2090), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n785), .A2(new_n792), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n738), .A2(G26), .ZN(new_n798));
  OR2_X1    g373(.A1(G104), .A2(G2105), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n799), .B(G2104), .C1(G116), .C2(new_n475), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT85), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT84), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n478), .A2(new_n802), .A3(G128), .A4(G2105), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n465), .A2(new_n467), .A3(G128), .A4(G2105), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT84), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n630), .A2(G140), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n801), .A2(new_n806), .A3(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n803), .A2(new_n805), .B1(G140), .B2(new_n630), .ZN(new_n811));
  NAND3_X1  g386(.A1(new_n811), .A2(KEYINPUT86), .A3(new_n801), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n798), .B1(new_n814), .B2(new_n738), .ZN(new_n815));
  MUX2_X1   g390(.A(new_n798), .B(new_n815), .S(KEYINPUT28), .Z(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(G2067), .ZN(new_n817));
  NOR3_X1   g392(.A1(new_n781), .A2(new_n797), .A3(new_n817), .ZN(new_n818));
  NAND4_X1  g393(.A1(new_n724), .A2(new_n728), .A3(new_n730), .A4(new_n818), .ZN(G150));
  INV_X1    g394(.A(G150), .ZN(G311));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  OAI22_X1  g397(.A1(new_n509), .A2(new_n821), .B1(new_n822), .B2(new_n512), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n526), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n504), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT92), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n824), .B(KEYINPUT92), .C1(new_n504), .C2(new_n825), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(G860), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT37), .Z(new_n831));
  NAND2_X1  g406(.A1(new_n611), .A2(G559), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT91), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT39), .ZN(new_n834));
  INV_X1    g409(.A(new_n826), .ZN(new_n835));
  NOR2_X1   g410(.A1(new_n835), .A2(new_n553), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(new_n829), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n553), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n834), .B(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(KEYINPUT90), .B(KEYINPUT38), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n839), .B(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n831), .B1(new_n841), .B2(G860), .ZN(G145));
  XOR2_X1   g417(.A(G160), .B(new_n634), .Z(new_n843));
  XOR2_X1   g418(.A(new_n843), .B(G162), .Z(new_n844));
  AND3_X1   g419(.A1(new_n811), .A2(KEYINPUT86), .A3(new_n801), .ZN(new_n845));
  AOI21_X1  g420(.A(KEYINPUT86), .B1(new_n811), .B2(new_n801), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n760), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n756), .A2(new_n758), .A3(new_n759), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n810), .A2(new_n848), .A3(new_n812), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT93), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n492), .A2(new_n494), .A3(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n850), .B1(new_n492), .B2(new_n494), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AND3_X1   g429(.A1(new_n847), .A2(new_n849), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n847), .B2(new_n849), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n747), .B1(new_n855), .B2(new_n856), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n630), .A2(KEYINPUT94), .A3(G142), .ZN(new_n858));
  AND2_X1   g433(.A1(new_n483), .A2(G130), .ZN(new_n859));
  AOI21_X1  g434(.A(KEYINPUT94), .B1(new_n630), .B2(G142), .ZN(new_n860));
  NOR3_X1   g435(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  OR2_X1    g436(.A1(G106), .A2(G2105), .ZN(new_n862));
  OAI211_X1 g437(.A(new_n862), .B(G2104), .C1(G118), .C2(new_n475), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n861), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n700), .A2(new_n626), .ZN(new_n865));
  INV_X1    g440(.A(new_n626), .ZN(new_n866));
  NAND4_X1  g441(.A1(new_n866), .A2(new_n696), .A3(new_n697), .A4(new_n699), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n864), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n861), .A2(new_n865), .A3(new_n867), .A4(new_n863), .ZN(new_n870));
  AND3_X1   g445(.A1(new_n869), .A2(KEYINPUT95), .A3(new_n870), .ZN(new_n871));
  AOI21_X1  g446(.A(KEYINPUT95), .B1(new_n869), .B2(new_n870), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n853), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n874), .A2(new_n851), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n845), .A2(new_n846), .A3(new_n760), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n848), .B1(new_n810), .B2(new_n812), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(new_n745), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n847), .A2(new_n849), .A3(new_n854), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  AND3_X1   g456(.A1(new_n857), .A2(new_n873), .A3(new_n881), .ZN(new_n882));
  AOI21_X1  g457(.A(new_n873), .B1(new_n857), .B2(new_n881), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n844), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  INV_X1    g460(.A(new_n844), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n869), .A2(new_n870), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n887), .B1(new_n857), .B2(new_n881), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n888), .B2(KEYINPUT96), .ZN(new_n889));
  INV_X1    g464(.A(new_n887), .ZN(new_n890));
  NOR3_X1   g465(.A1(new_n855), .A2(new_n856), .A3(new_n745), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n746), .B1(new_n878), .B2(new_n880), .ZN(new_n892));
  OAI211_X1 g467(.A(KEYINPUT96), .B(new_n890), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n857), .A2(new_n873), .A3(new_n881), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n884), .B(new_n885), .C1(new_n889), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n896), .A2(KEYINPUT97), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n898));
  INV_X1    g473(.A(KEYINPUT96), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n900), .A2(new_n894), .A3(new_n886), .A4(new_n893), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT97), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n901), .A2(new_n902), .A3(new_n885), .A4(new_n884), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n897), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g480(.A(new_n838), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n622), .B(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(G299), .A2(new_n610), .ZN(new_n908));
  NAND4_X1  g483(.A1(new_n569), .A2(new_n606), .A3(new_n571), .A4(new_n609), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n907), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n908), .A2(new_n914), .A3(new_n909), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n914), .B1(new_n908), .B2(new_n909), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT98), .B1(new_n910), .B2(KEYINPUT41), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n912), .B1(new_n907), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g496(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(KEYINPUT42), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g499(.A(G288), .B(G166), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(new_n591), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(G290), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  NOR3_X1   g504(.A1(new_n922), .A2(new_n923), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(G868), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(G868), .B2(new_n837), .ZN(G295));
  OAI21_X1  g507(.A(new_n931), .B1(G868), .B2(new_n837), .ZN(G331));
  INV_X1    g508(.A(KEYINPUT99), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n934), .B1(G301), .B2(G168), .ZN(new_n935));
  AOI211_X1 g510(.A(KEYINPUT99), .B(G286), .C1(new_n573), .C2(new_n575), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(G168), .A2(new_n546), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n906), .B1(new_n937), .B2(new_n939), .ZN(new_n940));
  NOR4_X1   g515(.A1(new_n935), .A2(new_n936), .A3(new_n838), .A4(new_n938), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n911), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(G301), .A2(G168), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT99), .ZN(new_n944));
  NAND3_X1  g519(.A1(G301), .A2(new_n934), .A3(G168), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n939), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n946), .A2(new_n838), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n937), .A2(new_n906), .A3(new_n939), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n947), .A2(new_n919), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n927), .B1(new_n942), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n942), .A2(new_n927), .A3(new_n949), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT100), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g528(.A1(new_n942), .A2(new_n949), .A3(KEYINPUT100), .A4(new_n927), .ZN(new_n954));
  AOI211_X1 g529(.A(G37), .B(new_n950), .C1(new_n953), .C2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  AOI21_X1  g531(.A(G37), .B1(new_n953), .B2(new_n954), .ZN(new_n957));
  OR2_X1    g532(.A1(new_n915), .A2(new_n916), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n947), .A2(new_n948), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(KEYINPUT101), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT101), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n947), .A2(new_n948), .A3(new_n961), .A4(new_n958), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n960), .A2(new_n942), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n929), .ZN(new_n964));
  AND3_X1   g539(.A1(new_n957), .A2(KEYINPUT43), .A3(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT44), .B1(new_n956), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n953), .A2(new_n954), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT43), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n967), .A2(new_n964), .A3(new_n968), .A4(new_n885), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n969), .B1(new_n955), .B2(new_n968), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n966), .B1(new_n971), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n495), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n977));
  XNOR2_X1  g552(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n976), .B(new_n977), .C1(new_n978), .C2(new_n974), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n735), .ZN(new_n980));
  OR2_X1    g555(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n974), .A2(KEYINPUT50), .ZN(new_n982));
  NAND4_X1  g557(.A1(new_n981), .A2(new_n772), .A3(new_n977), .A4(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(G8), .A3(G286), .ZN(new_n985));
  NAND2_X1  g560(.A1(G286), .A2(G8), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n986), .B1(KEYINPUT122), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(G8), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n980), .B2(new_n983), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT121), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  AOI211_X1 g567(.A(KEYINPUT121), .B(new_n989), .C1(new_n980), .C2(new_n983), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n988), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n986), .A2(KEYINPUT122), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT51), .B(new_n985), .C1(new_n994), .C2(new_n995), .ZN(new_n996));
  OR2_X1    g571(.A1(new_n990), .A2(new_n988), .ZN(new_n997));
  OAI211_X1 g572(.A(KEYINPUT45), .B(new_n973), .C1(new_n852), .C2(new_n853), .ZN(new_n998));
  INV_X1    g573(.A(new_n977), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n974), .B2(new_n978), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n998), .A2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT105), .B1(new_n1001), .B2(G1971), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT106), .B(G2090), .Z(new_n1003));
  NAND4_X1  g578(.A1(new_n981), .A2(new_n977), .A3(new_n982), .A4(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1971), .B1(new_n998), .B2(new_n1000), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT105), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT55), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1009), .B1(G166), .B2(new_n989), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT107), .ZN(new_n1011));
  NAND3_X1  g586(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1013), .B(new_n1009), .C1(G166), .C2(new_n989), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1011), .A2(new_n1012), .A3(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT108), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1008), .A2(new_n1016), .A3(G8), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1004), .ZN(new_n1018));
  OAI21_X1  g593(.A(G8), .B1(new_n1018), .B2(new_n1005), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1015), .ZN(new_n1020));
  INV_X1    g595(.A(G1981), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n591), .A2(new_n1021), .ZN(new_n1022));
  OAI21_X1  g597(.A(G1981), .B1(new_n587), .B2(new_n590), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT49), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n977), .A2(new_n495), .A3(new_n973), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1022), .A2(KEYINPUT49), .A3(new_n1023), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1026), .A2(G8), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n581), .A2(G1976), .A3(new_n582), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1027), .A2(G8), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT52), .ZN(new_n1032));
  XNOR2_X1  g607(.A(KEYINPUT109), .B(G1976), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT52), .B1(G288), .B2(new_n1033), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1034), .A2(new_n1027), .A3(G8), .A4(new_n1030), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1029), .A2(new_n1032), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT113), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT113), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1029), .A2(new_n1032), .A3(new_n1035), .A4(new_n1038), .ZN(new_n1039));
  AOI22_X1  g614(.A1(new_n1019), .A2(new_n1020), .B1(new_n1037), .B2(new_n1039), .ZN(new_n1040));
  AND2_X1   g615(.A1(new_n1017), .A2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n996), .A2(new_n997), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1001), .A2(new_n753), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n981), .A2(new_n977), .A3(new_n982), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1043), .A2(new_n1044), .B1(new_n727), .B2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n753), .A2(KEYINPUT53), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n875), .A2(new_n973), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1048), .B2(new_n978), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1049), .A2(new_n977), .A3(new_n998), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1051), .A2(KEYINPUT125), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT125), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1046), .A2(new_n1053), .A3(new_n1050), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1052), .A2(G171), .A3(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1046), .B1(new_n1047), .B2(new_n979), .ZN(new_n1056));
  INV_X1    g631(.A(G301), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g633(.A(KEYINPUT54), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g634(.A1(new_n1051), .A2(new_n1057), .ZN(new_n1060));
  AOI21_X1  g635(.A(KEYINPUT54), .B1(new_n1060), .B2(KEYINPUT124), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(KEYINPUT123), .A3(new_n1057), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT123), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(KEYINPUT124), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1066), .B1(new_n1051), .B2(new_n1057), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1061), .A2(new_n1062), .A3(new_n1065), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1042), .B1(new_n1059), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  XNOR2_X1  g645(.A(KEYINPUT56), .B(G2072), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1001), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1045), .A2(new_n791), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  XOR2_X1   g650(.A(G299), .B(KEYINPUT57), .Z(new_n1076));
  AND2_X1   g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1070), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1074), .B(new_n1076), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1080), .A2(KEYINPUT61), .ZN(new_n1081));
  INV_X1    g656(.A(G2067), .ZN(new_n1082));
  INV_X1    g657(.A(new_n1027), .ZN(new_n1083));
  AOI22_X1  g658(.A1(new_n1045), .A2(new_n784), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AND2_X1   g659(.A1(new_n1084), .A2(new_n610), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n610), .ZN(new_n1086));
  OAI21_X1  g661(.A(KEYINPUT60), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n610), .A2(KEYINPUT60), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1084), .A2(new_n1088), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1079), .A2(new_n1081), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  AND2_X1   g667(.A1(new_n1027), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT117), .B(G1996), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n998), .A2(new_n1000), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(KEYINPUT118), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT118), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n998), .A2(new_n1000), .A3(new_n1097), .A4(new_n1094), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1093), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(new_n1099), .B(KEYINPUT119), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1091), .B1(new_n1100), .B2(new_n554), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1093), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(KEYINPUT119), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1099), .A2(new_n1106), .ZN(new_n1107));
  AND4_X1   g682(.A1(new_n1091), .A2(new_n1105), .A3(new_n554), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g683(.A(KEYINPUT59), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1100), .A2(new_n1091), .A3(new_n554), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1105), .A2(new_n554), .A3(new_n1107), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT120), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1110), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1090), .B1(new_n1109), .B2(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1078), .A2(new_n1086), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1116), .A2(new_n1077), .ZN(new_n1117));
  XNOR2_X1  g692(.A(new_n1117), .B(KEYINPUT116), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1069), .B1(new_n1115), .B2(new_n1118), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n990), .A2(G168), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1017), .A2(new_n1040), .A3(new_n1120), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT114), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT63), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT114), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1017), .A2(new_n1040), .A3(new_n1120), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1122), .A2(new_n1123), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(new_n1036), .ZN(new_n1127));
  AND3_X1   g702(.A1(new_n1017), .A2(KEYINPUT63), .A3(new_n1127), .ZN(new_n1128));
  AND2_X1   g703(.A1(new_n1008), .A2(G8), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1128), .B(new_n1120), .C1(new_n1015), .C2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1126), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(G1976), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1029), .A2(new_n1132), .A3(new_n716), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1133), .A2(KEYINPUT111), .A3(new_n1022), .ZN(new_n1134));
  NOR2_X1   g709(.A1(new_n1083), .A2(new_n989), .ZN(new_n1135));
  OR2_X1    g710(.A1(new_n1135), .A2(KEYINPUT110), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1135), .A2(KEYINPUT110), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1133), .A2(new_n1022), .ZN(new_n1139));
  OAI211_X1 g714(.A(new_n1137), .B(new_n1138), .C1(KEYINPUT111), .C2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1140), .B1(new_n1036), .B2(new_n1017), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT112), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT112), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1140), .B(new_n1143), .C1(new_n1036), .C2(new_n1017), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1131), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT115), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n996), .A2(new_n997), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT62), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1065), .A2(new_n1062), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n996), .A2(KEYINPUT62), .A3(new_n997), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1151), .A2(new_n1152), .A3(new_n1041), .A4(new_n1153), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1131), .A2(new_n1145), .A3(KEYINPUT115), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1119), .A2(new_n1148), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1048), .A2(new_n978), .ZN(new_n1157));
  NOR2_X1   g732(.A1(new_n1157), .A2(new_n999), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1158), .A2(G1996), .A3(new_n848), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT104), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n813), .B(new_n1082), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1161), .B1(G1996), .B2(new_n848), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1160), .B1(new_n1158), .B2(new_n1162), .ZN(new_n1163));
  AND2_X1   g738(.A1(new_n700), .A2(new_n702), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n700), .A2(new_n702), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1158), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(G1986), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n692), .A2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1169), .A2(KEYINPUT103), .ZN(new_n1170));
  NAND2_X1  g745(.A1(G290), .A2(G1986), .ZN(new_n1171));
  MUX2_X1   g746(.A(KEYINPUT103), .B(new_n1170), .S(new_n1171), .Z(new_n1172));
  AOI21_X1  g747(.A(new_n1167), .B1(new_n1158), .B2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1156), .A2(new_n1173), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n814), .A2(new_n1082), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(KEYINPUT126), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT126), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1175), .A2(new_n1179), .A3(new_n1176), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1178), .A2(new_n1158), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1158), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT46), .ZN(new_n1183));
  OR3_X1    g758(.A1(new_n1182), .A2(new_n1183), .A3(G1996), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1161), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1158), .B1(new_n1185), .B2(new_n848), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1183), .B1(new_n1182), .B2(G1996), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1184), .A2(new_n1186), .A3(new_n1187), .ZN(new_n1188));
  XNOR2_X1  g763(.A(new_n1188), .B(KEYINPUT47), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1182), .A2(new_n1169), .ZN(new_n1190));
  XOR2_X1   g765(.A(new_n1190), .B(KEYINPUT48), .Z(new_n1191));
  NAND3_X1  g766(.A1(new_n1163), .A2(new_n1166), .A3(new_n1191), .ZN(new_n1192));
  AND3_X1   g767(.A1(new_n1181), .A2(new_n1189), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1174), .A2(new_n1193), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g769(.A(G401), .ZN(new_n1196));
  NOR2_X1   g770(.A1(G229), .A2(new_n461), .ZN(new_n1197));
  NAND4_X1  g771(.A1(new_n904), .A2(new_n1196), .A3(new_n667), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g772(.A(new_n950), .ZN(new_n1199));
  NAND3_X1  g773(.A1(new_n967), .A2(new_n885), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g774(.A1(new_n1200), .A2(KEYINPUT43), .ZN(new_n1201));
  AOI211_X1 g775(.A(KEYINPUT127), .B(new_n1198), .C1(new_n1201), .C2(new_n969), .ZN(new_n1202));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n1203));
  INV_X1    g777(.A(new_n1198), .ZN(new_n1204));
  AOI21_X1  g778(.A(new_n1203), .B1(new_n970), .B2(new_n1204), .ZN(new_n1205));
  NOR2_X1   g779(.A1(new_n1202), .A2(new_n1205), .ZN(G308));
  INV_X1    g780(.A(new_n969), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n968), .B1(new_n957), .B2(new_n1199), .ZN(new_n1208));
  OAI21_X1  g782(.A(new_n1204), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1209));
  NAND2_X1  g783(.A1(new_n1209), .A2(KEYINPUT127), .ZN(new_n1210));
  NAND3_X1  g784(.A1(new_n970), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1211));
  NAND2_X1  g785(.A1(new_n1210), .A2(new_n1211), .ZN(G225));
endmodule


