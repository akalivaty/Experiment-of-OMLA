//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 0 1 1 0 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n251, new_n252,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n259, new_n260,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1267, new_n1268, new_n1269,
    new_n1270;
  OR3_X1    g0000(.A1(KEYINPUT64), .A2(G58), .A3(G68), .ZN(new_n201));
  OAI21_X1  g0001(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g0003(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G50), .ZN(new_n205));
  INV_X1    g0005(.A(G77), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(G353));
  OAI21_X1  g0008(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0009(.A(G250), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(G257), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n210), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n204), .A2(G50), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n222), .A2(G20), .ZN(new_n223));
  OAI22_X1  g0023(.A1(new_n219), .A2(KEYINPUT0), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT0), .B2(new_n219), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT66), .Z(new_n226));
  INV_X1    g0026(.A(G87), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  OAI22_X1  g0028(.A1(new_n227), .A2(new_n210), .B1(new_n228), .B2(new_n217), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(G68), .B2(G238), .ZN(new_n230));
  INV_X1    g0030(.A(G107), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n230), .B1(new_n231), .B2(new_n218), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(G116), .B2(G270), .ZN(new_n233));
  INV_X1    g0033(.A(G50), .ZN(new_n234));
  INV_X1    g0034(.A(G226), .ZN(new_n235));
  INV_X1    g0035(.A(G244), .ZN(new_n236));
  OAI221_X1 g0036(.A(new_n233), .B1(new_n234), .B2(new_n235), .C1(new_n206), .C2(new_n236), .ZN(new_n237));
  INV_X1    g0037(.A(G58), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  NOR2_X1   g0039(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g0040(.A(new_n214), .B1(new_n237), .B2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT1), .ZN(new_n242));
  NOR2_X1   g0042(.A1(new_n226), .A2(new_n242), .ZN(G361));
  XOR2_X1   g0043(.A(G250), .B(G257), .Z(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT67), .B(KEYINPUT68), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT2), .B(G226), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n239), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G238), .B(G244), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n248), .B(new_n252), .Z(G358));
  XNOR2_X1  g0053(.A(G68), .B(G77), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT69), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n255), .B(new_n234), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n256), .B(G58), .ZN(new_n257));
  XNOR2_X1  g0057(.A(G87), .B(G116), .ZN(new_n258));
  XNOR2_X1  g0058(.A(G97), .B(G107), .ZN(new_n259));
  XNOR2_X1  g0059(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g0060(.A(new_n257), .B(new_n260), .ZN(G351));
  INV_X1    g0061(.A(KEYINPUT3), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT70), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n263), .A2(new_n265), .A3(KEYINPUT70), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n271), .A2(new_n206), .ZN(new_n272));
  AND2_X1   g0072(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n273));
  NOR2_X1   g0073(.A1(KEYINPUT71), .A2(G1698), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G222), .ZN(new_n276));
  INV_X1    g0076(.A(G223), .ZN(new_n277));
  INV_X1    g0077(.A(G1698), .ZN(new_n278));
  OAI22_X1  g0078(.A1(new_n275), .A2(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n272), .B1(new_n271), .B2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT72), .ZN(new_n281));
  OR2_X1    g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n222), .B1(new_n264), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n280), .A2(new_n281), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n282), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n288));
  INV_X1    g0088(.A(G274), .ZN(new_n289));
  OR2_X1    g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n288), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n287), .B(new_n290), .C1(new_n235), .C2(new_n291), .ZN(new_n292));
  OR2_X1    g0092(.A1(new_n292), .A2(G179), .ZN(new_n293));
  OR2_X1    g0093(.A1(KEYINPUT8), .A2(G58), .ZN(new_n294));
  NAND2_X1  g0094(.A1(KEYINPUT8), .A2(G58), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  NOR2_X1   g0097(.A1(new_n264), .A2(G20), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  AOI22_X1  g0099(.A1(new_n297), .A2(new_n298), .B1(G150), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g0100(.A(new_n300), .B1(new_n205), .B2(new_n212), .ZN(new_n301));
  NAND3_X1  g0101(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(new_n221), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT73), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n301), .A2(new_n304), .B1(new_n234), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n304), .A2(new_n306), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n211), .A2(G20), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(G50), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n292), .A2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n293), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n292), .A2(G200), .ZN(new_n316));
  XNOR2_X1  g0116(.A(new_n311), .B(KEYINPUT9), .ZN(new_n317));
  INV_X1    g0117(.A(G190), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n292), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n322), .ZN(new_n323));
  INV_X1    g0123(.A(G238), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n275), .A2(new_n235), .B1(new_n239), .B2(new_n278), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n270), .A2(new_n325), .B1(G33), .B2(G97), .ZN(new_n326));
  OAI221_X1 g0126(.A(new_n290), .B1(new_n324), .B2(new_n291), .C1(new_n326), .C2(new_n284), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(KEYINPUT13), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(G200), .ZN(new_n331));
  INV_X1    g0131(.A(G68), .ZN(new_n332));
  AOI22_X1  g0132(.A1(new_n298), .A2(G77), .B1(G20), .B2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n299), .ZN(new_n334));
  OAI21_X1  g0134(.A(new_n333), .B1(new_n234), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n304), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT11), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT75), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n305), .B(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(KEYINPUT12), .A3(new_n332), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n306), .A2(KEYINPUT12), .ZN(new_n342));
  INV_X1    g0142(.A(new_n303), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n339), .A2(new_n343), .A3(new_n309), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT12), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n342), .B1(new_n345), .B2(G68), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n337), .A2(new_n341), .A3(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT77), .ZN(new_n348));
  XNOR2_X1  g0148(.A(new_n347), .B(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n328), .A2(G190), .A3(new_n329), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n331), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT78), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT17), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT80), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n355), .B1(new_n262), .B2(G33), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT79), .B(G33), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n356), .B1(new_n357), .B2(new_n262), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT79), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G33), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n264), .A2(KEYINPUT79), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n355), .B(KEYINPUT3), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n275), .A2(new_n277), .B1(new_n235), .B2(new_n278), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n363), .A2(new_n364), .B1(G33), .B2(G87), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n365), .A2(new_n284), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n290), .B1(new_n291), .B2(new_n239), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(G190), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n297), .A2(new_n309), .ZN(new_n370));
  XOR2_X1   g0170(.A(new_n370), .B(KEYINPUT83), .Z(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n308), .B1(new_n306), .B2(new_n296), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT16), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n238), .A2(new_n332), .ZN(new_n374));
  OAI21_X1  g0174(.A(G20), .B1(new_n203), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n299), .A2(G159), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n358), .A2(new_n212), .A3(new_n362), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT81), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n378), .A2(KEYINPUT81), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n263), .A2(KEYINPUT80), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n264), .A2(KEYINPUT79), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n359), .A2(G33), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n384), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n388));
  AOI211_X1 g0188(.A(KEYINPUT80), .B(new_n262), .C1(new_n385), .C2(new_n386), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT82), .ZN(new_n391));
  NAND4_X1  g0191(.A1(new_n390), .A2(new_n391), .A3(KEYINPUT7), .A4(new_n212), .ZN(new_n392));
  OAI21_X1  g0192(.A(KEYINPUT82), .B1(new_n378), .B2(new_n379), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n382), .A2(new_n383), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  AOI211_X1 g0194(.A(new_n373), .B(new_n377), .C1(new_n394), .C2(G68), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n379), .B1(new_n270), .B2(G20), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n265), .B1(new_n387), .B2(KEYINPUT3), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(KEYINPUT7), .A3(new_n212), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n377), .B1(new_n399), .B2(G68), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n303), .B1(new_n400), .B2(KEYINPUT16), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n369), .B(new_n372), .C1(new_n395), .C2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(G200), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n368), .A2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n354), .B1(new_n402), .B2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n372), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n377), .B1(new_n394), .B2(G68), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT16), .ZN(new_n408));
  INV_X1    g0208(.A(new_n401), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n406), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(new_n404), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n410), .A2(KEYINPUT17), .A3(new_n411), .A4(new_n369), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n372), .B1(new_n395), .B2(new_n401), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n368), .A2(G179), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n312), .B2(new_n368), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(KEYINPUT18), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT18), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n405), .B(new_n412), .C1(new_n416), .C2(new_n417), .ZN(new_n418));
  OAI22_X1  g0218(.A1(new_n275), .A2(new_n239), .B1(new_n324), .B2(new_n278), .ZN(new_n419));
  NOR2_X1   g0219(.A1(new_n271), .A2(new_n419), .ZN(new_n420));
  XOR2_X1   g0220(.A(KEYINPUT74), .B(G107), .Z(new_n421));
  INV_X1    g0221(.A(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n285), .B1(new_n270), .B2(new_n422), .ZN(new_n423));
  OAI221_X1 g0223(.A(new_n290), .B1(new_n236), .B2(new_n291), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(new_n312), .ZN(new_n425));
  XOR2_X1   g0225(.A(KEYINPUT15), .B(G87), .Z(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n298), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n296), .A2(new_n334), .B1(new_n212), .B2(new_n206), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n303), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n340), .A2(new_n206), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n431), .B(new_n432), .C1(new_n206), .C2(new_n344), .ZN(new_n433));
  OAI211_X1 g0233(.A(new_n425), .B(new_n433), .C1(G179), .C2(new_n424), .ZN(new_n434));
  INV_X1    g0234(.A(new_n434), .ZN(new_n435));
  OR3_X1    g0235(.A1(new_n353), .A2(new_n418), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(KEYINPUT14), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n437), .B1(new_n330), .B2(G169), .ZN(new_n438));
  AOI211_X1 g0238(.A(KEYINPUT14), .B(new_n312), .C1(new_n328), .C2(new_n329), .ZN(new_n439));
  INV_X1    g0239(.A(G179), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n330), .A2(new_n440), .ZN(new_n441));
  NOR3_X1   g0241(.A1(new_n438), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n349), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n433), .B1(new_n424), .B2(G200), .ZN(new_n447));
  XNOR2_X1  g0247(.A(new_n447), .B(KEYINPUT76), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n424), .A2(new_n318), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NOR4_X1   g0251(.A1(new_n323), .A2(new_n436), .A3(new_n446), .A4(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT23), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n421), .B2(G20), .ZN(new_n455));
  INV_X1    g0255(.A(G116), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n387), .A2(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n212), .B2(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n454), .A2(new_n231), .A3(G20), .ZN(new_n459));
  XNOR2_X1  g0259(.A(new_n459), .B(KEYINPUT93), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT91), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n212), .A2(G87), .ZN(new_n462));
  INV_X1    g0262(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n363), .B2(new_n463), .ZN(new_n464));
  AOI211_X1 g0264(.A(KEYINPUT91), .B(new_n462), .C1(new_n358), .C2(new_n362), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT22), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n271), .A2(KEYINPUT22), .A3(new_n462), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n458), .B(new_n460), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT92), .B(KEYINPUT24), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g0271(.A(KEYINPUT91), .B1(new_n390), .B2(new_n462), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n363), .A2(new_n461), .A3(new_n463), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n472), .A2(KEYINPUT22), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n468), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(new_n470), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n458), .A4(new_n460), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n471), .A2(new_n303), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT94), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT94), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n471), .A2(new_n481), .A3(new_n303), .A4(new_n478), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n306), .A2(new_n231), .ZN(new_n484));
  XNOR2_X1  g0284(.A(new_n484), .B(KEYINPUT25), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n308), .B1(G1), .B2(new_n264), .ZN(new_n486));
  INV_X1    g0286(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(G107), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n483), .A2(new_n488), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n275), .A2(new_n210), .B1(new_n217), .B2(new_n278), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n363), .A2(new_n490), .B1(G294), .B2(new_n357), .ZN(new_n491));
  OR2_X1    g0291(.A1(new_n491), .A2(new_n284), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT5), .ZN(new_n493));
  OR3_X1    g0293(.A1(new_n493), .A2(KEYINPUT85), .A3(G41), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n493), .B1(KEYINPUT85), .B2(G41), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n211), .A2(G45), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  AND2_X1   g0297(.A1(new_n497), .A2(new_n284), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(G264), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n492), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n497), .A2(new_n289), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n312), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(G179), .B2(new_n503), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n489), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n456), .B1(new_n211), .B2(G33), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n339), .A2(new_n343), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n303), .B1(new_n212), .B2(G116), .ZN(new_n510));
  XNOR2_X1  g0310(.A(new_n510), .B(KEYINPUT89), .ZN(new_n511));
  NAND2_X1  g0311(.A1(G33), .A2(G283), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n212), .C1(G33), .C2(new_n228), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(KEYINPUT20), .A3(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(KEYINPUT20), .B1(new_n511), .B2(new_n513), .ZN(new_n516));
  OAI221_X1 g0316(.A(new_n509), .B1(G116), .B2(new_n339), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n273), .A2(new_n274), .ZN(new_n518));
  AOI22_X1  g0318(.A1(new_n518), .A2(G257), .B1(G264), .B2(G1698), .ZN(new_n519));
  INV_X1    g0319(.A(G303), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n390), .A2(new_n519), .B1(new_n520), .B2(new_n270), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n285), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n501), .B1(new_n498), .B2(G270), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n517), .A2(G169), .A3(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT90), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT21), .ZN(new_n528));
  INV_X1    g0328(.A(new_n524), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n517), .A2(G179), .A3(new_n529), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT21), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n524), .A2(new_n318), .ZN(new_n534));
  AOI211_X1 g0334(.A(new_n534), .B(new_n517), .C1(G200), .C2(new_n524), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n518), .A2(KEYINPUT4), .A3(G244), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n537), .B1(new_n210), .B2(new_n278), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(new_n270), .ZN(new_n539));
  AOI211_X1 g0339(.A(new_n236), .B(new_n275), .C1(new_n358), .C2(new_n362), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n539), .B(new_n512), .C1(new_n540), .C2(KEYINPUT4), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n285), .ZN(new_n542));
  INV_X1    g0342(.A(new_n501), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n498), .A2(G257), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n228), .A2(new_n231), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n231), .A2(KEYINPUT6), .A3(G97), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI22_X1  g0352(.A1(new_n552), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n553));
  XNOR2_X1  g0353(.A(new_n553), .B(KEYINPUT84), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n399), .A2(new_n422), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n343), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n305), .A2(G97), .ZN(new_n557));
  INV_X1    g0357(.A(new_n557), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n558), .B1(new_n486), .B2(new_n228), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n546), .B(new_n560), .C1(new_n318), .C2(new_n545), .ZN(new_n561));
  INV_X1    g0361(.A(new_n559), .ZN(new_n562));
  AND2_X1   g0362(.A1(new_n554), .A2(new_n555), .ZN(new_n563));
  OAI211_X1 g0363(.A(KEYINPUT86), .B(new_n562), .C1(new_n563), .C2(new_n343), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n556), .B2(new_n559), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n542), .A2(G179), .A3(new_n543), .A4(new_n544), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n541), .A2(new_n285), .B1(G257), .B2(new_n498), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n312), .B1(new_n569), .B2(new_n543), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n564), .B(new_n566), .C1(new_n568), .C2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n363), .A2(new_n212), .A3(G68), .ZN(new_n572));
  XNOR2_X1  g0372(.A(KEYINPUT87), .B(G87), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n421), .A2(new_n573), .A3(new_n228), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT19), .ZN(new_n575));
  NOR3_X1   g0375(.A1(new_n575), .A2(new_n264), .A3(new_n228), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n574), .B1(G20), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n575), .B1(new_n428), .B2(new_n228), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n572), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n303), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT88), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n340), .A2(new_n427), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n581), .B1(new_n580), .B2(new_n582), .ZN(new_n584));
  OR2_X1    g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  OAI22_X1  g0385(.A1(new_n275), .A2(new_n324), .B1(new_n236), .B2(new_n278), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n457), .B1(new_n363), .B2(new_n586), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n587), .A2(new_n284), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n496), .A2(new_n289), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n589), .B(new_n284), .C1(G250), .C2(new_n496), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G190), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n487), .A2(G87), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(G200), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n585), .A2(new_n593), .A3(new_n594), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n487), .A2(new_n426), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n583), .B2(new_n584), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n592), .A2(new_n440), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n598), .B(new_n599), .C1(G169), .C2(new_n592), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n561), .A2(new_n571), .A3(new_n596), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n503), .A2(G200), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n502), .A2(G190), .ZN(new_n603));
  NAND4_X1  g0403(.A1(new_n483), .A2(new_n488), .A3(new_n602), .A4(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n507), .A2(new_n536), .A3(new_n601), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n453), .A2(new_n605), .ZN(G372));
  AOI21_X1  g0406(.A(new_n505), .B1(new_n483), .B2(new_n488), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n601), .B(new_n604), .C1(new_n607), .C2(new_n533), .ZN(new_n608));
  INV_X1    g0408(.A(new_n600), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n545), .A2(G169), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n560), .B1(new_n610), .B2(new_n567), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n596), .A2(new_n600), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n571), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n596), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n609), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n608), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n452), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g0419(.A(new_n619), .B(KEYINPUT95), .Z(new_n620));
  OR2_X1    g0420(.A1(new_n416), .A2(new_n417), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n446), .B1(new_n351), .B2(new_n435), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n405), .A2(new_n412), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n320), .A2(new_n321), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n315), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n620), .A2(new_n626), .ZN(G369));
  AND4_X1   g0427(.A1(new_n483), .A2(new_n488), .A3(new_n602), .A4(new_n603), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n211), .A2(new_n212), .A3(G13), .ZN(new_n629));
  OR2_X1    g0429(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(KEYINPUT27), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n630), .A2(G213), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(KEYINPUT96), .B(G343), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n483), .B2(new_n488), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n628), .A2(new_n607), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n607), .A2(new_n635), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT97), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n489), .A2(new_n635), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n507), .A2(new_n642), .A3(new_n604), .ZN(new_n643));
  INV_X1    g0443(.A(KEYINPUT97), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(new_n644), .A3(new_n639), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n641), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n517), .A2(new_n635), .ZN(new_n648));
  OR3_X1    g0448(.A1(new_n533), .A2(new_n535), .A3(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n533), .A2(new_n648), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(G330), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n647), .A2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n507), .A2(new_n635), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n533), .A2(new_n636), .ZN(new_n659));
  XNOR2_X1  g0459(.A(new_n659), .B(KEYINPUT98), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n646), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n657), .A2(new_n661), .ZN(G399));
  NOR2_X1   g0462(.A1(new_n216), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G1), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n574), .A2(G116), .ZN(new_n666));
  OAI22_X1  g0466(.A1(new_n665), .A2(new_n666), .B1(new_n220), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  NOR4_X1   g0468(.A1(new_n567), .A2(new_n524), .A3(new_n591), .A4(new_n500), .ZN(new_n669));
  OAI21_X1  g0469(.A(KEYINPUT30), .B1(new_n669), .B2(KEYINPUT99), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT99), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT30), .ZN(new_n672));
  AND3_X1   g0472(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n673), .A2(G179), .A3(new_n529), .A4(new_n592), .ZN(new_n674));
  OAI211_X1 g0474(.A(new_n671), .B(new_n672), .C1(new_n674), .C2(new_n500), .ZN(new_n675));
  NOR3_X1   g0475(.A1(new_n673), .A2(new_n529), .A3(new_n502), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n676), .A2(new_n440), .A3(new_n591), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n670), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n678), .A2(KEYINPUT31), .A3(new_n635), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(new_n635), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT31), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n679), .B(new_n682), .C1(new_n605), .C2(new_n635), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n635), .B1(new_n608), .B2(new_n617), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT29), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n561), .B(new_n604), .C1(new_n607), .C2(new_n533), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n571), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n596), .A2(new_n600), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n615), .ZN(new_n692));
  NAND3_X1  g0492(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n600), .B(KEYINPUT100), .Z(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(KEYINPUT26), .B2(new_n612), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n635), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n684), .B(new_n687), .C1(new_n696), .C2(new_n686), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n668), .B1(new_n698), .B2(G1), .ZN(G364));
  NAND3_X1  g0499(.A1(new_n212), .A2(G13), .A3(G45), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n664), .A2(G1), .A3(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(G13), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(new_n264), .A3(KEYINPUT103), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT103), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n704), .B1(G13), .B2(G33), .ZN(new_n705));
  AOI21_X1  g0505(.A(G20), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n652), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n221), .B1(G20), .B2(new_n312), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n212), .A2(G179), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n403), .A2(G190), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n318), .A2(new_n403), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n710), .ZN(new_n714));
  OAI221_X1 g0514(.A(new_n270), .B1(new_n231), .B2(new_n712), .C1(new_n573), .C2(new_n714), .ZN(new_n715));
  XOR2_X1   g0515(.A(new_n715), .B(KEYINPUT104), .Z(new_n716));
  NOR2_X1   g0516(.A1(G190), .A2(G200), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n710), .A2(new_n717), .ZN(new_n718));
  INV_X1    g0518(.A(G159), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT32), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n318), .A2(G179), .A3(G200), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(new_n212), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n720), .A2(new_n721), .B1(new_n228), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n212), .A2(new_n440), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(new_n713), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n711), .ZN(new_n727));
  OAI22_X1  g0527(.A1(new_n726), .A2(new_n234), .B1(new_n727), .B2(new_n332), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n716), .A2(new_n724), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n717), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G77), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n720), .A2(new_n721), .ZN(new_n733));
  INV_X1    g0533(.A(new_n725), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n734), .A2(new_n318), .A3(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G58), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n729), .A2(new_n732), .A3(new_n733), .A4(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G311), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n271), .B1(new_n738), .B2(new_n730), .ZN(new_n739));
  INV_X1    g0539(.A(new_n712), .ZN(new_n740));
  INV_X1    g0540(.A(new_n718), .ZN(new_n741));
  AOI22_X1  g0541(.A1(G283), .A2(new_n740), .B1(new_n741), .B2(G329), .ZN(new_n742));
  INV_X1    g0542(.A(G294), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  INV_X1    g0544(.A(new_n735), .ZN(new_n745));
  OAI221_X1 g0545(.A(new_n742), .B1(new_n743), .B2(new_n723), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n727), .ZN(new_n747));
  XNOR2_X1  g0547(.A(KEYINPUT105), .B(KEYINPUT33), .ZN(new_n748));
  INV_X1    g0548(.A(G317), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n748), .B(new_n749), .ZN(new_n750));
  AOI211_X1 g0550(.A(new_n739), .B(new_n746), .C1(new_n747), .C2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G326), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n751), .B1(new_n520), .B2(new_n714), .C1(new_n752), .C2(new_n726), .ZN(new_n753));
  AND2_X1   g0553(.A1(new_n737), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n257), .A2(G45), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT101), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n363), .A2(new_n216), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(G45), .B2(new_n220), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n758), .B1(G116), .B2(new_n215), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n271), .A2(new_n216), .ZN(new_n760));
  AOI21_X1  g0560(.A(new_n759), .B1(G355), .B2(new_n760), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT102), .Z(new_n762));
  NOR2_X1   g0562(.A1(new_n706), .A2(new_n708), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI221_X1 g0564(.A(new_n707), .B1(new_n709), .B2(new_n754), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n652), .A2(new_n653), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n655), .A2(new_n701), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n765), .A2(new_n767), .ZN(G396));
  NAND2_X1  g0568(.A1(new_n435), .A2(new_n636), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n448), .A2(new_n449), .B1(new_n433), .B2(new_n635), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n769), .B1(new_n770), .B2(new_n435), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n685), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g0573(.A(new_n635), .B(new_n771), .C1(new_n608), .C2(new_n617), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(new_n684), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(new_n701), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n703), .A2(new_n705), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n771), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n701), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(new_n708), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n206), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n735), .A2(G143), .B1(G159), .B2(new_n731), .ZN(new_n783));
  INV_X1    g0583(.A(G137), .ZN(new_n784));
  INV_X1    g0584(.A(G150), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n783), .B1(new_n784), .B2(new_n726), .C1(new_n785), .C2(new_n727), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT34), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n390), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n788), .B1(new_n238), .B2(new_n723), .ZN(new_n789));
  INV_X1    g0589(.A(G132), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n718), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n712), .A2(new_n332), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n786), .A2(new_n787), .B1(new_n234), .B2(new_n714), .ZN(new_n793));
  NOR4_X1   g0593(.A1(new_n789), .A2(new_n791), .A3(new_n792), .A4(new_n793), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n712), .A2(new_n227), .B1(new_n718), .B2(new_n738), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT106), .ZN(new_n796));
  OAI221_X1 g0596(.A(new_n796), .B1(new_n228), .B2(new_n723), .C1(new_n456), .C2(new_n730), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n714), .A2(new_n231), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n745), .A2(new_n743), .ZN(new_n799));
  INV_X1    g0599(.A(G283), .ZN(new_n800));
  OAI221_X1 g0600(.A(new_n271), .B1(new_n800), .B2(new_n727), .C1(new_n520), .C2(new_n726), .ZN(new_n801));
  NOR4_X1   g0601(.A1(new_n797), .A2(new_n798), .A3(new_n799), .A4(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n708), .B1(new_n794), .B2(new_n802), .ZN(new_n803));
  NAND4_X1  g0603(.A1(new_n779), .A2(new_n780), .A3(new_n782), .A4(new_n803), .ZN(new_n804));
  AND2_X1   g0604(.A1(new_n777), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(G384));
  OAI211_X1 g0606(.A(G20), .B(new_n222), .C1(new_n552), .C2(KEYINPUT35), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n456), .B(new_n807), .C1(KEYINPUT35), .C2(new_n552), .ZN(new_n808));
  XOR2_X1   g0608(.A(new_n808), .B(KEYINPUT36), .Z(new_n809));
  OAI21_X1  g0609(.A(G77), .B1(new_n238), .B2(new_n332), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n220), .A2(new_n810), .B1(G50), .B2(new_n332), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n811), .A2(G1), .A3(new_n702), .ZN(new_n812));
  INV_X1    g0612(.A(KEYINPUT40), .ZN(new_n813));
  INV_X1    g0613(.A(new_n632), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n407), .A2(KEYINPUT16), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n815), .A2(new_n304), .A3(new_n408), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n816), .A2(new_n372), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n418), .A2(new_n814), .A3(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n415), .A2(new_n814), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n816), .B2(new_n372), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n402), .A2(new_n404), .ZN(new_n821));
  OAI21_X1  g0621(.A(KEYINPUT37), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(KEYINPUT37), .ZN(new_n823));
  OAI221_X1 g0623(.A(new_n823), .B1(new_n402), .B2(new_n404), .C1(new_n410), .C2(new_n819), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n818), .A2(new_n825), .A3(KEYINPUT38), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT38), .B1(new_n818), .B2(new_n825), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT107), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n818), .A2(new_n825), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT38), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT107), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n818), .A2(new_n825), .A3(KEYINPUT38), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n349), .A2(new_n636), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n353), .B2(new_n443), .ZN(new_n837));
  INV_X1    g0637(.A(new_n836), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n445), .A2(new_n351), .A3(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n771), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n683), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n813), .B1(new_n835), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n840), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n410), .A2(new_n819), .ZN(new_n844));
  OAI21_X1  g0644(.A(KEYINPUT37), .B1(new_n844), .B2(new_n821), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n824), .A3(KEYINPUT108), .ZN(new_n846));
  INV_X1    g0646(.A(KEYINPUT108), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n847), .B(KEYINPUT37), .C1(new_n844), .C2(new_n821), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n418), .A2(new_n413), .A3(new_n814), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n830), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n833), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(KEYINPUT109), .B1(new_n683), .B2(new_n840), .ZN(new_n854));
  NOR4_X1   g0654(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT110), .A4(new_n813), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT110), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n843), .A2(new_n852), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT109), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n813), .B1(new_n841), .B2(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n856), .B1(new_n857), .B2(new_n859), .ZN(new_n860));
  OAI211_X1 g0660(.A(G330), .B(new_n842), .C1(new_n855), .C2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n452), .A2(G330), .A3(new_n683), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n863), .B(KEYINPUT111), .ZN(new_n864));
  AND2_X1   g0664(.A1(new_n828), .A2(new_n834), .ZN(new_n865));
  INV_X1    g0665(.A(new_n841), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT40), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n841), .A2(new_n858), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n868), .A2(KEYINPUT40), .A3(new_n843), .A4(new_n852), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(KEYINPUT110), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n857), .A2(new_n856), .A3(new_n859), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n867), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n872), .A2(new_n452), .A3(new_n683), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n864), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n621), .A2(new_n814), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n837), .A2(new_n839), .ZN(new_n877));
  INV_X1    g0677(.A(new_n769), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n877), .B1(new_n774), .B2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n835), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(KEYINPUT39), .B1(new_n851), .B2(new_n833), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT39), .ZN(new_n882));
  NOR3_X1   g0682(.A1(new_n826), .A2(new_n827), .A3(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n445), .A2(new_n635), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n881), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n880), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(new_n626), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n687), .B1(new_n696), .B2(new_n686), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n888), .B1(new_n889), .B2(new_n452), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n887), .B(new_n890), .Z(new_n891));
  XOR2_X1   g0691(.A(new_n874), .B(new_n891), .Z(new_n892));
  AOI21_X1  g0692(.A(new_n211), .B1(G13), .B2(new_n212), .ZN(new_n893));
  OAI211_X1 g0693(.A(new_n809), .B(new_n812), .C1(new_n892), .C2(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT112), .Z(G367));
  OR2_X1    g0695(.A1(new_n571), .A2(new_n635), .ZN(new_n896));
  AND3_X1   g0696(.A1(new_n643), .A2(new_n644), .A3(new_n639), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n644), .B1(new_n643), .B2(new_n639), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n660), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  OAI211_X1 g0699(.A(new_n571), .B(new_n561), .C1(new_n560), .C2(new_n636), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n611), .A2(new_n635), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g0702(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g0703(.A(KEYINPUT42), .B1(new_n899), .B2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n660), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n905), .B1(new_n641), .B2(new_n645), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT42), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n658), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OAI211_X1 g0708(.A(new_n896), .B(new_n904), .C1(new_n908), .C2(new_n903), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n656), .A2(new_n902), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n585), .A2(new_n594), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n911), .A2(new_n635), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n691), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n609), .A2(new_n911), .A3(new_n635), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n909), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n910), .B1(new_n909), .B2(new_n916), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n909), .A2(new_n916), .ZN(new_n923));
  INV_X1    g0723(.A(new_n910), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g0725(.A(new_n920), .B1(new_n925), .B2(new_n917), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  XNOR2_X1  g0727(.A(new_n663), .B(KEYINPUT41), .ZN(new_n928));
  INV_X1    g0728(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(KEYINPUT44), .B1(new_n661), .B2(new_n902), .ZN(new_n930));
  INV_X1    g0730(.A(new_n658), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n899), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT44), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n932), .A2(new_n933), .A3(new_n903), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT45), .B1(new_n661), .B2(new_n902), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT45), .ZN(new_n936));
  NOR4_X1   g0736(.A1(new_n906), .A2(new_n936), .A3(new_n658), .A4(new_n903), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n930), .B(new_n934), .C1(new_n935), .C2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(new_n656), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n933), .B1(new_n932), .B2(new_n903), .ZN(new_n940));
  AOI211_X1 g0740(.A(KEYINPUT44), .B(new_n902), .C1(new_n899), .C2(new_n931), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n936), .B1(new_n932), .B2(new_n903), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n661), .A2(KEYINPUT45), .A3(new_n902), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n942), .A2(new_n657), .A3(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n641), .A2(new_n645), .A3(new_n905), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n899), .A2(new_n654), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n654), .B1(new_n899), .B2(new_n947), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n698), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n939), .A2(new_n946), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n929), .B1(new_n953), .B2(new_n698), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n700), .A2(G1), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT113), .Z(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n927), .B1(new_n954), .B2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n757), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n248), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n763), .B1(new_n215), .B2(new_n427), .ZN(new_n961));
  INV_X1    g0761(.A(G143), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n726), .A2(new_n962), .B1(new_n727), .B2(new_n719), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n723), .A2(new_n332), .ZN(new_n964));
  NOR2_X1   g0764(.A1(new_n730), .A2(new_n234), .ZN(new_n965));
  OR3_X1    g0765(.A1(new_n963), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n745), .A2(new_n785), .B1(new_n712), .B2(new_n206), .ZN(new_n967));
  NOR3_X1   g0767(.A1(new_n966), .A2(new_n967), .A3(new_n271), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n968), .B1(new_n238), .B2(new_n714), .C1(new_n784), .C2(new_n718), .ZN(new_n969));
  XOR2_X1   g0769(.A(KEYINPUT114), .B(G311), .Z(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n390), .B1(new_n726), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n714), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n973), .A2(KEYINPUT46), .A3(G116), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n975), .B1(new_n714), .B2(new_n456), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n974), .B(new_n976), .C1(new_n743), .C2(new_n727), .ZN(new_n977));
  INV_X1    g0777(.A(KEYINPUT115), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n972), .B(new_n979), .C1(G317), .C2(new_n741), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n731), .A2(G283), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n735), .A2(G303), .ZN(new_n982));
  INV_X1    g0782(.A(new_n723), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n977), .A2(new_n978), .B1(new_n422), .B2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n712), .A2(new_n228), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n969), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT47), .Z(new_n988));
  OAI221_X1 g0788(.A(new_n780), .B1(new_n960), .B2(new_n961), .C1(new_n988), .C2(new_n709), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT116), .Z(new_n990));
  INV_X1    g0790(.A(new_n706), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n990), .B1(new_n991), .B2(new_n915), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n958), .A2(new_n992), .ZN(G387));
  OAI21_X1  g0793(.A(new_n697), .B1(new_n948), .B2(new_n949), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n951), .A2(new_n663), .A3(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n714), .A2(new_n206), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n983), .A2(new_n426), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n719), .B2(new_n726), .C1(new_n745), .C2(new_n234), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n998), .C1(new_n297), .C2(new_n747), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n731), .A2(G68), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n986), .B1(G150), .B2(new_n741), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n999), .A2(new_n363), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n726), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G322), .A2(new_n1003), .B1(new_n731), .B2(G303), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n727), .B2(new_n971), .C1(new_n749), .C2(new_n745), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT48), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n800), .B2(new_n723), .C1(new_n743), .C2(new_n714), .ZN(new_n1007));
  XOR2_X1   g0807(.A(new_n1007), .B(KEYINPUT49), .Z(new_n1008));
  OAI221_X1 g0808(.A(new_n390), .B1(new_n456), .B2(new_n712), .C1(new_n752), .C2(new_n718), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT117), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1002), .B1(new_n1008), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1011), .A2(new_n708), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n959), .B1(new_n252), .B2(G45), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1013), .B1(new_n666), .B2(new_n760), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n297), .A2(new_n234), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT50), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n332), .A2(new_n206), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1016), .A2(new_n666), .A3(G45), .A4(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1014), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n231), .B2(new_n216), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n780), .B1(new_n1020), .B2(new_n764), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1021), .B1(new_n647), .B2(new_n706), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n950), .A2(new_n957), .B1(new_n1012), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n995), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(KEYINPUT118), .ZN(new_n1025));
  INV_X1    g0825(.A(KEYINPUT118), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n995), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(G393));
  NOR2_X1   g0828(.A1(new_n938), .A2(new_n656), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n657), .B1(new_n942), .B2(new_n945), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n951), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1031), .A2(new_n663), .A3(new_n953), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n939), .A2(new_n946), .A3(new_n957), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT119), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n757), .A2(new_n260), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n763), .C1(new_n228), .C2(new_n215), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n903), .A2(new_n706), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  OR2_X1    g0837(.A1(new_n1036), .A2(new_n1034), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n735), .A2(G311), .B1(new_n1003), .B2(G317), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n271), .B1(new_n231), .B2(new_n712), .C1(new_n456), .C2(new_n723), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n730), .A2(new_n743), .B1(new_n718), .B2(new_n744), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n800), .B2(new_n714), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n727), .A2(new_n520), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n983), .A2(G77), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n234), .B2(new_n727), .C1(new_n296), .C2(new_n730), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n712), .A2(new_n227), .B1(new_n718), .B2(new_n962), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1047), .A2(new_n390), .A3(new_n1048), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n1049), .B1(new_n332), .B2(new_n714), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n735), .A2(G159), .B1(new_n1003), .B2(G150), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n1044), .A2(new_n1045), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n708), .ZN(new_n1054));
  NAND4_X1  g0854(.A1(new_n1037), .A2(new_n780), .A3(new_n1038), .A4(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1033), .A2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1032), .A2(new_n1056), .ZN(G390));
  NAND2_X1  g0857(.A1(new_n852), .A2(new_n882), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n831), .A2(KEYINPUT39), .A3(new_n833), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(new_n778), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(KEYINPUT54), .B(G143), .Z(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n1064), .A2(new_n730), .B1(new_n784), .B2(new_n727), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT121), .ZN(new_n1066));
  OAI211_X1 g0866(.A(new_n1066), .B(new_n270), .C1(new_n234), .C2(new_n712), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n714), .A2(new_n785), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT53), .Z(new_n1069));
  NOR2_X1   g0869(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n983), .A2(G159), .B1(G125), .B2(new_n741), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1070), .B(new_n1071), .C1(new_n790), .C2(new_n745), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(G128), .B2(new_n1003), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI221_X1 g0874(.A(new_n1046), .B1(new_n743), .B2(new_n718), .C1(new_n421), .C2(new_n727), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n792), .B(new_n1075), .C1(G97), .C2(new_n731), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n270), .B1(G116), .B2(new_n735), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI221_X1 g0878(.A(new_n1078), .B1(new_n227), .B2(new_n714), .C1(new_n800), .C2(new_n726), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n709), .B1(new_n1074), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g0880(.A1(new_n1062), .A2(new_n701), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n781), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1081), .B1(new_n297), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n884), .B1(new_n851), .B2(new_n833), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n770), .A2(new_n435), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n878), .B1(new_n696), .B2(new_n1086), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n877), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1084), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g0889(.A(KEYINPUT120), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n618), .A2(new_n636), .A3(new_n772), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1088), .B1(new_n1091), .B2(new_n769), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1092), .B2(new_n884), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n879), .A2(KEYINPUT120), .A3(new_n885), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n1093), .A2(new_n1094), .A3(new_n1060), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1089), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g0896(.A1(new_n683), .A2(G330), .A3(new_n772), .A4(new_n877), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1089), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1083), .B1(new_n1101), .B2(new_n956), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1088), .B1(new_n684), .B2(new_n771), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1103), .A2(new_n1097), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1105), .A2(new_n1087), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(new_n1103), .A2(new_n1097), .B1(new_n769), .B2(new_n1091), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n862), .B(new_n890), .C1(new_n1106), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1101), .A2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n1089), .A2(new_n1095), .A3(new_n1097), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1097), .B1(new_n1089), .B2(new_n1095), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1107), .B1(new_n1105), .B2(new_n1087), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n889), .A2(new_n452), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n626), .A3(new_n862), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n664), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1102), .B1(new_n1109), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(G378));
  INV_X1    g0919(.A(KEYINPUT57), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1115), .B1(new_n1112), .B2(new_n1116), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1058), .A2(new_n884), .A3(new_n1059), .ZN(new_n1122));
  XOR2_X1   g0922(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n322), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n322), .A2(new_n1124), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1126), .A2(new_n311), .A3(new_n814), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n311), .A2(new_n814), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1127), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1129), .B1(new_n1130), .B2(new_n1125), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1092), .A2(new_n828), .A3(new_n834), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1122), .A2(new_n1132), .A3(new_n1133), .A4(new_n876), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1132), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n880), .B2(new_n886), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n872), .A2(G330), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1134), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n861), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n1120), .B1(new_n1121), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1116), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1115), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1140), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1144), .A2(new_n1145), .A3(KEYINPUT57), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1141), .A2(new_n1146), .A3(new_n663), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1082), .A2(G50), .ZN(new_n1148));
  AOI211_X1 g0948(.A(new_n701), .B(new_n1148), .C1(new_n1132), .C2(new_n778), .ZN(new_n1149));
  INV_X1    g0949(.A(G124), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n264), .B1(new_n718), .B2(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1064), .A2(new_n714), .B1(new_n784), .B2(new_n730), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n735), .A2(G128), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n790), .B2(new_n727), .ZN(new_n1154));
  AOI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(G125), .C2(new_n1003), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1155), .B1(new_n785), .B2(new_n723), .ZN(new_n1156));
  AOI211_X1 g0956(.A(G41), .B(new_n1151), .C1(new_n1156), .C2(KEYINPUT59), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(KEYINPUT59), .B2(new_n1156), .C1(new_n719), .C2(new_n712), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n390), .B1(new_n745), .B2(new_n231), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n283), .B1(new_n712), .B2(new_n238), .C1(new_n206), .C2(new_n714), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n726), .A2(new_n456), .B1(new_n718), .B2(new_n800), .ZN(new_n1161));
  NOR4_X1   g0961(.A1(new_n1159), .A2(new_n964), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n1162), .B1(new_n228), .B2(new_n727), .C1(new_n427), .C2(new_n730), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT58), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1158), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n363), .A2(G33), .ZN(new_n1166));
  AOI21_X1  g0966(.A(G50), .B1(new_n1166), .B2(new_n283), .ZN(new_n1167));
  XOR2_X1   g0967(.A(new_n1167), .B(KEYINPUT122), .Z(new_n1168));
  OAI21_X1  g0968(.A(new_n708), .B1(new_n1165), .B2(new_n1168), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1149), .A2(new_n1169), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n1170), .B1(new_n1140), .B2(new_n956), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1147), .A2(new_n1172), .ZN(G375));
  NAND2_X1  g0973(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1174));
  AND2_X1   g0974(.A1(new_n1108), .A2(new_n1174), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n928), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT123), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1088), .A2(new_n778), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n781), .A2(new_n332), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n271), .B1(new_n745), .B2(new_n800), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1180), .B1(G303), .B2(new_n741), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(new_n422), .A2(new_n731), .B1(new_n747), .B2(G116), .ZN(new_n1182));
  OAI221_X1 g0982(.A(new_n1181), .B1(KEYINPUT124), .B2(new_n1182), .C1(new_n206), .C2(new_n712), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n1182), .A2(KEYINPUT124), .B1(G97), .B2(new_n973), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1184), .B(new_n997), .C1(new_n743), .C2(new_n726), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n730), .A2(new_n785), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n390), .B1(G128), .B2(new_n741), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n1064), .A2(new_n727), .B1(new_n790), .B2(new_n726), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G50), .B2(new_n983), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n973), .A2(G159), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n735), .A2(G137), .B1(G58), .B2(new_n740), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1187), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n1183), .A2(new_n1185), .B1(new_n1186), .B2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1193), .A2(new_n708), .ZN(new_n1194));
  NAND4_X1  g0994(.A1(new_n1178), .A2(new_n780), .A3(new_n1179), .A4(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1113), .B2(new_n956), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1177), .A2(new_n1197), .ZN(G381));
  AOI21_X1  g0998(.A(new_n1140), .B1(new_n1143), .B2(new_n1142), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n664), .B1(new_n1199), .B2(KEYINPUT57), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1171), .B1(new_n1200), .B2(new_n1141), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1118), .ZN(new_n1202));
  INV_X1    g1002(.A(G390), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1177), .A2(new_n805), .A3(new_n1203), .A4(new_n1197), .ZN(new_n1204));
  INV_X1    g1004(.A(G396), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1025), .A2(new_n1205), .A3(new_n1027), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1204), .A2(G387), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1202), .B1(new_n1207), .B2(KEYINPUT125), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(KEYINPUT125), .B2(new_n1207), .ZN(G407));
  OAI211_X1 g1009(.A(G407), .B(G213), .C1(new_n633), .C2(new_n1202), .ZN(G409));
  NAND3_X1  g1010(.A1(new_n958), .A2(new_n992), .A3(G390), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n995), .A2(new_n1023), .A3(new_n1026), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1026), .B1(new_n995), .B2(new_n1023), .ZN(new_n1213));
  OAI21_X1  g1013(.A(G396), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g1014(.A1(new_n1214), .A2(new_n1206), .A3(KEYINPUT127), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1211), .A2(new_n1215), .ZN(new_n1216));
  AND2_X1   g1016(.A1(new_n1214), .A2(new_n1206), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1217), .A2(new_n958), .A3(new_n992), .A4(G390), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(G387), .A2(new_n1203), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1220), .A2(new_n1215), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1144), .A2(new_n1145), .A3(new_n928), .ZN(new_n1224));
  AND3_X1   g1024(.A1(new_n1118), .A2(new_n1172), .A3(new_n1224), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G375), .B2(G378), .ZN(new_n1226));
  AOI21_X1  g1026(.A(KEYINPUT60), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1108), .A2(new_n1174), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n664), .B(new_n1227), .C1(new_n1228), .C2(KEYINPUT60), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(new_n1229), .A2(new_n805), .A3(new_n1196), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(KEYINPUT60), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1227), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n663), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(G384), .B1(new_n1233), .B2(new_n1197), .ZN(new_n1234));
  NOR2_X1   g1034(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n634), .A2(G213), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1226), .A2(KEYINPUT63), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(KEYINPUT61), .ZN(new_n1238));
  AND3_X1   g1038(.A1(new_n1223), .A2(new_n1237), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT63), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT126), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1118), .B1(new_n1147), .B2(new_n1172), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(new_n1225), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1118), .A2(new_n1172), .A3(new_n1224), .ZN(new_n1244));
  OAI211_X1 g1044(.A(KEYINPUT126), .B(new_n1244), .C1(new_n1201), .C2(new_n1118), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1245), .A3(new_n1236), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n634), .A2(G213), .A3(G2897), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1247), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n805), .B1(new_n1229), .B2(new_n1196), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1233), .A2(G384), .A3(new_n1197), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1247), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1248), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1240), .B1(new_n1246), .B2(new_n1253), .ZN(new_n1254));
  NAND4_X1  g1054(.A1(new_n1243), .A2(new_n1245), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1239), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1223), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1255), .A2(KEYINPUT62), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1244), .B(new_n1236), .C1(new_n1201), .C2(new_n1118), .ZN(new_n1260));
  AOI21_X1  g1060(.A(KEYINPUT61), .B1(new_n1253), .B2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1235), .ZN(new_n1262));
  OAI21_X1  g1062(.A(KEYINPUT62), .B1(new_n1260), .B2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1259), .B2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1257), .A2(new_n1265), .ZN(G405));
  INV_X1    g1066(.A(new_n1242), .ZN(new_n1267));
  AND3_X1   g1067(.A1(new_n1202), .A2(new_n1262), .A3(new_n1267), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1262), .B1(new_n1202), .B2(new_n1267), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(new_n1258), .ZN(G402));
endmodule


