//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 1 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:58 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G97), .ZN(new_n209));
  INV_X1    g0009(.A(G257), .ZN(new_n210));
  OAI22_X1  g0010(.A1(new_n207), .A2(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g0011(.A(new_n211), .B1(G87), .B2(G250), .ZN(new_n212));
  INV_X1    g0012(.A(G116), .ZN(new_n213));
  INV_X1    g0013(.A(G270), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G50), .B2(G226), .ZN(new_n216));
  INV_X1    g0016(.A(G58), .ZN(new_n217));
  INV_X1    g0017(.A(G232), .ZN(new_n218));
  INV_X1    g0018(.A(G107), .ZN(new_n219));
  INV_X1    g0019(.A(G264), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  OAI21_X1  g0024(.A(new_n203), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(G20), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(G50), .B1(G58), .B2(G68), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n226), .C1(new_n229), .C2(new_n231), .ZN(G361));
  XOR2_X1   g0032(.A(G226), .B(G232), .Z(new_n233));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT65), .B(G250), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n237), .B(new_n241), .Z(G358));
  XNOR2_X1  g0042(.A(KEYINPUT66), .B(G87), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n213), .ZN(new_n244));
  AND2_X1   g0044(.A1(G97), .A2(G107), .ZN(new_n245));
  NOR2_X1   g0045(.A1(G97), .A2(G107), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G68), .B(G77), .Z(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n227), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G58), .A2(G68), .ZN(new_n255));
  INV_X1    g0055(.A(G50), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n228), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT67), .ZN(new_n258));
  XNOR2_X1  g0058(.A(KEYINPUT8), .B(G58), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(G20), .ZN(new_n261));
  INV_X1    g0061(.A(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G150), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  OAI22_X1  g0065(.A1(new_n259), .A2(new_n262), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n254), .B1(new_n258), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(G13), .A3(G20), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n268), .A2(KEYINPUT68), .A3(G13), .A4(G20), .ZN(new_n272));
  AND2_X1   g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n256), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n254), .B1(new_n271), .B2(new_n272), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G1), .B2(new_n228), .ZN(new_n276));
  OAI211_X1 g0076(.A(new_n267), .B(new_n274), .C1(new_n256), .C2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT9), .ZN(new_n278));
  OR2_X1    g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n277), .A2(new_n278), .ZN(new_n280));
  XNOR2_X1  g0080(.A(KEYINPUT3), .B(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(G222), .A2(G1698), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G223), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n285), .B(new_n288), .C1(G77), .C2(new_n281), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n268), .B(G274), .C1(G41), .C2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(G226), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n287), .A2(new_n292), .ZN(new_n293));
  OAI211_X1 g0093(.A(new_n289), .B(new_n290), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(G200), .ZN(new_n295));
  INV_X1    g0095(.A(G190), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g0097(.A1(new_n279), .A2(new_n280), .A3(new_n295), .A4(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n298), .A2(KEYINPUT10), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n294), .A2(G179), .ZN(new_n303));
  INV_X1    g0103(.A(G169), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n294), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n303), .A2(new_n277), .A3(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(new_n276), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G77), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n271), .A2(new_n272), .ZN(new_n309));
  XOR2_X1   g0109(.A(KEYINPUT15), .B(G87), .Z(new_n310));
  NAND3_X1  g0110(.A1(new_n310), .A2(KEYINPUT70), .A3(new_n261), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT70), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT15), .B(G87), .ZN(new_n313));
  OAI21_X1  g0113(.A(new_n312), .B1(new_n313), .B2(new_n262), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  OAI22_X1  g0115(.A1(new_n259), .A2(new_n265), .B1(new_n228), .B2(new_n207), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n254), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  AND2_X1   g0117(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n318));
  NOR2_X1   g0118(.A1(new_n317), .A2(KEYINPUT71), .ZN(new_n319));
  OAI221_X1 g0119(.A(new_n308), .B1(G77), .B2(new_n309), .C1(new_n318), .C2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n281), .A2(G238), .A3(G1698), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n281), .A2(G232), .A3(new_n283), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G33), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(G107), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n321), .A2(new_n322), .A3(new_n327), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(KEYINPUT69), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n329), .A2(new_n288), .A3(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n290), .ZN(new_n332));
  INV_X1    g0132(.A(new_n293), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n332), .B1(new_n333), .B2(G244), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n335), .A2(new_n304), .ZN(new_n336));
  INV_X1    g0136(.A(G179), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n331), .A2(new_n337), .A3(new_n334), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n320), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n302), .A2(new_n306), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(new_n254), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n261), .A2(G77), .B1(G20), .B2(new_n222), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n264), .A2(G50), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n345), .B(KEYINPUT11), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n273), .A2(new_n222), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT12), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n307), .A2(G68), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n324), .A2(new_n325), .A3(G232), .A4(G1698), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(KEYINPUT73), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT73), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n281), .A2(new_n353), .A3(G232), .A4(G1698), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n281), .A2(G226), .A3(new_n283), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n356), .B1(new_n260), .B2(new_n209), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n288), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n290), .B1(new_n293), .B2(new_n223), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(KEYINPUT74), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT74), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n361), .B(new_n290), .C1(new_n293), .C2(new_n223), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n358), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT13), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT13), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n358), .A2(new_n363), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n350), .B1(new_n368), .B2(G200), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n365), .A2(G190), .A3(new_n367), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(KEYINPUT75), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT75), .ZN(new_n372));
  NAND4_X1  g0172(.A1(new_n365), .A2(new_n372), .A3(G190), .A4(new_n367), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n369), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT76), .ZN(new_n375));
  AND3_X1   g0175(.A1(new_n358), .A2(new_n363), .A3(new_n366), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n366), .B1(new_n358), .B2(new_n363), .ZN(new_n377));
  OAI21_X1  g0177(.A(G169), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT14), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n365), .A2(G179), .A3(new_n367), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n381), .B(G169), .C1(new_n376), .C2(new_n377), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n380), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n350), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT76), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n369), .A2(new_n371), .A3(new_n385), .A4(new_n373), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n375), .A2(new_n384), .A3(new_n386), .ZN(new_n387));
  OR2_X1    g0187(.A1(new_n387), .A2(KEYINPUT77), .ZN(new_n388));
  INV_X1    g0188(.A(new_n320), .ZN(new_n389));
  INV_X1    g0189(.A(G200), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n331), .B2(new_n334), .ZN(new_n391));
  INV_X1    g0191(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n389), .A2(KEYINPUT72), .A3(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT72), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n394), .B1(new_n320), .B2(new_n391), .ZN(new_n395));
  AND2_X1   g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n331), .A2(G190), .A3(new_n334), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n387), .A2(KEYINPUT77), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT18), .ZN(new_n399));
  INV_X1    g0199(.A(new_n259), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n273), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n401), .B1(new_n276), .B2(new_n400), .ZN(new_n402));
  XNOR2_X1  g0202(.A(KEYINPUT78), .B(G33), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n325), .B1(new_n403), .B2(KEYINPUT3), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT7), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(G20), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n326), .A2(new_n228), .ZN(new_n407));
  AOI22_X1  g0207(.A1(new_n404), .A2(new_n406), .B1(new_n407), .B2(new_n405), .ZN(new_n408));
  OAI21_X1  g0208(.A(KEYINPUT79), .B1(new_n408), .B2(new_n222), .ZN(new_n409));
  XNOR2_X1  g0209(.A(G58), .B(G68), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n410), .A2(G20), .B1(G159), .B2(new_n264), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n260), .A2(KEYINPUT78), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT78), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(G33), .ZN(new_n414));
  AOI21_X1  g0214(.A(KEYINPUT3), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n325), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n406), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n405), .B1(new_n281), .B2(G20), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT79), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(G68), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(new_n411), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n412), .A2(new_n414), .A3(KEYINPUT3), .ZN(new_n425));
  AOI21_X1  g0225(.A(G20), .B1(new_n425), .B2(new_n324), .ZN(new_n426));
  OAI21_X1  g0226(.A(G68), .B1(new_n426), .B2(new_n405), .ZN(new_n427));
  AOI211_X1 g0227(.A(KEYINPUT7), .B(G20), .C1(new_n425), .C2(new_n324), .ZN(new_n428));
  OAI211_X1 g0228(.A(KEYINPUT16), .B(new_n411), .C1(new_n427), .C2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n429), .A2(new_n254), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n402), .B1(new_n424), .B2(new_n430), .ZN(new_n431));
  OR2_X1    g0231(.A1(G223), .A2(G1698), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n291), .A2(G1698), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n425), .A2(new_n324), .A3(new_n432), .A4(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(G33), .A2(G87), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(new_n288), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n290), .B1(new_n293), .B2(new_n218), .ZN(new_n438));
  INV_X1    g0238(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n337), .A3(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT80), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n287), .B1(new_n434), .B2(new_n435), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n304), .B1(new_n442), .B2(new_n438), .ZN(new_n443));
  AND3_X1   g0243(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n441), .B1(new_n440), .B2(new_n443), .ZN(new_n445));
  NOR2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n399), .B1(new_n431), .B2(new_n446), .ZN(new_n447));
  AOI21_X1  g0247(.A(G169), .B1(new_n437), .B2(new_n439), .ZN(new_n448));
  NOR3_X1   g0248(.A1(new_n442), .A2(G179), .A3(new_n438), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT80), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n440), .A2(new_n441), .A3(new_n443), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n429), .A2(new_n254), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n423), .B2(new_n422), .ZN(new_n454));
  OAI211_X1 g0254(.A(new_n452), .B(KEYINPUT18), .C1(new_n454), .C2(new_n402), .ZN(new_n455));
  AND2_X1   g0255(.A1(new_n447), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n424), .A2(new_n430), .ZN(new_n457));
  INV_X1    g0257(.A(new_n402), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n437), .A2(new_n439), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n390), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(G190), .B2(new_n459), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n457), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT17), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n431), .A2(KEYINPUT17), .A3(new_n461), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n456), .A2(new_n466), .ZN(new_n467));
  AND4_X1   g0267(.A1(new_n341), .A2(new_n388), .A3(new_n398), .A4(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(G87), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n470), .A2(G20), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n425), .A2(new_n324), .A3(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT91), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n425), .A2(KEYINPUT91), .A3(new_n324), .A4(new_n471), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(KEYINPUT22), .A3(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT22), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n281), .A2(new_n477), .A3(new_n471), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n412), .A2(new_n414), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(new_n228), .A3(G116), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n219), .A2(G20), .ZN(new_n482));
  AOI21_X1  g0282(.A(new_n482), .B1(KEYINPUT92), .B2(KEYINPUT23), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT92), .A2(KEYINPUT23), .ZN(new_n484));
  MUX2_X1   g0284(.A(new_n483), .B(new_n482), .S(new_n484), .Z(new_n485));
  NAND3_X1  g0285(.A1(new_n479), .A2(new_n481), .A3(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT24), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n479), .A2(KEYINPUT24), .A3(new_n481), .A4(new_n485), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n488), .A2(new_n254), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(KEYINPUT83), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n268), .A2(G33), .ZN(new_n492));
  AND4_X1   g0292(.A1(new_n491), .A2(new_n309), .A3(new_n342), .A4(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n275), .B2(new_n492), .ZN(new_n494));
  OAI21_X1  g0294(.A(G107), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(KEYINPUT25), .B1(new_n309), .B2(G107), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n309), .A2(KEYINPUT25), .A3(G107), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n495), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n498), .A2(KEYINPUT93), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT93), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n495), .A2(new_n500), .A3(new_n496), .A4(new_n497), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G41), .ZN(new_n503));
  AND3_X1   g0303(.A1(new_n503), .A2(KEYINPUT85), .A3(KEYINPUT5), .ZN(new_n504));
  AOI21_X1  g0304(.A(KEYINPUT5), .B1(new_n503), .B2(KEYINPUT85), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n268), .A2(G45), .A3(G274), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(G250), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(new_n283), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n210), .A2(G1698), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n425), .A2(new_n324), .A3(new_n509), .A4(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n480), .A2(G294), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n288), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n287), .B1(new_n504), .B2(new_n505), .ZN(new_n515));
  INV_X1    g0315(.A(G45), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n287), .B1(G1), .B2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n220), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT94), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n514), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n287), .B1(new_n511), .B2(new_n512), .ZN(new_n522));
  OAI21_X1  g0322(.A(KEYINPUT94), .B1(new_n522), .B2(new_n518), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n507), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n507), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n514), .A2(new_n519), .A3(new_n525), .ZN(new_n526));
  OAI22_X1  g0326(.A1(new_n524), .A2(G200), .B1(G190), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n490), .A2(new_n502), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G169), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n524), .A2(G179), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n490), .A2(new_n502), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g0331(.A1(new_n528), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n425), .A2(G244), .A3(new_n283), .A4(new_n324), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT4), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n324), .A2(new_n325), .A3(G250), .A4(G1698), .ZN(new_n536));
  AND2_X1   g0336(.A1(KEYINPUT4), .A2(G244), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n324), .A2(new_n325), .A3(new_n537), .A4(new_n283), .ZN(new_n538));
  NAND2_X1  g0338(.A1(G33), .A2(G283), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n536), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT84), .ZN(new_n542));
  INV_X1    g0342(.A(KEYINPUT84), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n535), .A2(new_n543), .A3(new_n540), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n542), .A2(new_n288), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n515), .A2(new_n517), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n507), .B1(new_n546), .B2(G257), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(G200), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n209), .A2(G107), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT6), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(KEYINPUT81), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT81), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT6), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n550), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n555), .B1(new_n247), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G20), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n264), .A2(G77), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n219), .B1(new_n417), .B2(new_n418), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n254), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n557), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(new_n408), .B2(new_n219), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(KEYINPUT82), .A3(new_n254), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n275), .A2(new_n492), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(KEYINPUT83), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n275), .A2(new_n491), .A3(new_n492), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n564), .A2(new_n567), .B1(G97), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n309), .A2(G97), .ZN(new_n573));
  INV_X1    g0373(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n545), .A2(G190), .A3(new_n547), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n549), .A2(new_n572), .A3(new_n574), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n571), .A2(G97), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n562), .A2(new_n563), .ZN(new_n578));
  AOI21_X1  g0378(.A(KEYINPUT82), .B1(new_n566), .B2(new_n254), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n574), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n548), .A2(new_n304), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n545), .A2(new_n337), .A3(new_n547), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n580), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n576), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n214), .B1(new_n515), .B2(new_n517), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n210), .A2(new_n283), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n220), .A2(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n425), .A2(new_n324), .A3(new_n587), .A4(new_n588), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n326), .A2(G303), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g0391(.A(new_n586), .B(new_n525), .C1(new_n591), .C2(new_n287), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n592), .A2(new_n337), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n275), .A2(G116), .A3(new_n492), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n273), .A2(new_n213), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n213), .A2(G20), .ZN(new_n596));
  AOI21_X1  g0396(.A(G20), .B1(G33), .B2(G283), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n260), .A2(G97), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n597), .A2(new_n598), .A3(KEYINPUT90), .ZN(new_n599));
  AOI21_X1  g0399(.A(KEYINPUT90), .B1(new_n597), .B2(new_n598), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n254), .B(new_n596), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT20), .ZN(new_n602));
  AND2_X1   g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n601), .A2(new_n602), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n594), .B(new_n595), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n593), .A2(new_n605), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT89), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n287), .B1(new_n589), .B2(new_n590), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n608), .A2(new_n507), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n607), .B1(new_n609), .B2(new_n586), .ZN(new_n610));
  NOR4_X1   g0410(.A1(new_n608), .A2(new_n585), .A3(KEYINPUT89), .A4(new_n507), .ZN(new_n611));
  OAI21_X1  g0411(.A(G200), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n592), .A2(KEYINPUT89), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n609), .A2(new_n607), .A3(new_n586), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(G190), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n605), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n612), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  OAI211_X1 g0417(.A(G169), .B(new_n605), .C1(new_n610), .C2(new_n611), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT21), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n613), .A2(new_n614), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(KEYINPUT21), .A3(G169), .A4(new_n605), .ZN(new_n622));
  AND4_X1   g0422(.A1(new_n606), .A2(new_n617), .A3(new_n620), .A4(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT88), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT87), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n506), .B1(new_n517), .B2(new_n508), .ZN(new_n626));
  NOR2_X1   g0426(.A1(G238), .A2(G1698), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n627), .B1(new_n208), .B2(G1698), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n628), .A2(new_n425), .A3(new_n324), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n480), .A2(G116), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n626), .B1(new_n631), .B2(new_n288), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n625), .B1(new_n632), .B2(G190), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n287), .B1(new_n629), .B2(new_n630), .ZN(new_n634));
  NOR4_X1   g0434(.A1(new_n634), .A2(KEYINPUT87), .A3(new_n626), .A4(new_n296), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n624), .B1(new_n633), .B2(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(new_n626), .ZN(new_n637));
  INV_X1    g0437(.A(new_n324), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n403), .B2(KEYINPUT3), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n639), .A2(new_n628), .B1(G116), .B2(new_n480), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n637), .B(G190), .C1(new_n640), .C2(new_n287), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT87), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n632), .A2(new_n625), .A3(G190), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n642), .A2(new_n643), .A3(KEYINPUT88), .ZN(new_n644));
  INV_X1    g0444(.A(new_n632), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n309), .A2(new_n310), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n222), .A2(G20), .ZN(new_n649));
  NOR3_X1   g0449(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n650));
  AOI21_X1  g0450(.A(G20), .B1(G33), .B2(G97), .ZN(new_n651));
  OAI21_X1  g0451(.A(KEYINPUT19), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT19), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n261), .A2(new_n653), .A3(G97), .ZN(new_n654));
  AOI22_X1  g0454(.A1(new_n639), .A2(new_n649), .B1(new_n652), .B2(new_n654), .ZN(new_n655));
  OAI211_X1 g0455(.A(new_n648), .B(KEYINPUT86), .C1(new_n655), .C2(new_n342), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT86), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n652), .A2(new_n654), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n425), .A2(new_n324), .A3(new_n649), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n342), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n657), .B1(new_n660), .B2(new_n647), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n656), .A2(new_n661), .B1(new_n571), .B2(G87), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n636), .A2(new_n644), .A3(new_n646), .A4(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n656), .A2(new_n661), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n571), .A2(new_n310), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n632), .A2(new_n337), .ZN(new_n667));
  OAI211_X1 g0467(.A(new_n666), .B(new_n667), .C1(G169), .C2(new_n632), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n532), .A2(new_n584), .A3(new_n623), .A4(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n469), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g0472(.A(new_n672), .B(KEYINPUT95), .Z(G372));
  INV_X1    g0473(.A(new_n306), .ZN(new_n674));
  INV_X1    g0474(.A(new_n339), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(new_n374), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n384), .ZN(new_n677));
  AND4_X1   g0477(.A1(KEYINPUT17), .A2(new_n457), .A3(new_n458), .A4(new_n461), .ZN(new_n678));
  AOI21_X1  g0478(.A(KEYINPUT17), .B1(new_n431), .B2(new_n461), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n456), .B1(new_n677), .B2(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT98), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI22_X1  g0483(.A1(new_n681), .A2(new_n682), .B1(new_n301), .B2(new_n300), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n674), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n620), .A2(new_n622), .A3(new_n606), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n490), .A2(new_n502), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n530), .A2(new_n529), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT96), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n634), .A2(new_n691), .ZN(new_n692));
  AOI211_X1 g0492(.A(KEYINPUT96), .B(new_n287), .C1(new_n629), .C2(new_n630), .ZN(new_n693));
  OAI21_X1  g0493(.A(new_n637), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n304), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n695), .A2(new_n666), .A3(new_n667), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(G200), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n642), .A2(new_n643), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n697), .A2(new_n698), .A3(new_n662), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n696), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT97), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT97), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n528), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n690), .A2(new_n704), .A3(new_n584), .A4(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT26), .ZN(new_n707));
  INV_X1    g0507(.A(new_n583), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n704), .A2(new_n707), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT26), .B1(new_n669), .B2(new_n583), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n706), .A2(new_n696), .A3(new_n709), .A4(new_n710), .ZN(new_n711));
  INV_X1    g0511(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n685), .B1(new_n469), .B2(new_n712), .ZN(G369));
  INV_X1    g0513(.A(G13), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G20), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(new_n268), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n716), .A2(KEYINPUT27), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G213), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(G343), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n605), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n623), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n686), .B2(new_n722), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(G330), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n687), .A2(new_n721), .ZN(new_n726));
  AOI22_X1  g0526(.A1(new_n532), .A2(new_n726), .B1(new_n531), .B2(new_n721), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n686), .B2(new_n721), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n725), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n620), .A2(new_n622), .A3(new_n606), .ZN(new_n730));
  INV_X1    g0530(.A(new_n721), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n532), .A2(new_n730), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n531), .A2(new_n731), .ZN(new_n733));
  AND2_X1   g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n729), .A2(new_n734), .ZN(G399));
  INV_X1    g0535(.A(new_n204), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(G41), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n650), .A2(new_n213), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n738), .A2(G1), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(new_n230), .B2(new_n738), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n742), .B(KEYINPUT28), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT29), .ZN(new_n744));
  AND3_X1   g0544(.A1(new_n711), .A2(new_n744), .A3(new_n731), .ZN(new_n745));
  AND2_X1   g0545(.A1(new_n545), .A2(new_n547), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n521), .A2(new_n523), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n592), .A2(new_n645), .A3(new_n337), .ZN(new_n748));
  NAND4_X1  g0548(.A1(new_n746), .A2(KEYINPUT30), .A3(new_n747), .A4(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n545), .A2(new_n747), .A3(new_n547), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n593), .A2(new_n632), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND4_X1  g0553(.A1(new_n621), .A2(new_n548), .A3(new_n337), .A4(new_n694), .ZN(new_n754));
  OAI211_X1 g0554(.A(new_n749), .B(new_n753), .C1(new_n524), .C2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT31), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n755), .A2(new_n756), .A3(new_n721), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n756), .B1(new_n755), .B2(new_n721), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n671), .A2(new_n721), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n759), .A2(G330), .ZN(new_n760));
  NOR3_X1   g0560(.A1(new_n669), .A2(new_n583), .A3(KEYINPUT26), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n696), .A2(new_n699), .A3(new_n702), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n702), .B1(new_n696), .B2(new_n699), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n708), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g0564(.A(new_n761), .B1(new_n764), .B2(KEYINPUT26), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n765), .A2(new_n706), .A3(new_n696), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n744), .B1(new_n766), .B2(new_n731), .ZN(new_n767));
  NOR3_X1   g0567(.A1(new_n745), .A2(new_n760), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n743), .B1(new_n768), .B2(G1), .ZN(G364));
  NAND2_X1  g0569(.A1(new_n715), .A2(G45), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n738), .A2(G1), .A3(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n725), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n773), .B1(G330), .B2(new_n724), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n231), .A2(new_n516), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n639), .A2(new_n736), .ZN(new_n776));
  OAI211_X1 g0576(.A(new_n775), .B(new_n776), .C1(new_n251), .C2(new_n516), .ZN(new_n777));
  INV_X1    g0577(.A(G355), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n281), .A2(new_n204), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n777), .B1(G116), .B2(new_n204), .C1(new_n778), .C2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(G13), .A2(G33), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(G20), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n227), .B1(G20), .B2(new_n304), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  XOR2_X1   g0585(.A(new_n785), .B(KEYINPUT99), .Z(new_n786));
  AOI21_X1  g0586(.A(new_n771), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  XOR2_X1   g0587(.A(new_n787), .B(KEYINPUT100), .Z(new_n788));
  INV_X1    g0588(.A(new_n784), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n228), .A2(new_n296), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n337), .A2(G200), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n228), .A2(G190), .ZN(new_n794));
  NOR2_X1   g0594(.A1(G179), .A2(G200), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(G322), .A2(new_n793), .B1(new_n797), .B2(G329), .ZN(new_n798));
  INV_X1    g0598(.A(G294), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n228), .B1(new_n795), .B2(G190), .ZN(new_n800));
  OAI211_X1 g0600(.A(new_n798), .B(new_n326), .C1(new_n799), .C2(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n337), .A2(new_n390), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(G326), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n390), .A2(G179), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n794), .ZN(new_n806));
  INV_X1    g0606(.A(G283), .ZN(new_n807));
  OAI22_X1  g0607(.A1(new_n803), .A2(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  XOR2_X1   g0608(.A(KEYINPUT33), .B(G317), .Z(new_n809));
  NAND2_X1  g0609(.A1(new_n802), .A2(new_n794), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n794), .A2(new_n791), .ZN(new_n811));
  INV_X1    g0611(.A(G311), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n801), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(G303), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n790), .A2(new_n805), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G159), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n796), .A2(new_n818), .ZN(new_n819));
  XOR2_X1   g0619(.A(KEYINPUT101), .B(KEYINPUT32), .Z(new_n820));
  OAI22_X1  g0620(.A1(new_n819), .A2(new_n820), .B1(new_n207), .B2(new_n811), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n800), .A2(new_n209), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n803), .A2(new_n256), .B1(new_n806), .B2(new_n219), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n819), .A2(new_n820), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n222), .A2(new_n810), .B1(new_n816), .B2(new_n470), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G58), .B2(new_n793), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n281), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n817), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n783), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n788), .B1(new_n789), .B2(new_n829), .C1(new_n724), .C2(new_n830), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n774), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NOR2_X1   g0633(.A1(new_n339), .A2(new_n721), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n393), .A2(new_n397), .A3(new_n395), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n835), .B1(new_n389), .B2(new_n731), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n834), .B1(new_n836), .B2(new_n339), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n838), .B1(new_n712), .B2(new_n721), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n711), .A2(new_n731), .A3(new_n837), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(new_n760), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n842), .A2(new_n771), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n838), .A2(new_n781), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n784), .A2(new_n781), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n207), .ZN(new_n846));
  INV_X1    g0646(.A(new_n816), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n822), .B1(G107), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(new_n213), .B2(new_n811), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n326), .B1(new_n796), .B2(new_n812), .C1(new_n799), .C2(new_n792), .ZN(new_n850));
  OAI22_X1  g0650(.A1(new_n803), .A2(new_n815), .B1(new_n806), .B2(new_n470), .ZN(new_n851));
  NOR3_X1   g0651(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(new_n807), .B2(new_n810), .ZN(new_n853));
  INV_X1    g0653(.A(G132), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n639), .B1(new_n854), .B2(new_n796), .ZN(new_n855));
  INV_X1    g0655(.A(new_n811), .ZN(new_n856));
  AOI22_X1  g0656(.A1(G143), .A2(new_n793), .B1(new_n856), .B2(G159), .ZN(new_n857));
  INV_X1    g0657(.A(G137), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n857), .B1(new_n858), .B2(new_n803), .C1(new_n263), .C2(new_n810), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n806), .ZN(new_n862));
  AOI22_X1  g0662(.A1(G50), .A2(new_n847), .B1(new_n862), .B2(G68), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(new_n860), .C2(new_n859), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n800), .A2(new_n217), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n853), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  XOR2_X1   g0666(.A(new_n866), .B(KEYINPUT102), .Z(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n784), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n844), .A2(new_n772), .A3(new_n846), .A4(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n843), .A2(new_n869), .ZN(G384));
  NAND3_X1  g0670(.A1(new_n468), .A2(G330), .A3(new_n759), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT38), .ZN(new_n872));
  OAI21_X1  g0672(.A(KEYINPUT7), .B1(new_n639), .B2(G20), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n426), .A2(new_n405), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n873), .A2(new_n874), .A3(G68), .ZN(new_n875));
  AOI21_X1  g0675(.A(KEYINPUT16), .B1(new_n875), .B2(new_n411), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n458), .B1(new_n453), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n452), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n719), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n462), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n454), .A2(new_n402), .B1(new_n452), .B2(new_n879), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT37), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(new_n462), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n882), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n447), .A2(new_n455), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n880), .B1(new_n680), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n872), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n880), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n456), .B2(new_n466), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n882), .A2(new_n885), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n893));
  AND3_X1   g0693(.A1(new_n889), .A2(KEYINPUT105), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g0694(.A(KEYINPUT105), .B1(new_n889), .B2(new_n893), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n350), .A2(new_n721), .ZN(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n387), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n384), .A2(new_n374), .A3(new_n896), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n759), .A2(new_n837), .A3(new_n900), .ZN(new_n901));
  NOR3_X1   g0701(.A1(new_n894), .A2(new_n895), .A3(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(G330), .B1(new_n902), .B2(KEYINPUT40), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT107), .ZN(new_n904));
  AND3_X1   g0704(.A1(new_n891), .A2(KEYINPUT38), .A3(new_n892), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n431), .A2(new_n719), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n906), .B1(new_n456), .B2(new_n466), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n883), .A2(new_n462), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT37), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n885), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n907), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT40), .B1(new_n905), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n904), .B1(new_n912), .B2(new_n901), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n759), .A2(new_n837), .A3(new_n900), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT40), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n909), .A2(new_n885), .ZN(new_n916));
  INV_X1    g0716(.A(new_n906), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n917), .B1(new_n680), .B2(new_n887), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n872), .B1(new_n916), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n915), .B1(new_n919), .B2(new_n893), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n914), .A2(new_n920), .A3(KEYINPUT107), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n913), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n871), .B1(new_n903), .B2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n902), .A2(KEYINPUT40), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n913), .A2(new_n921), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n925), .A2(new_n468), .A3(new_n759), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n923), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n468), .B1(new_n745), .B2(new_n767), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n928), .A2(new_n685), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n927), .B(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n834), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n840), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(new_n900), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT104), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n894), .A2(new_n895), .ZN(new_n936));
  INV_X1    g0736(.A(new_n900), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(new_n840), .B2(new_n931), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n938), .A2(KEYINPUT104), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n935), .A2(new_n936), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(KEYINPUT106), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n911), .A2(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n889), .A2(new_n893), .ZN(new_n943));
  OAI21_X1  g0743(.A(KEYINPUT39), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT39), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n919), .A2(new_n941), .A3(new_n893), .A4(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n384), .A2(new_n721), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n947), .A2(new_n948), .B1(new_n456), .B2(new_n719), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n940), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n930), .B(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n268), .B2(new_n715), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n213), .B1(new_n557), .B2(KEYINPUT35), .ZN(new_n953));
  OAI211_X1 g0753(.A(new_n953), .B(new_n229), .C1(KEYINPUT35), .C2(new_n557), .ZN(new_n954));
  XNOR2_X1  g0754(.A(new_n954), .B(KEYINPUT36), .ZN(new_n955));
  OAI211_X1 g0755(.A(new_n231), .B(G77), .C1(new_n217), .C2(new_n222), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n956), .B(KEYINPUT103), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(G50), .B2(new_n222), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n958), .A2(G1), .A3(new_n714), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n952), .A2(new_n955), .A3(new_n959), .ZN(G367));
  NOR2_X1   g0760(.A1(new_n313), .A2(new_n204), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n241), .A2(new_n776), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n785), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n796), .A2(new_n858), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n810), .A2(new_n818), .B1(new_n811), .B2(new_n256), .ZN(new_n965));
  INV_X1    g0765(.A(new_n803), .ZN(new_n966));
  AOI211_X1 g0766(.A(new_n964), .B(new_n965), .C1(G143), .C2(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n793), .A2(G150), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n800), .A2(new_n222), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n969), .A2(new_n326), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n806), .A2(new_n207), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G58), .B2(new_n847), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n967), .A2(new_n968), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n816), .A2(new_n213), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n806), .A2(new_n209), .ZN(new_n976));
  INV_X1    g0776(.A(G317), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n796), .A2(new_n977), .ZN(new_n978));
  NOR4_X1   g0778(.A1(new_n975), .A2(new_n639), .A3(new_n976), .A4(new_n978), .ZN(new_n979));
  AOI22_X1  g0779(.A1(G311), .A2(new_n966), .B1(new_n793), .B2(G303), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n811), .A2(new_n807), .B1(new_n800), .B2(new_n219), .ZN(new_n981));
  XOR2_X1   g0781(.A(new_n981), .B(KEYINPUT110), .Z(new_n982));
  NAND3_X1  g0782(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n810), .A2(new_n799), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n973), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT47), .Z(new_n986));
  OAI221_X1 g0786(.A(new_n772), .B1(new_n961), .B2(new_n963), .C1(new_n986), .C2(new_n789), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n987), .B(KEYINPUT111), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n704), .B1(new_n662), .B2(new_n731), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n662), .A2(new_n731), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n989), .B1(new_n696), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n988), .B1(new_n830), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n770), .A2(G1), .ZN(new_n993));
  INV_X1    g0793(.A(new_n580), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n584), .B1(new_n994), .B2(new_n731), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n708), .A2(new_n721), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n995), .A2(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n734), .A2(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT44), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n734), .A2(new_n997), .ZN(new_n1000));
  XOR2_X1   g0800(.A(KEYINPUT108), .B(KEYINPUT45), .Z(new_n1001));
  XNOR2_X1  g0801(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n999), .A2(new_n729), .A3(new_n1002), .ZN(new_n1003));
  OR2_X1    g0803(.A1(new_n725), .A2(new_n728), .ZN(new_n1004));
  AND3_X1   g0804(.A1(new_n1004), .A2(new_n729), .A3(new_n732), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1003), .A2(new_n768), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT109), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1003), .A2(KEYINPUT109), .A3(new_n768), .A4(new_n1005), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(new_n768), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n737), .B(KEYINPUT41), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n993), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n997), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n1014), .A2(new_n732), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT42), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n583), .B1(new_n995), .B2(new_n689), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n731), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OR3_X1    g0819(.A1(new_n1019), .A2(KEYINPUT43), .A3(new_n991), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n729), .A2(new_n1014), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n1022), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n991), .A2(KEYINPUT43), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n1019), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AND3_X1   g0825(.A1(new_n1020), .A2(new_n1021), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1021), .B1(new_n1020), .B2(new_n1025), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n992), .B1(new_n1013), .B2(new_n1028), .ZN(G387));
  OR2_X1    g0829(.A1(new_n1005), .A2(new_n768), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1005), .A2(new_n768), .ZN(new_n1031));
  NAND3_X1  g0831(.A1(new_n1030), .A2(new_n737), .A3(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n810), .A2(new_n259), .B1(new_n800), .B2(new_n313), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(KEYINPUT112), .B(G150), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n976), .B(new_n1033), .C1(new_n797), .C2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n793), .A2(G50), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n803), .A2(new_n818), .B1(new_n816), .B2(new_n207), .ZN(new_n1037));
  AOI21_X1  g0837(.A(new_n1037), .B1(G68), .B2(new_n856), .ZN(new_n1038));
  NAND4_X1  g0838(.A1(new_n1035), .A2(new_n639), .A3(new_n1036), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g0839(.A(new_n810), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(G322), .A2(new_n966), .B1(new_n1040), .B2(G311), .ZN(new_n1041));
  OAI221_X1 g0841(.A(new_n1041), .B1(new_n815), .B2(new_n811), .C1(new_n977), .C2(new_n792), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT48), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n807), .B2(new_n800), .C1(new_n799), .C2(new_n816), .ZN(new_n1044));
  XOR2_X1   g0844(.A(new_n1044), .B(KEYINPUT49), .Z(new_n1045));
  INV_X1    g0845(.A(new_n639), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n213), .B2(new_n806), .C1(new_n804), .C2(new_n796), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1039), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n784), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n771), .B1(new_n727), .B2(new_n783), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n259), .A2(G50), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  AOI21_X1  g0853(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1053), .A2(new_n740), .A3(new_n1054), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n776), .B(new_n1055), .C1(new_n237), .C2(new_n516), .ZN(new_n1056));
  OAI221_X1 g0856(.A(new_n1056), .B1(G107), .B2(new_n204), .C1(new_n740), .C2(new_n779), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1051), .B1(new_n786), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n1005), .B2(new_n993), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1032), .A2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n999), .A2(new_n1002), .ZN(new_n1061));
  XOR2_X1   g0861(.A(new_n1061), .B(new_n729), .Z(new_n1062));
  NAND2_X1  g0862(.A1(new_n1062), .A2(new_n1031), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1063), .A2(new_n737), .A3(new_n1010), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n993), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1062), .A2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n771), .B1(new_n1014), .B2(new_n783), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n803), .A2(new_n977), .B1(new_n792), .B2(new_n812), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI22_X1  g0869(.A1(new_n810), .A2(new_n815), .B1(new_n811), .B2(new_n799), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n800), .A2(new_n213), .ZN(new_n1071));
  NOR3_X1   g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n847), .A2(G283), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n281), .B1(new_n862), .B2(G107), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n797), .A2(G322), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n816), .A2(new_n222), .B1(new_n806), .B2(new_n470), .ZN(new_n1077));
  AOI211_X1 g0877(.A(new_n1077), .B(new_n1046), .C1(G143), .C2(new_n797), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT113), .Z(new_n1079));
  OAI22_X1  g0879(.A1(new_n803), .A2(new_n263), .B1(new_n792), .B2(new_n818), .ZN(new_n1080));
  XOR2_X1   g0880(.A(new_n1080), .B(KEYINPUT51), .Z(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(G50), .B2(new_n1040), .ZN(new_n1082));
  OAI211_X1 g0882(.A(new_n1079), .B(new_n1082), .C1(new_n207), .C2(new_n800), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n811), .A2(new_n259), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1076), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n784), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n776), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n785), .B1(new_n209), .B2(new_n204), .C1(new_n248), .C2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1067), .A2(new_n1086), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1064), .A2(new_n1066), .A3(new_n1089), .ZN(G390));
  AOI21_X1  g0890(.A(new_n771), .B1(new_n259), .B2(new_n845), .ZN(new_n1091));
  XOR2_X1   g0891(.A(new_n1091), .B(KEYINPUT115), .Z(new_n1092));
  OAI22_X1  g0892(.A1(new_n816), .A2(new_n470), .B1(new_n796), .B2(new_n799), .ZN(new_n1093));
  AOI211_X1 g0893(.A(new_n281), .B(new_n1093), .C1(G107), .C2(new_n1040), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n862), .A2(G68), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n793), .A2(G116), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n803), .A2(new_n807), .B1(new_n800), .B2(new_n207), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1097), .B1(G97), .B2(new_n856), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .A4(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(G125), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n796), .A2(new_n1100), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT54), .B(G143), .Z(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  INV_X1    g0903(.A(G128), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1103), .A2(new_n811), .B1(new_n1104), .B2(new_n803), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n1101), .B(new_n1105), .C1(G132), .C2(new_n793), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n281), .B1(new_n806), .B2(new_n256), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT116), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n847), .A2(new_n1034), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n1109), .A2(KEYINPUT53), .B1(new_n818), .B2(new_n800), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(KEYINPUT53), .B2(new_n1109), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1106), .A2(new_n1108), .A3(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n810), .A2(new_n858), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1099), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1092), .B1(new_n1114), .B2(new_n784), .ZN(new_n1115));
  XOR2_X1   g0915(.A(new_n1115), .B(KEYINPUT117), .Z(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n947), .B2(new_n782), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n836), .A2(new_n339), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n766), .A2(new_n731), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n931), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n900), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n919), .A2(new_n893), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n948), .B(KEYINPUT114), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n944), .B(new_n946), .C1(new_n938), .C2(new_n948), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n760), .A2(new_n837), .A3(new_n900), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1117), .B1(new_n1131), .B2(new_n1065), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1130), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1127), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n928), .A2(new_n871), .A3(new_n685), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n759), .A2(G330), .A3(new_n837), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n937), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1127), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1139), .A2(new_n932), .ZN(new_n1140));
  NAND4_X1  g0940(.A1(new_n1127), .A2(new_n931), .A3(new_n1119), .A4(new_n1138), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1136), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n738), .B1(new_n1135), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1142), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1131), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1132), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(G378));
  XOR2_X1   g0947(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n302), .A2(new_n306), .ZN(new_n1150));
  INV_X1    g0950(.A(KEYINPUT55), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n302), .A2(KEYINPUT55), .A3(new_n306), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n277), .A2(new_n879), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1152), .A2(new_n1153), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1154), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1149), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1157), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1159), .A2(new_n1148), .A3(new_n1155), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1158), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n903), .B2(new_n922), .ZN(new_n1163));
  INV_X1    g0963(.A(G330), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT105), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT38), .B1(new_n891), .B2(new_n892), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1165), .B1(new_n905), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n889), .A2(new_n893), .A3(KEYINPUT105), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n914), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1164), .B1(new_n1169), .B2(new_n915), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1170), .A2(new_n925), .A3(new_n1161), .ZN(new_n1171));
  NAND4_X1  g0971(.A1(new_n1163), .A2(new_n949), .A3(new_n940), .A4(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1170), .A2(new_n925), .A3(new_n1161), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1161), .B1(new_n1170), .B2(new_n925), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n950), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1129), .A2(new_n1130), .A3(new_n1142), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1136), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1172), .A2(new_n1175), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n738), .B1(new_n1178), .B2(KEYINPUT57), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1172), .A2(new_n1175), .A3(KEYINPUT119), .ZN(new_n1180));
  AOI21_X1  g0980(.A(KEYINPUT119), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1136), .B1(new_n1135), .B2(new_n1182), .ZN(new_n1183));
  NOR3_X1   g0983(.A1(new_n1180), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1179), .B1(new_n1184), .B2(KEYINPUT57), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1162), .A2(new_n781), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(G77), .A2(new_n847), .B1(new_n1040), .B2(G97), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n1187), .B1(new_n217), .B2(new_n806), .C1(new_n219), .C2(new_n792), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(new_n811), .A2(new_n313), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n796), .A2(new_n807), .ZN(new_n1190));
  NOR4_X1   g0990(.A1(new_n1188), .A2(new_n969), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n966), .A2(G116), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1191), .A2(new_n503), .A3(new_n1046), .A4(new_n1192), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT58), .Z(new_n1194));
  OAI22_X1  g0994(.A1(new_n803), .A2(new_n1100), .B1(new_n800), .B2(new_n263), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(G132), .A2(new_n1040), .B1(new_n856), .B2(G137), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1196), .B1(new_n1104), .B2(new_n792), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1195), .B(new_n1197), .C1(new_n847), .C2(new_n1102), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT59), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G33), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(G41), .B1(new_n797), .B2(G124), .ZN(new_n1201));
  OAI211_X1 g1001(.A(new_n1200), .B(new_n1201), .C1(new_n818), .C2(new_n806), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n414), .ZN(new_n1204));
  AOI21_X1  g1004(.A(G41), .B1(new_n1204), .B2(KEYINPUT3), .ZN(new_n1205));
  OAI22_X1  g1005(.A1(new_n1202), .A2(new_n1203), .B1(G50), .B2(new_n1205), .ZN(new_n1206));
  OAI21_X1  g1006(.A(new_n784), .B1(new_n1194), .B2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n845), .A2(new_n256), .ZN(new_n1208));
  NAND4_X1  g1008(.A1(new_n1186), .A2(new_n772), .A3(new_n1207), .A4(new_n1208), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1210), .B1(new_n1211), .B2(new_n993), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1185), .A2(new_n1212), .ZN(G375));
  OAI22_X1  g1013(.A1(new_n803), .A2(new_n799), .B1(new_n811), .B2(new_n219), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G116), .B2(new_n1040), .ZN(new_n1215));
  XOR2_X1   g1015(.A(new_n1215), .B(KEYINPUT121), .Z(new_n1216));
  OAI22_X1  g1016(.A1(new_n313), .A2(new_n800), .B1(new_n796), .B2(new_n815), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1216), .A2(new_n281), .A3(new_n971), .A4(new_n1217), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n209), .B2(new_n816), .C1(new_n807), .C2(new_n792), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(new_n1219), .B(KEYINPUT122), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n816), .A2(new_n818), .B1(new_n796), .B2(new_n1104), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT123), .Z(new_n1222));
  NOR2_X1   g1022(.A1(new_n811), .A2(new_n263), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n792), .A2(new_n858), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n639), .B1(new_n217), .B2(new_n806), .C1(new_n854), .C2(new_n803), .ZN(new_n1225));
  NOR4_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1224), .A4(new_n1225), .ZN(new_n1226));
  OAI221_X1 g1026(.A(new_n1226), .B1(new_n256), .B2(new_n800), .C1(new_n810), .C2(new_n1103), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n789), .B1(new_n1220), .B2(new_n1227), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n771), .B(new_n1228), .C1(new_n222), .C2(new_n845), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n900), .A2(new_n782), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT120), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1182), .A2(new_n993), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1140), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n1012), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1232), .B1(new_n1234), .B2(new_n1142), .ZN(G381));
  OR2_X1    g1035(.A1(G381), .A2(G384), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1185), .A2(new_n1146), .A3(new_n1212), .ZN(new_n1237));
  AND3_X1   g1037(.A1(new_n1064), .A2(new_n1066), .A3(new_n1089), .ZN(new_n1238));
  OAI211_X1 g1038(.A(new_n1238), .B(new_n992), .C1(new_n1013), .C2(new_n1028), .ZN(new_n1239));
  NAND3_X1  g1039(.A1(new_n1032), .A2(new_n832), .A3(new_n1059), .ZN(new_n1240));
  OR4_X1    g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1239), .A4(new_n1240), .ZN(G407));
  OAI211_X1 g1041(.A(G407), .B(G213), .C1(G343), .C2(new_n1237), .ZN(G409));
  NAND2_X1  g1042(.A1(G387), .A2(G390), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1244), .A2(new_n1240), .ZN(new_n1245));
  XOR2_X1   g1045(.A(new_n1245), .B(KEYINPUT125), .Z(new_n1246));
  AND3_X1   g1046(.A1(new_n1239), .A2(new_n1243), .A3(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1246), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(new_n1146), .B1(new_n1185), .B2(new_n1212), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT119), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n950), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1252));
  AOI22_X1  g1052(.A1(new_n1163), .A2(new_n1171), .B1(new_n949), .B2(new_n940), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1251), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1176), .A2(new_n1177), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1172), .A2(new_n1175), .A3(KEYINPUT119), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1254), .A2(new_n1012), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n993), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1258));
  INV_X1    g1058(.A(KEYINPUT124), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(new_n1209), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1065), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1261));
  OAI21_X1  g1061(.A(KEYINPUT124), .B1(new_n1261), .B2(new_n1210), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1257), .A2(new_n1260), .A3(new_n1146), .A4(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n720), .A2(G213), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(KEYINPUT126), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1172), .A2(new_n1175), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1267), .A2(new_n1255), .A3(KEYINPUT57), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1268), .A2(new_n737), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT57), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1254), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1269), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1209), .B1(new_n1273), .B2(new_n1065), .ZN(new_n1274));
  OAI21_X1  g1074(.A(G378), .B1(new_n1272), .B2(new_n1274), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT126), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1275), .A2(new_n1276), .A3(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1266), .A2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT60), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n738), .B1(new_n1233), .B2(new_n1280), .ZN(new_n1281));
  OAI211_X1 g1081(.A(new_n1281), .B(new_n1144), .C1(new_n1280), .C2(new_n1233), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1232), .ZN(new_n1283));
  INV_X1    g1083(.A(G384), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1282), .A2(G384), .A3(new_n1232), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1285), .A2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1287), .ZN(new_n1290));
  NAND3_X1  g1090(.A1(new_n1275), .A2(new_n1276), .A3(new_n1290), .ZN(new_n1291));
  AOI22_X1  g1091(.A1(new_n1279), .A2(new_n1289), .B1(new_n1288), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n720), .A2(G213), .A3(G2897), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1287), .B(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1266), .A2(new_n1278), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  OAI21_X1  g1097(.A(new_n1249), .B1(new_n1292), .B2(new_n1297), .ZN(new_n1298));
  AND2_X1   g1098(.A1(new_n1290), .A2(KEYINPUT63), .ZN(new_n1299));
  NOR3_X1   g1099(.A1(new_n1250), .A2(KEYINPUT126), .A3(new_n1265), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1277), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT127), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT127), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1279), .A2(new_n1304), .A3(new_n1299), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1296), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1294), .B1(new_n1250), .B2(new_n1265), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(KEYINPUT63), .ZN(new_n1308));
  AOI21_X1  g1108(.A(new_n1306), .B1(new_n1308), .B2(new_n1291), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1303), .A2(new_n1305), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1298), .A2(new_n1310), .ZN(G405));
  NAND2_X1  g1111(.A1(new_n1275), .A2(new_n1237), .ZN(new_n1312));
  XNOR2_X1  g1112(.A(new_n1312), .B(new_n1287), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(new_n1313), .B(new_n1249), .ZN(G402));
endmodule


