//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:11 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n634, new_n635, new_n637, new_n638, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n854, new_n855, new_n856, new_n857,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT64), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n452), .B(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT66), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  OR2_X1    g034(.A1(new_n454), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n455), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G567), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n466), .A2(new_n467), .A3(G101), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(KEYINPUT3), .B(G2104), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(G137), .A3(new_n469), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  OAI21_X1  g052(.A(G125), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n469), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n475), .A2(new_n480), .ZN(G160));
  INV_X1    g056(.A(new_n477), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(G2105), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n469), .B1(new_n482), .B2(new_n483), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G124), .ZN(new_n487));
  OR2_X1    g062(.A1(G100), .A2(G2105), .ZN(new_n488));
  OAI211_X1 g063(.A(new_n488), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n485), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(new_n490), .ZN(G162));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n476), .C2(new_n477), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(G138), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G2105), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n499), .B1(new_n476), .B2(new_n477), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT4), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT4), .ZN(new_n502));
  OAI211_X1 g077(.A(new_n499), .B(new_n502), .C1(new_n477), .C2(new_n476), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n497), .B1(new_n501), .B2(new_n503), .ZN(G164));
  AND2_X1   g079(.A1(KEYINPUT5), .A2(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT5), .A2(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G62), .ZN(new_n508));
  INV_X1    g083(.A(G75), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(G88), .B1(new_n505), .B2(new_n506), .ZN(new_n512));
  NAND2_X1  g087(.A1(G50), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g089(.A(G651), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(KEYINPUT6), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT68), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n518), .B2(G651), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n515), .A2(KEYINPUT68), .A3(KEYINPUT6), .ZN(new_n520));
  AOI21_X1  g095(.A(new_n516), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n511), .A2(G651), .B1(new_n514), .B2(new_n521), .ZN(G166));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  OAI21_X1  g098(.A(G543), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AOI211_X1 g099(.A(KEYINPUT69), .B(new_n516), .C1(new_n519), .C2(new_n520), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G51), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT70), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT7), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n529), .B(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(KEYINPUT5), .A2(G543), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n521), .A2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n534), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n527), .A2(new_n531), .A3(new_n537), .A4(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  NAND2_X1  g115(.A1(new_n526), .A2(G52), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G64), .ZN(new_n543));
  OAI21_X1  g118(.A(new_n542), .B1(new_n507), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n536), .A2(G90), .B1(G651), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n541), .A2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  NAND2_X1  g122(.A1(new_n526), .A2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n507), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n536), .A2(G81), .B1(G651), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  NAND4_X1  g130(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND4_X1  g133(.A1(G319), .A2(G483), .A3(G661), .A4(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n519), .A2(new_n520), .ZN(new_n560));
  INV_X1    g135(.A(new_n516), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(KEYINPUT69), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n521), .A2(new_n523), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n563), .A2(G53), .A3(G543), .A4(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n565), .A2(KEYINPUT9), .ZN(new_n566));
  INV_X1    g141(.A(new_n524), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n567), .A2(new_n568), .A3(G53), .A4(new_n564), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n507), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  INV_X1    g149(.A(G91), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n575), .B2(new_n535), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT71), .B1(new_n570), .B2(new_n577), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT71), .ZN(new_n579));
  AOI211_X1 g154(.A(new_n579), .B(new_n576), .C1(new_n566), .C2(new_n569), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n578), .A2(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n514), .A2(new_n521), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n508), .B1(new_n532), .B2(new_n533), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n509), .A2(new_n510), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n582), .A2(new_n585), .ZN(G303));
  NAND3_X1  g161(.A1(new_n521), .A2(G87), .A3(new_n534), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n534), .B2(G74), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n589), .B1(new_n526), .B2(G49), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(G288));
  OAI21_X1  g166(.A(G61), .B1(new_n505), .B2(new_n506), .ZN(new_n592));
  NAND2_X1  g167(.A1(G73), .A2(G543), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n515), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT72), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n534), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n596));
  OAI22_X1  g171(.A1(new_n594), .A2(new_n595), .B1(new_n596), .B2(new_n562), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n592), .A2(new_n593), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(G651), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(KEYINPUT72), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(new_n601), .ZN(G305));
  AOI22_X1  g177(.A1(new_n534), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n603));
  NOR2_X1   g178(.A1(new_n603), .A2(new_n515), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT73), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n536), .A2(G85), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(new_n608));
  INV_X1    g183(.A(new_n526), .ZN(new_n609));
  XNOR2_X1  g184(.A(KEYINPUT74), .B(G47), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n608), .A2(new_n612), .ZN(G290));
  NAND2_X1  g188(.A1(G301), .A2(G868), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n521), .A2(G92), .A3(new_n534), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT10), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n526), .A2(G54), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n534), .A2(G66), .ZN(new_n618));
  NAND2_X1  g193(.A1(G79), .A2(G543), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT75), .ZN(new_n620));
  OAI21_X1  g195(.A(G651), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n616), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n614), .B1(new_n623), .B2(G868), .ZN(G284));
  OAI21_X1  g199(.A(new_n614), .B1(new_n623), .B2(G868), .ZN(G321));
  INV_X1    g200(.A(G868), .ZN(new_n626));
  NOR2_X1   g201(.A1(G286), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n570), .A2(new_n577), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(new_n579), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n570), .A2(KEYINPUT71), .A3(new_n577), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g206(.A(new_n627), .B1(new_n631), .B2(new_n626), .ZN(G297));
  AOI21_X1  g207(.A(new_n627), .B1(new_n631), .B2(new_n626), .ZN(G280));
  INV_X1    g208(.A(G860), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n622), .B1(G559), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT76), .ZN(G148));
  OR2_X1    g211(.A1(new_n622), .A2(G559), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(G868), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n638), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g214(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g215(.A1(new_n473), .A2(new_n466), .ZN(new_n641));
  XOR2_X1   g216(.A(KEYINPUT77), .B(KEYINPUT12), .Z(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT13), .ZN(new_n644));
  INV_X1    g219(.A(G2100), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n644), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n484), .A2(G135), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n486), .A2(G123), .ZN(new_n649));
  NOR2_X1   g224(.A1(new_n469), .A2(G111), .ZN(new_n650));
  OAI21_X1  g225(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n648), .B(new_n649), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  INV_X1    g227(.A(G2096), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n646), .A2(new_n647), .A3(new_n654), .ZN(G156));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2443), .B(G2446), .ZN(new_n657));
  XOR2_X1   g232(.A(new_n656), .B(new_n657), .Z(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(KEYINPUT15), .B(G2435), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(G2438), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2427), .B(G2430), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(KEYINPUT14), .ZN(new_n664));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n661), .A2(new_n662), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1341), .B(G1348), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n666), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n670), .B1(new_n666), .B2(new_n668), .ZN(new_n673));
  OAI21_X1  g248(.A(new_n659), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n666), .A2(new_n668), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n676), .A2(new_n658), .A3(new_n671), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT78), .B(KEYINPUT16), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n674), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n679), .A2(G14), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n678), .B1(new_n674), .B2(new_n677), .ZN(new_n681));
  OAI21_X1  g256(.A(KEYINPUT80), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n674), .A2(new_n677), .ZN(new_n683));
  INV_X1    g258(.A(new_n678), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT80), .ZN(new_n686));
  NAND4_X1  g261(.A1(new_n685), .A2(new_n686), .A3(G14), .A4(new_n679), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n682), .A2(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(G401));
  INV_X1    g264(.A(KEYINPUT18), .ZN(new_n690));
  XOR2_X1   g265(.A(G2084), .B(G2090), .Z(new_n691));
  XNOR2_X1  g266(.A(G2067), .B(G2678), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(KEYINPUT17), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n691), .A2(new_n692), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n696), .B(new_n645), .ZN(new_n697));
  XOR2_X1   g272(.A(G2072), .B(G2078), .Z(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n693), .B2(KEYINPUT18), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(new_n653), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n697), .B(new_n700), .ZN(G227));
  XNOR2_X1  g276(.A(G1971), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(KEYINPUT81), .B(KEYINPUT19), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1956), .B(G2474), .ZN(new_n705));
  XNOR2_X1  g280(.A(G1961), .B(G1966), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n704), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n705), .B(new_n706), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n705), .A2(new_n706), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  AND2_X1   g285(.A1(new_n710), .A2(KEYINPUT20), .ZN(new_n711));
  NOR2_X1   g286(.A1(new_n710), .A2(KEYINPUT20), .ZN(new_n712));
  OAI221_X1 g287(.A(new_n707), .B1(new_n704), .B2(new_n708), .C1(new_n711), .C2(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(G1991), .B(G1996), .Z(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(G1981), .B(G1986), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n717), .B(new_n718), .ZN(G229));
  INV_X1    g294(.A(G16), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G24), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT83), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G290), .B2(G16), .ZN(new_n723));
  INV_X1    g298(.A(G1986), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n723), .A2(new_n724), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n484), .A2(G131), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n486), .A2(G119), .ZN(new_n728));
  NOR2_X1   g303(.A1(new_n469), .A2(G107), .ZN(new_n729));
  OAI21_X1  g304(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n730), .ZN(new_n731));
  MUX2_X1   g306(.A(G25), .B(new_n731), .S(G29), .Z(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT82), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n732), .B(new_n734), .ZN(new_n735));
  NOR3_X1   g310(.A1(new_n725), .A2(new_n726), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n601), .A2(G16), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G6), .B2(G16), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT32), .B(G1981), .Z(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n738), .A2(new_n739), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n720), .A2(G22), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G166), .B2(new_n720), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(G1971), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(G1971), .ZN(new_n745));
  NAND4_X1  g320(.A1(new_n740), .A2(new_n741), .A3(new_n744), .A4(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n720), .A2(G23), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(new_n590), .B2(new_n720), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT33), .B(G1976), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n746), .A2(KEYINPUT34), .A3(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(KEYINPUT34), .B1(new_n746), .B2(new_n750), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n736), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(KEYINPUT84), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n754), .A2(KEYINPUT36), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT85), .Z(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n753), .A2(new_n757), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n623), .A2(G16), .ZN(new_n761));
  OAI211_X1 g336(.A(new_n761), .B(G1348), .C1(G4), .C2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  NOR2_X1   g338(.A1(G164), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G27), .B2(new_n763), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(G2078), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(G2078), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n765), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n770), .A2(KEYINPUT94), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n763), .A2(G33), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT88), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT25), .ZN(new_n775));
  AND2_X1   g350(.A1(new_n473), .A2(G127), .ZN(new_n776));
  AND2_X1   g351(.A1(G115), .A2(G2104), .ZN(new_n777));
  OAI21_X1  g352(.A(G2105), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(KEYINPUT89), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n484), .A2(G139), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n778), .B2(KEYINPUT89), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n772), .B1(new_n783), .B2(new_n763), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n784), .A2(G2072), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n762), .A2(new_n768), .A3(new_n771), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n763), .B1(KEYINPUT24), .B2(G34), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(KEYINPUT24), .B2(G34), .ZN(new_n788));
  INV_X1    g363(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G160), .B2(new_n763), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n790), .A2(G2084), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(KEYINPUT93), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n763), .A2(G35), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G162), .B2(new_n763), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT29), .B(G2090), .Z(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n792), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(new_n784), .A2(G2072), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n763), .A2(G26), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT28), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n484), .A2(G140), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n486), .A2(G128), .ZN(new_n802));
  OR2_X1    g377(.A1(G104), .A2(G2105), .ZN(new_n803));
  OAI211_X1 g378(.A(new_n803), .B(G2104), .C1(G116), .C2(new_n469), .ZN(new_n804));
  NAND3_X1  g379(.A1(new_n801), .A2(new_n802), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n805), .A2(G29), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(KEYINPUT87), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(KEYINPUT87), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n800), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(G2067), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n809), .B(new_n810), .ZN(new_n811));
  AND2_X1   g386(.A1(new_n763), .A2(G32), .ZN(new_n812));
  AOI22_X1  g387(.A1(new_n484), .A2(G141), .B1(G105), .B2(new_n466), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n486), .A2(G129), .ZN(new_n814));
  NAND3_X1  g389(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(KEYINPUT26), .Z(new_n816));
  NAND3_X1  g391(.A1(new_n813), .A2(new_n814), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g392(.A(new_n812), .B1(new_n817), .B2(G29), .ZN(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT27), .B(G1996), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT30), .B(G28), .ZN(new_n821));
  OR2_X1    g396(.A1(KEYINPUT31), .A2(G11), .ZN(new_n822));
  NAND2_X1  g397(.A1(KEYINPUT31), .A2(G11), .ZN(new_n823));
  AOI22_X1  g398(.A1(new_n821), .A2(new_n763), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n652), .B2(new_n763), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(new_n818), .B2(new_n819), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n790), .A2(G2084), .ZN(new_n827));
  AND3_X1   g402(.A1(new_n820), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n797), .A2(new_n798), .A3(new_n811), .A4(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(G1961), .ZN(new_n830));
  NOR2_X1   g405(.A1(G5), .A2(G16), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT90), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G301), .B2(new_n720), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT91), .ZN(new_n834));
  AOI211_X1 g409(.A(new_n786), .B(new_n829), .C1(new_n830), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n720), .A2(G20), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT23), .ZN(new_n837));
  OAI21_X1  g412(.A(new_n837), .B1(new_n631), .B2(new_n720), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(G1956), .Z(new_n839));
  NOR2_X1   g414(.A1(new_n834), .A2(new_n830), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT92), .Z(new_n841));
  NOR2_X1   g416(.A1(G16), .A2(G19), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n842), .B1(new_n554), .B2(G16), .ZN(new_n843));
  XOR2_X1   g418(.A(KEYINPUT86), .B(G1341), .Z(new_n844));
  XNOR2_X1  g419(.A(new_n843), .B(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n720), .A2(G21), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n846), .B1(G168), .B2(new_n720), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G1966), .ZN(new_n848));
  INV_X1    g423(.A(G1348), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n761), .B1(G4), .B2(G16), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n845), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n835), .A2(new_n839), .A3(new_n841), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n760), .A2(new_n852), .ZN(G311));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT95), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n854), .A2(new_n855), .A3(new_n758), .A4(new_n759), .ZN(new_n856));
  OAI21_X1  g431(.A(KEYINPUT95), .B1(new_n760), .B2(new_n852), .ZN(new_n857));
  AND2_X1   g432(.A1(new_n856), .A2(new_n857), .ZN(G150));
  NAND2_X1  g433(.A1(new_n623), .A2(G559), .ZN(new_n859));
  XOR2_X1   g434(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(G80), .A2(G543), .ZN(new_n862));
  INV_X1    g437(.A(G67), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n862), .B1(new_n507), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g439(.A1(new_n864), .A2(KEYINPUT97), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n515), .B1(new_n864), .B2(KEYINPUT97), .ZN(new_n866));
  AOI22_X1  g441(.A1(new_n865), .A2(new_n866), .B1(G93), .B2(new_n536), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n526), .A2(G55), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(new_n553), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n553), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(new_n861), .B(new_n872), .Z(new_n873));
  OR2_X1    g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n874), .A2(new_n634), .A3(new_n875), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n869), .A2(G860), .ZN(new_n877));
  XOR2_X1   g452(.A(new_n877), .B(KEYINPUT37), .Z(new_n878));
  NAND2_X1  g453(.A1(new_n876), .A2(new_n878), .ZN(G145));
  INV_X1    g454(.A(KEYINPUT98), .ZN(new_n880));
  XOR2_X1   g455(.A(G164), .B(new_n805), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n484), .A2(G142), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n486), .A2(G130), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n469), .A2(G118), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n885));
  OAI211_X1 g460(.A(new_n882), .B(new_n883), .C1(new_n884), .C2(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n881), .B(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n817), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n783), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n817), .B1(new_n780), .B2(new_n782), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n731), .B(new_n643), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n890), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n893), .B1(new_n890), .B2(new_n891), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n888), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(new_n896), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n898), .A2(new_n887), .A3(new_n894), .ZN(new_n899));
  XOR2_X1   g474(.A(G160), .B(new_n652), .Z(new_n900));
  XNOR2_X1  g475(.A(new_n900), .B(new_n490), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n897), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(G37), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n901), .B1(new_n897), .B2(new_n899), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n880), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n905), .ZN(new_n907));
  NAND4_X1  g482(.A1(new_n907), .A2(KEYINPUT98), .A3(new_n903), .A4(new_n902), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g485(.A1(G290), .A2(new_n601), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n607), .A2(new_n601), .A3(new_n611), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(new_n590), .B(G166), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT100), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n917));
  INV_X1    g492(.A(new_n914), .ZN(new_n918));
  AOI21_X1  g493(.A(G305), .B1(new_n608), .B2(new_n612), .ZN(new_n919));
  OAI21_X1  g494(.A(new_n918), .B1(new_n919), .B2(new_n912), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n915), .A2(new_n917), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n921), .A2(KEYINPUT101), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT101), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n915), .A2(new_n920), .A3(new_n923), .A4(new_n917), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n916), .A2(KEYINPUT42), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n922), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g502(.A(new_n926), .B1(new_n922), .B2(new_n924), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n631), .A2(new_n622), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT99), .ZN(new_n931));
  AOI21_X1  g506(.A(new_n931), .B1(G299), .B2(new_n623), .ZN(new_n932));
  NOR4_X1   g507(.A1(new_n578), .A2(new_n580), .A3(KEYINPUT99), .A4(new_n622), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  XNOR2_X1  g509(.A(new_n872), .B(new_n637), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(G299), .A2(new_n623), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n930), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT41), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n939), .B1(new_n631), .B2(new_n622), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n941), .B1(new_n932), .B2(new_n933), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n935), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(new_n929), .A2(new_n936), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n943), .A2(new_n936), .ZN(new_n945));
  NOR3_X1   g520(.A1(new_n945), .A2(new_n927), .A3(new_n928), .ZN(new_n946));
  OAI21_X1  g521(.A(G868), .B1(new_n944), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n869), .A2(new_n626), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n947), .A2(new_n948), .ZN(G295));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n948), .ZN(G331));
  INV_X1    g525(.A(KEYINPUT43), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT102), .ZN(new_n952));
  NAND2_X1  g527(.A1(G301), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n541), .A2(KEYINPUT102), .A3(new_n545), .ZN(new_n954));
  AND3_X1   g529(.A1(new_n953), .A2(G286), .A3(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G286), .B1(new_n953), .B2(new_n954), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n872), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(new_n954), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT102), .B1(new_n541), .B2(new_n545), .ZN(new_n959));
  OAI21_X1  g534(.A(G168), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n953), .A2(G286), .A3(new_n954), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n871), .A3(new_n961), .A4(new_n870), .ZN(new_n962));
  AND2_X1   g537(.A1(new_n957), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n940), .A2(new_n942), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n915), .A2(new_n920), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n957), .A2(new_n962), .ZN(new_n967));
  OAI211_X1 g542(.A(new_n967), .B(new_n930), .C1(new_n932), .C2(new_n933), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n903), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n966), .B1(new_n964), .B2(new_n968), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n951), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n967), .A2(new_n939), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n965), .B1(new_n973), .B2(new_n938), .ZN(new_n974));
  OAI221_X1 g549(.A(new_n930), .B1(new_n932), .B2(new_n933), .C1(new_n967), .C2(new_n939), .ZN(new_n975));
  AOI21_X1  g550(.A(G37), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n964), .A2(new_n968), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n976), .B1(new_n966), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n972), .B1(new_n978), .B2(new_n951), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(KEYINPUT44), .ZN(new_n980));
  OAI21_X1  g555(.A(KEYINPUT43), .B1(new_n970), .B2(new_n971), .ZN(new_n981));
  OAI211_X1 g556(.A(new_n976), .B(new_n951), .C1(new_n966), .C2(new_n977), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n980), .A2(new_n985), .ZN(G397));
  INV_X1    g561(.A(KEYINPUT55), .ZN(new_n987));
  INV_X1    g562(.A(G8), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(G166), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT45), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n993), .B1(G164), .B2(G1384), .ZN(new_n994));
  INV_X1    g569(.A(G40), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n475), .A2(new_n480), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1384), .ZN(new_n997));
  INV_X1    g572(.A(new_n503), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n502), .B1(new_n473), .B2(new_n499), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(KEYINPUT45), .B(new_n997), .C1(new_n1000), .C2(new_n497), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n994), .A2(new_n996), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(G1971), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT50), .ZN(new_n1006));
  OAI211_X1 g581(.A(new_n1006), .B(new_n997), .C1(new_n1000), .C2(new_n497), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT112), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n501), .A2(new_n503), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n492), .A2(new_n496), .ZN(new_n1011));
  AOI21_X1  g586(.A(G1384), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1012), .A2(KEYINPUT112), .A3(new_n1006), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1009), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n996), .B1(new_n1012), .B2(new_n1006), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  OAI211_X1 g592(.A(new_n996), .B(KEYINPUT111), .C1(new_n1012), .C2(new_n1006), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G2090), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1005), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT108), .B(G8), .Z(new_n1022));
  OAI21_X1  g597(.A(new_n992), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n1024), .A2(new_n1007), .A3(new_n1020), .A4(new_n996), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1004), .A2(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT107), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n989), .A2(new_n1027), .A3(new_n990), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1027), .B1(new_n989), .B2(new_n990), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1026), .A2(new_n1030), .A3(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n567), .A2(G49), .A3(new_n564), .ZN(new_n1033));
  INV_X1    g608(.A(new_n589), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(new_n1034), .A3(G1976), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1022), .B1(new_n996), .B2(new_n1012), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1032), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(new_n1022), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n997), .B1(new_n1000), .B2(new_n497), .ZN(new_n1039));
  INV_X1    g614(.A(new_n480), .ZN(new_n1040));
  NAND4_X1  g615(.A1(new_n1040), .A2(G40), .A3(new_n474), .A4(new_n472), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1038), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(G1981), .B1(new_n597), .B2(new_n600), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n599), .A2(KEYINPUT72), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n594), .A2(new_n595), .ZN(new_n1045));
  NAND2_X1  g620(.A1(G48), .A2(G543), .ZN(new_n1046));
  INV_X1    g621(.A(G86), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n507), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n521), .ZN(new_n1049));
  XNOR2_X1  g624(.A(KEYINPUT110), .B(G1981), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1044), .A2(new_n1045), .A3(new_n1049), .A4(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT49), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1043), .A2(KEYINPUT49), .A3(new_n1051), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1037), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1032), .B1(new_n590), .B2(G1976), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(KEYINPUT109), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT109), .ZN(new_n1059));
  OAI211_X1 g634(.A(new_n1059), .B(new_n1032), .C1(new_n590), .C2(G1976), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1058), .A2(new_n1060), .A3(new_n1036), .A4(new_n1035), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1031), .A2(new_n1056), .A3(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT122), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1023), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(G1966), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1002), .A2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G2084), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1024), .A2(new_n1007), .A3(new_n1067), .A4(new_n996), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n988), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g644(.A1(G168), .A2(new_n1022), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT51), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(G286), .B2(new_n1038), .ZN(new_n1072));
  AOI21_X1  g647(.A(new_n1022), .B1(new_n1066), .B2(new_n1068), .ZN(new_n1073));
  OAI21_X1  g648(.A(new_n1072), .B1(new_n1073), .B2(KEYINPUT119), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1066), .A2(new_n1068), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1075), .A2(KEYINPUT119), .A3(new_n1038), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1074), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1075), .A2(new_n1070), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NOR4_X1   g654(.A1(G164), .A2(new_n1008), .A3(KEYINPUT50), .A4(G1384), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT112), .B1(new_n1012), .B2(new_n1006), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT111), .B1(new_n1024), .B2(new_n996), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1018), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n1082), .B(new_n1020), .C1(new_n1083), .C2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n1004), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n991), .B1(new_n1086), .B2(new_n1038), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1031), .A2(new_n1056), .A3(new_n1061), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT122), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT53), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n994), .A2(new_n1001), .A3(new_n769), .A4(new_n996), .ZN(new_n1091));
  AOI21_X1  g666(.A(G171), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NOR3_X1   g667(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1093));
  OAI21_X1  g668(.A(KEYINPUT113), .B1(new_n1015), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT113), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1024), .A2(new_n1007), .A3(new_n1095), .A4(new_n996), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1094), .A2(new_n830), .A3(new_n1096), .ZN(new_n1097));
  AND2_X1   g672(.A1(new_n994), .A2(new_n1001), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1098), .A2(KEYINPUT53), .A3(new_n769), .A4(new_n996), .ZN(new_n1099));
  AND3_X1   g674(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(KEYINPUT120), .B1(new_n1097), .B2(new_n1099), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1092), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1091), .A2(new_n1090), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n769), .A2(KEYINPUT53), .A3(G40), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT121), .B1(new_n478), .B2(new_n479), .ZN(new_n1106));
  NOR2_X1   g681(.A1(new_n1106), .A2(new_n469), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n478), .A2(KEYINPUT121), .A3(new_n479), .ZN(new_n1108));
  AOI211_X1 g683(.A(new_n1105), .B(new_n475), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1098), .A2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1097), .A2(new_n1104), .A3(new_n1110), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1103), .B1(new_n1111), .B2(G171), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1102), .A2(new_n1112), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1064), .A2(new_n1079), .A3(new_n1089), .A4(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1104), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1115), .A2(G171), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1111), .A2(G171), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT54), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT123), .B1(new_n1114), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT120), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1097), .A2(KEYINPUT120), .A3(new_n1099), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1125), .B2(new_n1104), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1103), .B1(new_n1126), .B2(new_n1117), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1063), .B1(new_n1023), .B2(new_n1062), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1087), .A2(new_n1088), .A3(KEYINPUT122), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT123), .ZN(new_n1131));
  AOI22_X1  g706(.A1(new_n1077), .A2(new_n1078), .B1(new_n1102), .B2(new_n1112), .ZN(new_n1132));
  NAND4_X1  g707(.A1(new_n1127), .A2(new_n1130), .A3(new_n1131), .A4(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT57), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1134), .B1(new_n570), .B2(new_n577), .ZN(new_n1135));
  AOI211_X1 g710(.A(KEYINPUT57), .B(new_n576), .C1(new_n566), .C2(new_n569), .ZN(new_n1136));
  OR2_X1    g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1138));
  AOI21_X1  g713(.A(G1956), .B1(new_n1138), .B2(new_n1082), .ZN(new_n1139));
  XOR2_X1   g714(.A(KEYINPUT56), .B(G2072), .Z(new_n1140));
  NOR2_X1   g715(.A1(new_n1002), .A2(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1141), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1143), .B(new_n1144), .C1(new_n1019), .C2(G1956), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1142), .A2(new_n1145), .A3(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT61), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1144), .B1(new_n1019), .B2(G1956), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1149), .A2(KEYINPUT117), .A3(new_n1137), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1147), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1148), .B1(new_n1149), .B2(new_n1137), .ZN(new_n1152));
  XOR2_X1   g727(.A(KEYINPUT58), .B(G1341), .Z(new_n1153));
  OAI21_X1  g728(.A(new_n1153), .B1(new_n1039), .B2(new_n1041), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(KEYINPUT116), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT116), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1156), .B(new_n1153), .C1(new_n1039), .C2(new_n1041), .ZN(new_n1157));
  OAI211_X1 g732(.A(new_n1155), .B(new_n1157), .C1(G1996), .C2(new_n1002), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n554), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(KEYINPUT59), .ZN(new_n1160));
  INV_X1    g735(.A(KEYINPUT59), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1158), .A2(new_n1161), .A3(new_n554), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1152), .A2(new_n1145), .B1(new_n1160), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1094), .A2(new_n849), .A3(new_n1096), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n996), .A2(new_n1012), .A3(new_n810), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(KEYINPUT60), .B1(new_n622), .B2(KEYINPUT118), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n622), .A2(KEYINPUT118), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT60), .ZN(new_n1171));
  AOI22_X1  g746(.A1(new_n1166), .A2(new_n1171), .B1(KEYINPUT118), .B2(new_n622), .ZN(new_n1172));
  OAI21_X1  g747(.A(new_n1170), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1151), .A2(new_n1163), .A3(new_n1173), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1166), .A2(KEYINPUT114), .A3(new_n623), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1142), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(KEYINPUT114), .B1(new_n1166), .B2(new_n623), .ZN(new_n1177));
  OAI211_X1 g752(.A(KEYINPUT115), .B(new_n1145), .C1(new_n1176), .C2(new_n1177), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1145), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT115), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1174), .A2(new_n1178), .A3(new_n1181), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1120), .A2(new_n1133), .A3(new_n1182), .ZN(new_n1183));
  AND3_X1   g758(.A1(new_n1073), .A2(KEYINPUT63), .A3(G168), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n988), .B1(new_n1004), .B2(new_n1025), .ZN(new_n1185));
  OAI211_X1 g760(.A(new_n1062), .B(new_n1184), .C1(new_n991), .C2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1073), .A2(G168), .ZN(new_n1187));
  NOR3_X1   g762(.A1(new_n1087), .A2(new_n1088), .A3(new_n1187), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1186), .B1(new_n1188), .B2(KEYINPUT63), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1190), .ZN(new_n1191));
  OR2_X1    g766(.A1(G288), .A2(G1976), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n1051), .B1(new_n1191), .B2(new_n1192), .ZN(new_n1193));
  AND2_X1   g768(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1194));
  INV_X1    g769(.A(new_n1031), .ZN(new_n1195));
  AOI22_X1  g770(.A1(new_n1036), .A2(new_n1193), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1189), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g772(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1198));
  NOR3_X1   g773(.A1(new_n1198), .A2(new_n1128), .A3(new_n1129), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1116), .B1(new_n1079), .B2(KEYINPUT62), .ZN(new_n1200));
  AOI21_X1  g775(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1183), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g777(.A1(new_n608), .A2(new_n724), .A3(new_n612), .ZN(new_n1203));
  AND2_X1   g778(.A1(new_n1203), .A2(KEYINPUT103), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n994), .A2(new_n1041), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1205), .B1(new_n1203), .B2(KEYINPUT103), .ZN(new_n1206));
  OR2_X1    g781(.A1(new_n1204), .A2(new_n1206), .ZN(new_n1207));
  NAND3_X1  g782(.A1(G290), .A2(G1986), .A3(new_n1205), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  XOR2_X1   g784(.A(new_n1209), .B(KEYINPUT104), .Z(new_n1210));
  XNOR2_X1  g785(.A(new_n805), .B(new_n810), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n817), .A2(G1996), .ZN(new_n1212));
  INV_X1    g787(.A(G1996), .ZN(new_n1213));
  NAND2_X1  g788(.A1(new_n889), .A2(new_n1213), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1211), .A2(new_n1212), .A3(new_n1214), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1215), .A2(new_n1205), .ZN(new_n1216));
  XNOR2_X1  g791(.A(new_n1216), .B(KEYINPUT105), .ZN(new_n1217));
  INV_X1    g792(.A(new_n733), .ZN(new_n1218));
  XNOR2_X1  g793(.A(new_n731), .B(new_n1218), .ZN(new_n1219));
  INV_X1    g794(.A(KEYINPUT106), .ZN(new_n1220));
  OR2_X1    g795(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1219), .A2(new_n1220), .ZN(new_n1222));
  NAND3_X1  g797(.A1(new_n1221), .A2(new_n1205), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1217), .A2(new_n1223), .ZN(new_n1224));
  NOR2_X1   g799(.A1(new_n1210), .A2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1202), .A2(new_n1225), .ZN(new_n1226));
  INV_X1    g801(.A(KEYINPUT48), .ZN(new_n1227));
  OR2_X1    g802(.A1(new_n1207), .A2(new_n1227), .ZN(new_n1228));
  AOI21_X1  g803(.A(new_n1224), .B1(new_n1207), .B2(new_n1227), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g805(.A1(new_n731), .A2(new_n1218), .ZN(new_n1231));
  NAND2_X1  g806(.A1(new_n1217), .A2(new_n1231), .ZN(new_n1232));
  OR2_X1    g807(.A1(new_n805), .A2(G2067), .ZN(new_n1233));
  NAND2_X1  g808(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1234), .A2(new_n1205), .ZN(new_n1235));
  OAI21_X1  g810(.A(new_n1230), .B1(KEYINPUT124), .B2(new_n1235), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1235), .A2(KEYINPUT124), .ZN(new_n1237));
  NAND2_X1  g812(.A1(new_n1205), .A2(new_n1213), .ZN(new_n1238));
  XNOR2_X1  g813(.A(new_n1238), .B(KEYINPUT46), .ZN(new_n1239));
  NAND2_X1  g814(.A1(new_n1211), .A2(new_n889), .ZN(new_n1240));
  NAND2_X1  g815(.A1(new_n1240), .A2(new_n1205), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1239), .A2(new_n1241), .ZN(new_n1242));
  XNOR2_X1  g817(.A(new_n1242), .B(KEYINPUT47), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1237), .A2(new_n1243), .ZN(new_n1244));
  OAI21_X1  g819(.A(KEYINPUT125), .B1(new_n1236), .B2(new_n1244), .ZN(new_n1245));
  INV_X1    g820(.A(new_n1235), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT124), .ZN(new_n1247));
  AOI22_X1  g822(.A1(new_n1246), .A2(new_n1247), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1248));
  INV_X1    g823(.A(KEYINPUT125), .ZN(new_n1249));
  NAND4_X1  g824(.A1(new_n1248), .A2(new_n1249), .A3(new_n1237), .A4(new_n1243), .ZN(new_n1250));
  NAND2_X1  g825(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g826(.A1(new_n1226), .A2(new_n1251), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g827(.A(G229), .B1(new_n906), .B2(new_n908), .ZN(new_n1254));
  NOR2_X1   g828(.A1(G227), .A2(new_n463), .ZN(new_n1255));
  AOI21_X1  g829(.A(KEYINPUT126), .B1(new_n688), .B2(new_n1255), .ZN(new_n1256));
  INV_X1    g830(.A(KEYINPUT126), .ZN(new_n1257));
  INV_X1    g831(.A(new_n1255), .ZN(new_n1258));
  AOI211_X1 g832(.A(new_n1257), .B(new_n1258), .C1(new_n682), .C2(new_n687), .ZN(new_n1259));
  OAI21_X1  g833(.A(new_n1254), .B1(new_n1256), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g834(.A(new_n1260), .B1(new_n981), .B2(new_n982), .ZN(G308));
  OAI211_X1 g835(.A(new_n983), .B(new_n1254), .C1(new_n1256), .C2(new_n1259), .ZN(G225));
endmodule


