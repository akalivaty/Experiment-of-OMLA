//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n544, new_n545, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n561, new_n562, new_n563,
    new_n564, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n575, new_n576, new_n578, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n639, new_n640, new_n641, new_n644, new_n646, new_n647,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n852, new_n853, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1206, new_n1207, new_n1208;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT64), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT65), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT66), .Z(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n459));
  INV_X1    g034(.A(new_n453), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n459), .B1(G567), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n458), .A2(KEYINPUT67), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(new_n463), .ZN(G319));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G101), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n469));
  INV_X1    g044(.A(G2105), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT68), .ZN(new_n473));
  NAND3_X1  g048(.A1(new_n473), .A2(new_n465), .A3(KEYINPUT3), .ZN(new_n474));
  NAND4_X1  g049(.A1(new_n469), .A2(new_n470), .A3(new_n472), .A4(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n467), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND3_X1  g052(.A1(new_n468), .A2(new_n472), .A3(G125), .ZN(new_n478));
  NAND2_X1  g053(.A1(G113), .A2(G2104), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n470), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g056(.A(new_n481), .B(KEYINPUT69), .ZN(G160));
  AND2_X1   g057(.A1(new_n474), .A2(new_n472), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n483), .A2(G2105), .A3(new_n469), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G124), .ZN(new_n486));
  INV_X1    g061(.A(new_n475), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n487), .A2(KEYINPUT70), .A3(G136), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT70), .ZN(new_n489));
  INV_X1    g064(.A(G136), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n489), .B1(new_n475), .B2(new_n490), .ZN(new_n491));
  OR2_X1    g066(.A1(G100), .A2(G2105), .ZN(new_n492));
  OAI211_X1 g067(.A(new_n492), .B(G2104), .C1(G112), .C2(new_n470), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n486), .A2(new_n488), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G162));
  INV_X1    g070(.A(G114), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(G2105), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  XNOR2_X1  g073(.A(new_n497), .B(new_n498), .ZN(new_n499));
  OAI21_X1  g074(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G126), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n484), .B2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  OAI21_X1  g080(.A(KEYINPUT4), .B1(new_n475), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n468), .A2(new_n472), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n507), .A2(G2105), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n505), .A2(KEYINPUT4), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(KEYINPUT72), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  OAI211_X1 g086(.A(new_n511), .B(KEYINPUT4), .C1(new_n475), .C2(new_n505), .ZN(new_n512));
  AOI21_X1  g087(.A(new_n504), .B1(new_n510), .B2(new_n512), .ZN(G164));
  INV_X1    g088(.A(KEYINPUT73), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n514), .A2(G651), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n517));
  OAI21_X1  g092(.A(KEYINPUT6), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT6), .A2(G651), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  AND2_X1   g095(.A1(KEYINPUT5), .A2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(KEYINPUT5), .A2(G543), .ZN(new_n522));
  OAI21_X1  g097(.A(G88), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(G50), .A2(G543), .ZN(new_n524));
  AOI22_X1  g099(.A1(new_n518), .A2(new_n520), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT73), .B(G651), .ZN(new_n526));
  OAI21_X1  g101(.A(G62), .B1(new_n521), .B2(new_n522), .ZN(new_n527));
  NAND2_X1  g102(.A1(G75), .A2(G543), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n525), .A2(KEYINPUT74), .A3(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n532));
  OAI21_X1  g107(.A(new_n520), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n523), .A2(new_n524), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n527), .A2(new_n528), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n516), .A2(KEYINPUT73), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n514), .A2(G651), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n536), .A2(new_n539), .ZN(new_n540));
  AOI21_X1  g115(.A(new_n531), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n530), .A2(new_n541), .ZN(G303));
  INV_X1    g117(.A(G303), .ZN(G166));
  AOI21_X1  g118(.A(new_n532), .B1(new_n537), .B2(new_n538), .ZN(new_n544));
  OAI21_X1  g119(.A(G543), .B1(new_n544), .B2(new_n519), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G51), .ZN(new_n547));
  NOR2_X1   g122(.A1(new_n521), .A2(new_n522), .ZN(new_n548));
  AOI21_X1  g123(.A(new_n548), .B1(new_n518), .B2(new_n520), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G89), .ZN(new_n550));
  NAND3_X1  g125(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n551));
  OR2_X1    g126(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(KEYINPUT7), .ZN(new_n553));
  OR2_X1    g128(.A1(KEYINPUT5), .A2(G543), .ZN(new_n554));
  NAND2_X1  g129(.A1(KEYINPUT5), .A2(G543), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g131(.A1(G63), .A2(G651), .ZN(new_n557));
  AOI22_X1  g132(.A1(new_n552), .A2(new_n553), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n547), .A2(new_n550), .A3(new_n558), .ZN(G286));
  INV_X1    g134(.A(G286), .ZN(G168));
  NAND2_X1  g135(.A1(new_n546), .A2(G52), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n549), .A2(G90), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n556), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n526), .ZN(new_n564));
  AND3_X1   g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(G171));
  XOR2_X1   g140(.A(KEYINPUT75), .B(G43), .Z(new_n566));
  NAND2_X1  g141(.A1(new_n546), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n549), .A2(G81), .ZN(new_n568));
  AOI22_X1  g143(.A1(new_n556), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n569));
  OR2_X1    g144(.A1(new_n569), .A2(new_n526), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n567), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G860), .ZN(G153));
  NAND4_X1  g148(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g149(.A1(G1), .A2(G3), .ZN(new_n575));
  XNOR2_X1  g150(.A(new_n575), .B(KEYINPUT8), .ZN(new_n576));
  NAND4_X1  g151(.A1(G319), .A2(G483), .A3(G661), .A4(new_n576), .ZN(G188));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n546), .A2(new_n578), .A3(G53), .ZN(new_n579));
  INV_X1    g154(.A(G53), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT9), .B1(new_n545), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(G78), .A2(G543), .ZN(new_n583));
  INV_X1    g158(.A(G65), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n548), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n549), .A2(G91), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n582), .A2(new_n586), .A3(new_n587), .ZN(G299));
  INV_X1    g163(.A(G171), .ZN(G301));
  OAI211_X1 g164(.A(G49), .B(G543), .C1(new_n544), .C2(new_n519), .ZN(new_n590));
  OAI211_X1 g165(.A(G87), .B(new_n556), .C1(new_n544), .C2(new_n519), .ZN(new_n591));
  OAI21_X1  g166(.A(G651), .B1(new_n556), .B2(G74), .ZN(new_n592));
  NAND3_X1  g167(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(G288));
  OAI211_X1 g168(.A(G48), .B(G543), .C1(new_n544), .C2(new_n519), .ZN(new_n594));
  OAI211_X1 g169(.A(G86), .B(new_n556), .C1(new_n544), .C2(new_n519), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n596), .B1(new_n554), .B2(new_n555), .ZN(new_n597));
  AND2_X1   g172(.A1(G73), .A2(G543), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n539), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(G305));
  OAI211_X1 g175(.A(G47), .B(G543), .C1(new_n544), .C2(new_n519), .ZN(new_n601));
  OAI211_X1 g176(.A(G85), .B(new_n556), .C1(new_n544), .C2(new_n519), .ZN(new_n602));
  INV_X1    g177(.A(G60), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n554), .B2(new_n555), .ZN(new_n604));
  AND2_X1   g179(.A1(G72), .A2(G543), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n539), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(G290));
  INV_X1    g182(.A(KEYINPUT78), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT76), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n545), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n533), .A2(KEYINPUT76), .A3(G543), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n611), .A2(G54), .A3(new_n612), .ZN(new_n613));
  OAI211_X1 g188(.A(G92), .B(new_n556), .C1(new_n544), .C2(new_n519), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT10), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g191(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .A4(new_n556), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  AOI22_X1  g193(.A1(new_n556), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n619), .A2(new_n516), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(new_n621));
  AND4_X1   g196(.A1(new_n609), .A2(new_n613), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  INV_X1    g197(.A(G54), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n623), .B1(new_n545), .B2(new_n610), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n620), .B1(new_n624), .B2(new_n612), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n609), .B1(new_n625), .B2(new_n618), .ZN(new_n626));
  OAI21_X1  g201(.A(new_n608), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n613), .A2(new_n618), .A3(new_n621), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n628), .A2(KEYINPUT77), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n625), .A2(new_n609), .A3(new_n618), .ZN(new_n630));
  NAND3_X1  g205(.A1(new_n629), .A2(KEYINPUT78), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g206(.A1(new_n627), .A2(new_n631), .ZN(new_n632));
  INV_X1    g207(.A(G868), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(G171), .A2(G868), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT79), .ZN(G284));
  INV_X1    g212(.A(new_n636), .ZN(G321));
  NAND2_X1  g213(.A1(G286), .A2(G868), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n587), .A2(new_n586), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n581), .B2(new_n579), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n639), .B1(new_n641), .B2(G868), .ZN(G297));
  XNOR2_X1  g217(.A(G297), .B(KEYINPUT80), .ZN(G280));
  INV_X1    g218(.A(G559), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n632), .B1(new_n644), .B2(G860), .ZN(G148));
  NAND3_X1  g220(.A1(new_n627), .A2(new_n644), .A3(new_n631), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n646), .A2(G868), .ZN(new_n647));
  OAI21_X1  g222(.A(new_n647), .B1(G868), .B2(new_n572), .ZN(G323));
  XNOR2_X1  g223(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g224(.A1(new_n508), .A2(G2104), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT13), .ZN(new_n653));
  INV_X1    g228(.A(G2100), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  OAI21_X1  g230(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n656));
  INV_X1    g231(.A(G111), .ZN(new_n657));
  AOI22_X1  g232(.A1(new_n656), .A2(KEYINPUT82), .B1(new_n657), .B2(G2105), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(KEYINPUT82), .B2(new_n656), .ZN(new_n659));
  INV_X1    g234(.A(G135), .ZN(new_n660));
  INV_X1    g235(.A(G123), .ZN(new_n661));
  OAI221_X1 g236(.A(new_n659), .B1(new_n660), .B2(new_n475), .C1(new_n484), .C2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(G2096), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n655), .A2(new_n664), .ZN(G156));
  XNOR2_X1  g240(.A(KEYINPUT15), .B(G2435), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT84), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G2427), .B(G2430), .Z(new_n669));
  OR2_X1    g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n670), .A2(KEYINPUT14), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT85), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2451), .B(G2454), .ZN(new_n674));
  XNOR2_X1  g249(.A(G2443), .B(G2446), .ZN(new_n675));
  XOR2_X1   g250(.A(new_n674), .B(new_n675), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n673), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n678));
  XOR2_X1   g253(.A(new_n677), .B(new_n678), .Z(new_n679));
  XNOR2_X1  g254(.A(G1341), .B(G1348), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n679), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(KEYINPUT86), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT86), .ZN(new_n684));
  NAND3_X1  g259(.A1(new_n679), .A2(new_n684), .A3(new_n681), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g261(.A(G14), .ZN(new_n687));
  INV_X1    g262(.A(new_n679), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n680), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n686), .A2(new_n689), .ZN(G401));
  INV_X1    g265(.A(KEYINPUT18), .ZN(new_n691));
  XOR2_X1   g266(.A(G2084), .B(G2090), .Z(new_n692));
  XNOR2_X1  g267(.A(G2067), .B(G2678), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(KEYINPUT17), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n692), .A2(new_n693), .ZN(new_n696));
  OAI21_X1  g271(.A(new_n691), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(new_n654), .ZN(new_n698));
  XOR2_X1   g273(.A(G2072), .B(G2078), .Z(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n694), .B2(KEYINPUT18), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(new_n663), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(G227));
  XNOR2_X1  g277(.A(G1956), .B(G2474), .ZN(new_n703));
  XNOR2_X1  g278(.A(G1961), .B(G1966), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1971), .B(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n703), .A2(new_n704), .A3(KEYINPUT88), .ZN(new_n710));
  NAND3_X1  g285(.A1(new_n706), .A2(new_n709), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT20), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n703), .A2(new_n704), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n705), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(new_n714), .B(new_n713), .S(new_n709), .Z(new_n715));
  NAND2_X1  g290(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(G1991), .B(G1996), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1981), .B(G1986), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(new_n722), .ZN(G229));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n724), .A2(G23), .ZN(new_n725));
  INV_X1    g300(.A(G288), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n724), .ZN(new_n727));
  XOR2_X1   g302(.A(new_n727), .B(KEYINPUT90), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT33), .B(G1976), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n728), .A2(new_n729), .ZN(new_n731));
  NOR2_X1   g306(.A1(G6), .A2(G16), .ZN(new_n732));
  AND3_X1   g307(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n732), .B1(new_n733), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT32), .B(G1981), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(KEYINPUT89), .B(G16), .Z(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n738), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  NAND4_X1  g317(.A1(new_n730), .A2(new_n731), .A3(new_n736), .A4(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(KEYINPUT34), .ZN(new_n745));
  NOR2_X1   g320(.A1(G25), .A2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G119), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n470), .A2(G107), .ZN(new_n748));
  OAI21_X1  g323(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n749));
  OAI22_X1  g324(.A1(new_n484), .A2(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(G131), .B2(new_n487), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n746), .B1(new_n751), .B2(G29), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT35), .B(G1991), .Z(new_n753));
  XOR2_X1   g328(.A(new_n752), .B(new_n753), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n738), .A2(G24), .ZN(new_n755));
  AND3_X1   g330(.A1(new_n601), .A2(new_n602), .A3(new_n606), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n738), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(G1986), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n754), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n744), .A2(new_n745), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT36), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n724), .A2(G4), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(new_n632), .B2(new_n724), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(G1348), .Z(new_n764));
  NAND2_X1  g339(.A1(new_n724), .A2(G21), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(G168), .B2(new_n724), .ZN(new_n766));
  INV_X1    g341(.A(G1966), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n738), .A2(G19), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(new_n572), .B2(new_n738), .ZN(new_n770));
  INV_X1    g345(.A(G1341), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(G2084), .ZN(new_n773));
  NAND2_X1  g348(.A1(G160), .A2(G29), .ZN(new_n774));
  INV_X1    g349(.A(G29), .ZN(new_n775));
  INV_X1    g350(.A(KEYINPUT24), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n775), .B1(new_n776), .B2(G34), .ZN(new_n777));
  AND2_X1   g352(.A1(new_n777), .A2(KEYINPUT91), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n776), .A2(G34), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n779), .B1(new_n777), .B2(KEYINPUT91), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n774), .B1(new_n778), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n768), .B(new_n772), .C1(new_n773), .C2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n775), .A2(G26), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT28), .ZN(new_n784));
  INV_X1    g359(.A(G128), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n470), .A2(G116), .ZN(new_n786));
  OAI21_X1  g361(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n787));
  OAI22_X1  g362(.A1(new_n484), .A2(new_n785), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n487), .A2(G140), .ZN(new_n789));
  OR2_X1    g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n784), .B1(new_n791), .B2(new_n775), .ZN(new_n792));
  INV_X1    g367(.A(G2067), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n792), .B(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n775), .A2(G33), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n470), .A2(G103), .A3(G2104), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT25), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n468), .A2(new_n472), .A3(G127), .ZN(new_n798));
  NAND2_X1  g373(.A1(G115), .A2(G2104), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n470), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI211_X1 g375(.A(new_n797), .B(new_n800), .C1(G139), .C2(new_n487), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(new_n775), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(G2072), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT31), .B(G11), .ZN(new_n804));
  INV_X1    g379(.A(G28), .ZN(new_n805));
  AOI21_X1  g380(.A(G29), .B1(new_n805), .B2(KEYINPUT30), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n807), .A2(KEYINPUT94), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n807), .A2(KEYINPUT94), .B1(KEYINPUT30), .B2(new_n805), .ZN(new_n809));
  OAI221_X1 g384(.A(new_n804), .B1(new_n808), .B2(new_n809), .C1(new_n662), .C2(new_n775), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G2072), .B2(new_n802), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n724), .A2(G5), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(G171), .B2(new_n724), .ZN(new_n813));
  INV_X1    g388(.A(G1961), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n794), .A2(new_n803), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(G2090), .ZN(new_n817));
  NOR2_X1   g392(.A1(G29), .A2(G35), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G162), .B2(G29), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  AOI211_X1 g396(.A(new_n782), .B(new_n816), .C1(new_n817), .C2(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n738), .A2(G20), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(KEYINPUT23), .Z(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G299), .B2(G16), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1956), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(new_n821), .B2(new_n817), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(KEYINPUT96), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n775), .A2(G32), .ZN(new_n829));
  NAND3_X1  g404(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT26), .ZN(new_n831));
  OR2_X1    g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  AOI22_X1  g408(.A1(new_n832), .A2(new_n833), .B1(G105), .B2(new_n466), .ZN(new_n834));
  INV_X1    g409(.A(G129), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n484), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G141), .B2(new_n487), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT92), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n829), .B1(new_n839), .B2(new_n775), .ZN(new_n840));
  XNOR2_X1  g415(.A(KEYINPUT27), .B(G1996), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT93), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g418(.A1(new_n840), .A2(new_n842), .B1(new_n773), .B2(new_n781), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n775), .A2(G27), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(G164), .B2(new_n775), .ZN(new_n846));
  INV_X1    g421(.A(G2078), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  AND3_X1   g423(.A1(new_n843), .A2(new_n844), .A3(new_n848), .ZN(new_n849));
  AND4_X1   g424(.A1(new_n764), .A2(new_n822), .A3(new_n828), .A4(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n761), .A2(new_n850), .ZN(G311));
  AND3_X1   g426(.A1(new_n761), .A2(KEYINPUT97), .A3(new_n850), .ZN(new_n852));
  AOI21_X1  g427(.A(KEYINPUT97), .B1(new_n761), .B2(new_n850), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n853), .ZN(G150));
  NAND2_X1  g429(.A1(new_n632), .A2(G559), .ZN(new_n855));
  XOR2_X1   g430(.A(KEYINPUT98), .B(KEYINPUT38), .Z(new_n856));
  XNOR2_X1  g431(.A(new_n855), .B(new_n856), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n556), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n858), .A2(new_n526), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n859), .B(KEYINPUT99), .Z(new_n860));
  AOI22_X1  g435(.A1(new_n546), .A2(G55), .B1(new_n549), .B2(G93), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n571), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n859), .B(KEYINPUT99), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n572), .A2(new_n864), .A3(new_n861), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n857), .B(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT39), .ZN(new_n869));
  AOI21_X1  g444(.A(G860), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n870), .B1(new_n869), .B2(new_n868), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n860), .A2(new_n862), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(G860), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT37), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n871), .A2(new_n875), .ZN(G145));
  XOR2_X1   g451(.A(KEYINPUT100), .B(G37), .Z(new_n877));
  XNOR2_X1  g452(.A(G164), .B(new_n790), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n487), .A2(G142), .ZN(new_n879));
  INV_X1    g454(.A(G130), .ZN(new_n880));
  NOR2_X1   g455(.A1(new_n470), .A2(G118), .ZN(new_n881));
  OAI21_X1  g456(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n882));
  OAI221_X1 g457(.A(new_n879), .B1(new_n880), .B2(new_n484), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n878), .B(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n751), .B(new_n652), .ZN(new_n885));
  OR2_X1    g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n884), .A2(new_n885), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n837), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(new_n801), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n838), .B2(new_n801), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(G160), .B(G162), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(new_n662), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n891), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n886), .A2(new_n887), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n892), .A2(new_n895), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g474(.A(new_n895), .B1(new_n892), .B2(new_n897), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n877), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n646), .A2(new_n867), .ZN(new_n905));
  NAND4_X1  g480(.A1(new_n866), .A2(new_n644), .A3(new_n627), .A4(new_n631), .ZN(new_n906));
  INV_X1    g481(.A(new_n628), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n907), .A2(new_n641), .ZN(new_n908));
  NOR2_X1   g483(.A1(G299), .A2(new_n628), .ZN(new_n909));
  NOR2_X1   g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND3_X1   g485(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(KEYINPUT41), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n912), .B1(new_n908), .B2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n907), .A2(new_n641), .ZN(new_n914));
  NAND2_X1  g489(.A1(G299), .A2(new_n628), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT41), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n917), .B1(new_n905), .B2(new_n906), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n904), .B1(new_n911), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n905), .A2(new_n906), .ZN(new_n920));
  INV_X1    g495(.A(new_n917), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n905), .A2(new_n906), .A3(new_n910), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(KEYINPUT104), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT103), .ZN(new_n925));
  OAI21_X1  g500(.A(KEYINPUT74), .B1(new_n525), .B2(new_n529), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n535), .A2(new_n540), .A3(new_n531), .ZN(new_n927));
  AND3_X1   g502(.A1(new_n926), .A2(new_n927), .A3(G305), .ZN(new_n928));
  AOI21_X1  g503(.A(G305), .B1(new_n926), .B2(new_n927), .ZN(new_n929));
  AND2_X1   g504(.A1(G288), .A2(G290), .ZN(new_n930));
  NOR2_X1   g505(.A1(G288), .A2(G290), .ZN(new_n931));
  OAI22_X1  g506(.A1(new_n928), .A2(new_n929), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n733), .B1(new_n530), .B2(new_n541), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n726), .A2(new_n756), .ZN(new_n934));
  NAND2_X1  g509(.A1(G288), .A2(G290), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n926), .A2(new_n927), .A3(G305), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n933), .A2(new_n934), .A3(new_n935), .A4(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(KEYINPUT101), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n932), .A2(new_n937), .A3(KEYINPUT101), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n932), .A2(new_n937), .A3(KEYINPUT102), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n942), .A2(KEYINPUT42), .ZN(new_n943));
  INV_X1    g518(.A(new_n937), .ZN(new_n944));
  AOI22_X1  g519(.A1(new_n933), .A2(new_n936), .B1(new_n934), .B2(new_n935), .ZN(new_n945));
  NOR4_X1   g520(.A1(new_n944), .A2(new_n945), .A3(KEYINPUT102), .A4(KEYINPUT42), .ZN(new_n946));
  INV_X1    g521(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n925), .B1(new_n943), .B2(new_n947), .ZN(new_n948));
  AOI211_X1 g523(.A(KEYINPUT103), .B(new_n946), .C1(new_n942), .C2(KEYINPUT42), .ZN(new_n949));
  OAI211_X1 g524(.A(new_n919), .B(new_n924), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n922), .A2(new_n923), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT42), .ZN(new_n953));
  AND3_X1   g528(.A1(new_n932), .A2(KEYINPUT101), .A3(new_n937), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n954), .A2(new_n938), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n955), .B2(new_n941), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT103), .B1(new_n956), .B2(new_n946), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n943), .A2(new_n925), .A3(new_n947), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n952), .A2(new_n957), .A3(new_n904), .A4(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G868), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n903), .B1(new_n951), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n873), .A2(new_n633), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n950), .A2(KEYINPUT105), .A3(G868), .A4(new_n959), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n961), .A2(new_n962), .A3(new_n963), .ZN(G295));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n962), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n948), .A2(new_n949), .ZN(new_n966));
  INV_X1    g541(.A(new_n919), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n633), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(KEYINPUT105), .B1(new_n968), .B2(new_n950), .ZN(new_n969));
  OAI21_X1  g544(.A(KEYINPUT106), .B1(new_n965), .B2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n961), .A2(new_n971), .A3(new_n962), .A4(new_n963), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n970), .A2(new_n972), .ZN(G331));
  INV_X1    g548(.A(KEYINPUT107), .ZN(new_n974));
  OAI21_X1  g549(.A(G286), .B1(G171), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G171), .A2(new_n974), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n975), .B(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n866), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n910), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n977), .A2(new_n867), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(KEYINPUT108), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n977), .A2(new_n983), .A3(new_n867), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n980), .B1(new_n982), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n917), .B1(new_n979), .B2(new_n981), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n955), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n979), .A2(new_n910), .A3(new_n981), .ZN(new_n988));
  AOI22_X1  g563(.A1(new_n982), .A2(new_n984), .B1(new_n866), .B2(new_n978), .ZN(new_n989));
  OAI221_X1 g564(.A(new_n988), .B1(new_n954), .B2(new_n938), .C1(new_n989), .C2(new_n917), .ZN(new_n990));
  AND4_X1   g565(.A1(KEYINPUT43), .A2(new_n987), .A3(new_n990), .A4(new_n877), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n988), .B1(new_n989), .B2(new_n917), .ZN(new_n992));
  AOI21_X1  g567(.A(G37), .B1(new_n992), .B2(new_n955), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT43), .B1(new_n993), .B2(new_n990), .ZN(new_n994));
  OAI21_X1  g569(.A(KEYINPUT44), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT43), .ZN(new_n996));
  AND4_X1   g571(.A1(new_n996), .A2(new_n987), .A3(new_n990), .A4(new_n877), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n996), .B1(new_n993), .B2(new_n990), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n995), .B1(new_n999), .B2(KEYINPUT44), .ZN(G397));
  NOR2_X1   g575(.A1(G164), .A2(G1384), .ZN(new_n1001));
  AND2_X1   g576(.A1(new_n1001), .A2(KEYINPUT109), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1003), .B1(new_n1001), .B2(KEYINPUT109), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n481), .A2(G40), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g581(.A(new_n790), .B(G2067), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(G1996), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(new_n1009), .B2(new_n837), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n1009), .B2(new_n839), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n751), .B(new_n753), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT112), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g589(.A1(G290), .A2(G1986), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT110), .Z(new_n1016));
  NAND2_X1  g591(.A1(G290), .A2(G1986), .ZN(new_n1017));
  XOR2_X1   g592(.A(new_n1017), .B(KEYINPUT111), .Z(new_n1018));
  OR2_X1    g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1006), .B1(new_n1014), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G8), .ZN(new_n1021));
  NOR2_X1   g596(.A1(G166), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n1022), .A2(KEYINPUT55), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(KEYINPUT55), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n510), .A2(new_n512), .ZN(new_n1026));
  INV_X1    g601(.A(new_n504), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G1384), .ZN(new_n1029));
  AOI21_X1  g604(.A(KEYINPUT45), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1005), .ZN(new_n1031));
  NOR2_X1   g606(.A1(new_n1003), .A2(G1384), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1031), .B1(G164), .B2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n741), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(KEYINPUT50), .A2(G1384), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1005), .B1(new_n1028), .B2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1038));
  XNOR2_X1  g613(.A(KEYINPUT113), .B(G2090), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1037), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1021), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1043), .B2(new_n1042), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1021), .B1(new_n1001), .B2(new_n1031), .ZN(new_n1046));
  INV_X1    g621(.A(G1976), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1046), .B1(new_n1047), .B2(G288), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(KEYINPUT52), .ZN(new_n1049));
  NAND2_X1  g624(.A1(G305), .A2(G1981), .ZN(new_n1050));
  OR2_X1    g625(.A1(G305), .A2(G1981), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(KEYINPUT114), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1051), .B(KEYINPUT114), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1057), .A2(KEYINPUT49), .A3(new_n1050), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1056), .A2(new_n1046), .A3(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(KEYINPUT52), .B1(G288), .B2(new_n1047), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1046), .B(new_n1060), .C1(new_n1047), .C2(G288), .ZN(new_n1061));
  AND3_X1   g636(.A1(new_n1049), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1041), .A2(new_n1025), .ZN(new_n1063));
  AND2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n767), .B1(new_n1030), .B2(new_n1034), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1037), .A2(new_n773), .A3(new_n1038), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT116), .ZN(new_n1068));
  NOR2_X1   g643(.A1(G286), .A2(new_n1021), .ZN(new_n1069));
  AND3_X1   g644(.A1(new_n1067), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1068), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1045), .A2(new_n1064), .A3(new_n1073), .A4(KEYINPUT63), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT63), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT115), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1025), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1042), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(KEYINPUT115), .B1(new_n1041), .B2(new_n1025), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1078), .A2(new_n1062), .A3(new_n1079), .A4(new_n1063), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1075), .B1(new_n1080), .B2(new_n1072), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1074), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1005), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n1003), .B1(G164), .B2(G1384), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n847), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT53), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n814), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1083), .A2(KEYINPUT53), .A3(new_n847), .A4(new_n1084), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1080), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(G8), .B1(new_n1067), .B2(G286), .ZN(new_n1094));
  AOI21_X1  g669(.A(G168), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1095));
  OAI21_X1  g670(.A(KEYINPUT51), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT51), .ZN(new_n1097));
  OAI211_X1 g672(.A(new_n1097), .B(G8), .C1(new_n1067), .C2(G286), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT62), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT62), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1096), .A2(new_n1098), .A3(new_n1101), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1093), .A2(new_n1100), .A3(new_n1102), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1059), .A2(new_n1047), .A3(new_n726), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1057), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1063), .ZN(new_n1106));
  AOI22_X1  g681(.A1(new_n1105), .A2(new_n1046), .B1(new_n1062), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1082), .A2(new_n1103), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT122), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n477), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n477), .A2(new_n1109), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT123), .B(G2078), .Z(new_n1112));
  NAND2_X1  g687(.A1(KEYINPUT53), .A2(G40), .ZN(new_n1113));
  NOR3_X1   g688(.A1(new_n480), .A2(new_n1112), .A3(new_n1113), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1110), .A2(new_n1111), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1115), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1116), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1117), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1092), .B1(G171), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n1120));
  AOI22_X1  g695(.A1(new_n1119), .A2(new_n1120), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1080), .ZN(new_n1122));
  OAI21_X1  g697(.A(KEYINPUT124), .B1(new_n1091), .B2(G171), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1118), .A2(G171), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1118), .A2(KEYINPUT124), .A3(G171), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(KEYINPUT54), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(G1956), .ZN(new_n1128));
  AOI21_X1  g703(.A(KEYINPUT118), .B1(new_n1088), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT118), .ZN(new_n1130));
  AOI211_X1 g705(.A(new_n1130), .B(G1956), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1131));
  OR2_X1    g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n641), .B(KEYINPUT57), .ZN(new_n1133));
  XNOR2_X1  g708(.A(KEYINPUT56), .B(G2072), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1083), .A2(new_n1084), .A3(new_n1134), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1132), .A2(KEYINPUT119), .A3(new_n1133), .A4(new_n1135), .ZN(new_n1136));
  OAI211_X1 g711(.A(new_n1133), .B(new_n1135), .C1(new_n1129), .C2(new_n1131), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT119), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g714(.A(KEYINPUT61), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1121), .A2(new_n1122), .A3(new_n1127), .A4(new_n1141), .ZN(new_n1142));
  AOI21_X1  g717(.A(G1348), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1001), .A2(new_n1031), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n1144), .A2(G2067), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n622), .A2(new_n626), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1146), .A2(new_n1149), .A3(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(KEYINPUT60), .B(new_n1148), .C1(new_n1143), .C2(new_n1145), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1083), .A2(new_n1009), .A3(new_n1084), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1083), .A2(KEYINPUT120), .A3(new_n1009), .A4(new_n1084), .ZN(new_n1157));
  XNOR2_X1  g732(.A(KEYINPUT121), .B(KEYINPUT58), .ZN(new_n1158));
  XNOR2_X1  g733(.A(new_n1158), .B(new_n771), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1144), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n1161), .A2(new_n572), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT59), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT59), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1164), .A3(new_n572), .ZN(new_n1165));
  AOI21_X1  g740(.A(new_n1153), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1135), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1133), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1169), .A2(KEYINPUT61), .A3(new_n1137), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1169), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1166), .A2(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  NOR2_X1   g748(.A1(new_n1142), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1020), .B1(new_n1108), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(KEYINPUT127), .ZN(new_n1176));
  AND2_X1   g751(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT126), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1177), .A2(new_n1178), .A3(KEYINPUT46), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1180));
  INV_X1    g755(.A(KEYINPUT46), .ZN(new_n1181));
  OAI21_X1  g756(.A(KEYINPUT126), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1179), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1008), .A2(new_n837), .ZN(new_n1184));
  AOI22_X1  g759(.A1(new_n1180), .A2(new_n1181), .B1(new_n1006), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1176), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1186), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1178), .B1(new_n1177), .B2(KEYINPUT46), .ZN(new_n1188));
  NOR3_X1   g763(.A1(new_n1180), .A2(KEYINPUT126), .A3(new_n1181), .ZN(new_n1189));
  OAI211_X1 g764(.A(new_n1176), .B(new_n1185), .C1(new_n1188), .C2(new_n1189), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1187), .A2(KEYINPUT47), .A3(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(KEYINPUT47), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1190), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1192), .B1(new_n1193), .B2(new_n1186), .ZN(new_n1194));
  AOI21_X1  g769(.A(KEYINPUT48), .B1(new_n1006), .B2(new_n1016), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1195), .B1(new_n1014), .B2(new_n1006), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1006), .A2(KEYINPUT48), .A3(new_n1016), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n751), .A2(new_n753), .ZN(new_n1198));
  XNOR2_X1  g773(.A(new_n1198), .B(KEYINPUT125), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1011), .A2(new_n1199), .ZN(new_n1200));
  OAI21_X1  g775(.A(new_n1200), .B1(G2067), .B2(new_n790), .ZN(new_n1201));
  AOI22_X1  g776(.A1(new_n1196), .A2(new_n1197), .B1(new_n1201), .B2(new_n1006), .ZN(new_n1202));
  AND3_X1   g777(.A1(new_n1191), .A2(new_n1194), .A3(new_n1202), .ZN(new_n1203));
  NAND2_X1  g778(.A1(new_n1175), .A2(new_n1203), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g779(.A1(new_n463), .A2(G227), .ZN(new_n1206));
  NAND2_X1  g780(.A1(new_n722), .A2(new_n1206), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n1207), .B1(new_n686), .B2(new_n689), .ZN(new_n1208));
  OAI211_X1 g782(.A(new_n1208), .B(new_n901), .C1(new_n998), .C2(new_n997), .ZN(G225));
  INV_X1    g783(.A(G225), .ZN(G308));
endmodule


