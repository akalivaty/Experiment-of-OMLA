//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G237), .ZN(new_n189));
  INV_X1    g003(.A(G953), .ZN(new_n190));
  AND4_X1   g004(.A1(G143), .A2(new_n189), .A3(new_n190), .A4(G214), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  AOI21_X1  g006(.A(G143), .B1(new_n192), .B2(G214), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT18), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G140), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G125), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G140), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n197), .A2(new_n199), .A3(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n194), .A2(new_n195), .B1(new_n201), .B2(new_n203), .ZN(new_n204));
  OAI211_X1 g018(.A(KEYINPUT18), .B(G131), .C1(new_n191), .C2(new_n193), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  OAI21_X1  g020(.A(G131), .B1(new_n191), .B2(new_n193), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(KEYINPUT17), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n194), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(new_n207), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n209), .B1(new_n212), .B2(KEYINPUT17), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT16), .ZN(new_n214));
  OR3_X1    g028(.A1(new_n198), .A2(KEYINPUT16), .A3(G140), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G146), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT71), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n214), .A2(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n202), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n216), .A2(new_n221), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n218), .A2(new_n220), .A3(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n206), .B1(new_n213), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g038(.A(G113), .B(G122), .ZN(new_n225));
  INV_X1    g039(.A(G104), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n225), .B(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  OAI211_X1 g043(.A(new_n227), .B(new_n206), .C1(new_n213), .C2(new_n223), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n188), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G475), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT82), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT19), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n200), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n197), .A2(new_n199), .A3(KEYINPUT19), .ZN(new_n237));
  AOI21_X1  g051(.A(G146), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n238), .A2(new_n217), .ZN(new_n239));
  AOI22_X1  g053(.A1(new_n239), .A2(new_n212), .B1(new_n205), .B2(new_n204), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n234), .B1(new_n240), .B2(new_n227), .ZN(new_n241));
  INV_X1    g055(.A(new_n237), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT19), .B1(new_n197), .B2(new_n199), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n202), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n191), .A2(new_n193), .A3(G131), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n244), .B(new_n216), .C1(new_n208), .C2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(new_n206), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT82), .A3(new_n228), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n241), .A2(new_n230), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT83), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n251), .A2(new_n252), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  AND4_X1   g068(.A1(KEYINPUT83), .A2(new_n249), .A3(new_n252), .A4(new_n253), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n233), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G478), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(KEYINPUT15), .ZN(new_n258));
  INV_X1    g072(.A(G116), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G122), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT85), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(new_n261), .A3(KEYINPUT14), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n261), .B1(new_n260), .B2(KEYINPUT14), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G122), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G116), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n267), .B1(new_n260), .B2(KEYINPUT14), .ZN(new_n268));
  OAI21_X1  g082(.A(G107), .B1(new_n265), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G107), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n260), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G128), .ZN(new_n274));
  INV_X1    g088(.A(G128), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(G143), .ZN(new_n276));
  INV_X1    g090(.A(G134), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n276), .A3(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n274), .A2(new_n276), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G134), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n272), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n267), .A2(new_n260), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G107), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n271), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT13), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n285), .B1(new_n275), .B2(G143), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n276), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n274), .A2(new_n285), .ZN(new_n288));
  OAI21_X1  g102(.A(G134), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n284), .A2(new_n289), .A3(new_n278), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT84), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n269), .A2(new_n281), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n284), .A2(new_n289), .A3(KEYINPUT84), .A4(new_n278), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  INV_X1    g108(.A(G217), .ZN(new_n295));
  NOR3_X1   g109(.A1(new_n294), .A2(new_n295), .A3(G953), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n292), .A2(new_n293), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n290), .A2(new_n291), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n260), .A2(KEYINPUT14), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT85), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n268), .B1(new_n300), .B2(new_n262), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n281), .B1(new_n270), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(new_n302), .A3(new_n293), .ZN(new_n303));
  INV_X1    g117(.A(new_n296), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n297), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n188), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n258), .B1(new_n307), .B2(KEYINPUT86), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT86), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n306), .B2(new_n188), .ZN(new_n310));
  AOI211_X1 g124(.A(KEYINPUT86), .B(G902), .C1(new_n297), .C2(new_n305), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n308), .B1(new_n312), .B2(new_n258), .ZN(new_n313));
  INV_X1    g127(.A(G952), .ZN(new_n314));
  NOR2_X1   g128(.A1(new_n314), .A2(G953), .ZN(new_n315));
  INV_X1    g129(.A(G234), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n315), .B1(new_n316), .B2(new_n189), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI211_X1 g132(.A(new_n188), .B(new_n190), .C1(G234), .C2(G237), .ZN(new_n319));
  XNOR2_X1  g133(.A(KEYINPUT21), .B(G898), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NOR3_X1   g135(.A1(new_n256), .A2(new_n313), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(G221), .B1(new_n294), .B2(G902), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G469), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n325), .A2(new_n188), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT1), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n202), .A2(G143), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n273), .A2(G146), .ZN(new_n329));
  AND4_X1   g143(.A1(new_n327), .A2(new_n328), .A3(new_n329), .A4(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n331));
  XNOR2_X1  g145(.A(G143), .B(G146), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n327), .A3(G128), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT75), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n273), .A2(KEYINPUT1), .A3(G146), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n332), .B2(G128), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n331), .A2(new_n335), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n270), .A2(G104), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n226), .A2(G107), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g156(.A1(new_n342), .A2(G101), .ZN(new_n343));
  OAI21_X1  g157(.A(KEYINPUT3), .B1(new_n226), .B2(G107), .ZN(new_n344));
  AOI21_X1  g158(.A(G101), .B1(new_n226), .B2(G107), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT3), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(new_n270), .A3(G104), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT74), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT74), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n344), .A2(new_n345), .A3(new_n347), .A4(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n343), .B1(new_n349), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n339), .A2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT10), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n349), .A2(new_n351), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT4), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n347), .A3(new_n341), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n358), .B2(G101), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n328), .A2(new_n329), .ZN(new_n361));
  NAND2_X1  g175(.A1(KEYINPUT0), .A2(G128), .ZN(new_n362));
  OR2_X1    g176(.A1(KEYINPUT0), .A2(G128), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n361), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n332), .A2(KEYINPUT0), .A3(G128), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n358), .A2(new_n357), .A3(G101), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n360), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT11), .B1(new_n277), .B2(G137), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT11), .ZN(new_n370));
  INV_X1    g184(.A(G137), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(G134), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT64), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n374), .B1(new_n371), .B2(G134), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n277), .A2(KEYINPUT64), .A3(G137), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n373), .A2(new_n210), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n210), .B1(new_n379), .B2(new_n373), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT65), .ZN(new_n382));
  AOI21_X1  g196(.A(G128), .B1(new_n328), .B2(new_n329), .ZN(new_n383));
  INV_X1    g197(.A(new_n336), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n336), .B(KEYINPUT65), .C1(new_n332), .C2(G128), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(new_n333), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n352), .A2(new_n387), .A3(KEYINPUT10), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n355), .A2(new_n368), .A3(new_n381), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n353), .B1(new_n387), .B2(new_n352), .ZN(new_n390));
  INV_X1    g204(.A(new_n381), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT12), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT76), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n392), .B1(new_n381), .B2(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n390), .A2(new_n391), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n390), .B2(new_n391), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n389), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(G110), .B(G140), .ZN(new_n398));
  INV_X1    g212(.A(G227), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(G953), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n398), .B(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n389), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n355), .A2(new_n368), .A3(new_n388), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(new_n391), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n397), .A2(new_n401), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n326), .B1(new_n407), .B2(G469), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n395), .A2(new_n396), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n409), .A2(new_n403), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n402), .B1(new_n406), .B2(new_n389), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n325), .B(new_n188), .C1(new_n410), .C2(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n324), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G210), .B1(G237), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n343), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n356), .A2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT2), .B(G113), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  OR2_X1    g233(.A1(KEYINPUT66), .A2(G119), .ZN(new_n420));
  NAND2_X1  g234(.A1(KEYINPUT66), .A2(G119), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n420), .A2(G116), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n259), .A2(G119), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND3_X1   g238(.A1(new_n422), .A2(KEYINPUT5), .A3(new_n423), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT5), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n420), .A2(new_n426), .A3(G116), .A4(new_n421), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(G113), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n424), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n417), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n422), .A2(new_n423), .ZN(new_n431));
  OAI211_X1 g245(.A(G113), .B(new_n427), .C1(new_n431), .C2(new_n426), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n352), .A2(new_n424), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  XNOR2_X1  g248(.A(G110), .B(G122), .ZN(new_n435));
  XOR2_X1   g249(.A(new_n435), .B(KEYINPUT8), .Z(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT79), .B1(new_n434), .B2(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT79), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n439), .B(new_n436), .C1(new_n430), .C2(new_n433), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n190), .A2(G224), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT80), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n443), .A2(KEYINPUT80), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n330), .B1(new_n337), .B2(new_n382), .ZN(new_n448));
  AOI21_X1  g262(.A(G125), .B1(new_n448), .B2(new_n386), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n364), .A2(new_n365), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n450), .A2(new_n198), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n446), .B(new_n447), .C1(new_n449), .C2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n451), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n387), .A2(new_n198), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n445), .A4(new_n444), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT77), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n457), .B1(new_n417), .B2(new_n429), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n431), .A2(new_n418), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n424), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n360), .A2(new_n460), .A3(new_n367), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n352), .A2(new_n432), .A3(KEYINPUT77), .A4(new_n424), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n461), .A3(new_n435), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n456), .A2(new_n463), .ZN(new_n464));
  OAI211_X1 g278(.A(KEYINPUT81), .B(new_n188), .C1(new_n441), .C2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n453), .A2(new_n454), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n466), .B(new_n442), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n458), .A2(new_n462), .A3(new_n461), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n435), .A2(KEYINPUT78), .ZN(new_n469));
  AOI22_X1  g283(.A1(KEYINPUT6), .A2(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n468), .A2(KEYINPUT6), .A3(new_n469), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n467), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n463), .B(new_n456), .C1(new_n438), .C2(new_n440), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT81), .B1(new_n474), .B2(new_n188), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n415), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n188), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g293(.A1(new_n479), .A2(new_n414), .A3(new_n472), .A4(new_n465), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  AND4_X1   g295(.A1(new_n187), .A2(new_n322), .A3(new_n413), .A4(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n371), .A2(G134), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n277), .A2(G137), .ZN(new_n484));
  OAI21_X1  g298(.A(G131), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n377), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n387), .ZN(new_n487));
  INV_X1    g301(.A(new_n460), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n366), .B1(new_n378), .B2(new_n380), .ZN(new_n489));
  AND3_X1   g303(.A1(new_n487), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n377), .A2(new_n485), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n448), .B2(new_n386), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G131), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n450), .B1(new_n494), .B2(new_n377), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT30), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT30), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n487), .A2(new_n489), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n490), .B1(new_n499), .B2(new_n460), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT67), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT31), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n192), .A2(G210), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT27), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT26), .B(G101), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n500), .A2(new_n501), .A3(new_n502), .A4(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT30), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n497), .B1(new_n487), .B2(new_n489), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n460), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n487), .A2(new_n489), .A3(new_n488), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n510), .A2(new_n502), .A3(new_n511), .A4(new_n506), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT67), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n488), .B1(new_n487), .B2(new_n489), .ZN(new_n514));
  OAI21_X1  g328(.A(KEYINPUT28), .B1(new_n490), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n515), .A2(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n506), .ZN(new_n519));
  AOI21_X1  g333(.A(KEYINPUT31), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n488), .B1(new_n496), .B2(new_n498), .ZN(new_n521));
  NOR3_X1   g335(.A1(new_n521), .A2(new_n490), .A3(new_n519), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n507), .B(new_n513), .C1(new_n520), .C2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G472), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n523), .A2(new_n524), .A3(new_n188), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT32), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT32), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n523), .A2(new_n527), .A3(new_n524), .A4(new_n188), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n515), .A2(new_n506), .A3(new_n517), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT29), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n188), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND4_X1  g346(.A1(new_n515), .A2(KEYINPUT68), .A3(new_n506), .A4(new_n517), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n519), .B1(new_n521), .B2(new_n490), .ZN(new_n534));
  AND3_X1   g348(.A1(new_n533), .A2(new_n534), .A3(new_n531), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT68), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n530), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n532), .B1(new_n535), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g352(.A(KEYINPUT69), .B1(new_n538), .B2(new_n524), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT69), .ZN(new_n540));
  INV_X1    g354(.A(new_n537), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n533), .A2(new_n534), .A3(new_n531), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g357(.A(new_n540), .B(G472), .C1(new_n543), .C2(new_n532), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n539), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n529), .A2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT25), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n420), .A2(new_n421), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G128), .ZN(new_n549));
  OR2_X1    g363(.A1(G119), .A2(G128), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT24), .B(G110), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(KEYINPUT23), .A3(new_n550), .ZN(new_n553));
  AOI21_X1  g367(.A(G128), .B1(new_n420), .B2(new_n421), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(KEYINPUT23), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n552), .B1(new_n555), .B2(G110), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n556), .A2(new_n216), .A3(new_n203), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n551), .B1(new_n549), .B2(new_n550), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT70), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n555), .A2(G110), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n223), .A3(new_n560), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT22), .B(G137), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n190), .A2(G221), .A3(G234), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n562), .B(new_n563), .Z(new_n564));
  AND3_X1   g378(.A1(new_n557), .A2(new_n561), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n557), .B2(new_n561), .ZN(new_n566));
  NOR3_X1   g380(.A1(new_n565), .A2(new_n566), .A3(G902), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n547), .B1(new_n567), .B2(KEYINPUT72), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n295), .B1(G234), .B2(new_n188), .ZN(new_n569));
  INV_X1    g383(.A(new_n566), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n557), .A2(new_n561), .A3(new_n564), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n188), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT72), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT25), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n568), .A2(new_n569), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n565), .A2(new_n566), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n569), .A2(G902), .ZN(new_n577));
  XOR2_X1   g391(.A(new_n577), .B(KEYINPUT73), .Z(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n575), .A2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n482), .A2(new_n546), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(new_n582), .B(G101), .ZN(G3));
  INV_X1    g397(.A(KEYINPUT88), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT87), .ZN(new_n585));
  AND3_X1   g399(.A1(new_n476), .A2(new_n585), .A3(new_n480), .ZN(new_n586));
  OAI211_X1 g400(.A(KEYINPUT87), .B(new_n415), .C1(new_n473), .C2(new_n475), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n187), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n584), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n476), .A2(new_n480), .A3(new_n585), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n590), .A2(KEYINPUT88), .A3(new_n187), .A4(new_n587), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(KEYINPUT90), .B(G478), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n307), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n296), .B1(new_n292), .B2(new_n293), .ZN(new_n595));
  AND4_X1   g409(.A1(new_n293), .A2(new_n298), .A3(new_n302), .A4(new_n296), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT33), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT33), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n297), .A2(new_n305), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n257), .A2(G902), .ZN(new_n601));
  AOI21_X1  g415(.A(KEYINPUT89), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT89), .ZN(new_n603));
  INV_X1    g417(.A(new_n601), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n603), .B(new_n604), .C1(new_n597), .C2(new_n599), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n594), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n256), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n321), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n524), .B1(new_n523), .B2(new_n188), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n525), .ZN(new_n611));
  INV_X1    g425(.A(new_n413), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n611), .A2(new_n612), .A3(new_n580), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n592), .A2(new_n608), .A3(new_n613), .ZN(new_n614));
  XOR2_X1   g428(.A(KEYINPUT34), .B(G104), .Z(new_n615));
  XNOR2_X1  g429(.A(new_n614), .B(new_n615), .ZN(G6));
  NOR2_X1   g430(.A1(KEYINPUT91), .A2(KEYINPUT20), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n617), .B1(new_n249), .B2(new_n253), .ZN(new_n618));
  NAND2_X1  g432(.A1(KEYINPUT91), .A2(KEYINPUT20), .ZN(new_n619));
  XOR2_X1   g433(.A(new_n619), .B(KEYINPUT92), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n618), .B(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n321), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n313), .A3(new_n233), .A4(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT93), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n623), .B(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n592), .A2(new_n613), .A3(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT35), .B(G107), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  NAND2_X1  g442(.A1(new_n557), .A2(new_n561), .ZN(new_n629));
  INV_X1    g443(.A(new_n564), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n630), .A2(KEYINPUT36), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n632), .A2(new_n578), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n575), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n610), .A2(new_n634), .A3(new_n525), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT94), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n610), .A2(new_n634), .A3(KEYINPUT94), .A4(new_n525), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n482), .A3(new_n638), .ZN(new_n639));
  XNOR2_X1  g453(.A(KEYINPUT37), .B(G110), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(KEYINPUT95), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n639), .B(new_n641), .ZN(G12));
  INV_X1    g456(.A(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n318), .B1(new_n319), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n621), .A2(new_n313), .A3(new_n233), .A4(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n546), .A2(new_n634), .A3(new_n647), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n589), .A2(new_n413), .A3(new_n591), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n650), .B(new_n275), .ZN(G30));
  INV_X1    g465(.A(KEYINPUT100), .ZN(new_n652));
  AND2_X1   g466(.A1(new_n575), .A2(new_n633), .ZN(new_n653));
  AND2_X1   g467(.A1(new_n256), .A2(new_n313), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n653), .A2(new_n187), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT99), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g471(.A(KEYINPUT96), .B(KEYINPUT38), .Z(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT97), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n481), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n500), .A2(new_n519), .ZN(new_n662));
  OR2_X1    g476(.A1(new_n490), .A2(new_n514), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n188), .B1(new_n663), .B2(new_n506), .ZN(new_n664));
  OAI21_X1  g478(.A(G472), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n529), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT98), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n652), .B1(new_n661), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n666), .B(KEYINPUT98), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n670), .A2(KEYINPUT100), .A3(new_n660), .A4(new_n657), .ZN(new_n671));
  XOR2_X1   g485(.A(new_n644), .B(KEYINPUT39), .Z(new_n672));
  NAND2_X1  g486(.A1(new_n413), .A2(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(new_n673), .B(KEYINPUT40), .Z(new_n674));
  NAND3_X1  g488(.A1(new_n669), .A2(new_n671), .A3(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  NAND3_X1  g490(.A1(new_n606), .A2(new_n256), .A3(new_n645), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n546), .A2(new_n634), .A3(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n649), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(new_n202), .ZN(G48));
  OAI21_X1  g495(.A(new_n188), .B1(new_n410), .B2(new_n411), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n683), .A2(new_n323), .A3(new_n412), .ZN(new_n684));
  INV_X1    g498(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n546), .A2(new_n581), .A3(new_n685), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n589), .A2(new_n591), .A3(new_n608), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XOR2_X1   g502(.A(KEYINPUT41), .B(G113), .Z(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(KEYINPUT101), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n688), .B(new_n690), .ZN(G15));
  NAND3_X1  g505(.A1(new_n625), .A2(new_n589), .A3(new_n591), .ZN(new_n692));
  NOR2_X1   g506(.A1(new_n692), .A2(new_n686), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n259), .ZN(G18));
  AOI21_X1  g508(.A(new_n653), .B1(new_n529), .B2(new_n545), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n592), .A2(new_n322), .A3(new_n695), .A4(new_n685), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G119), .ZN(G21));
  NAND3_X1  g511(.A1(new_n589), .A2(new_n591), .A3(new_n654), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n523), .A2(new_n188), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(KEYINPUT102), .ZN(new_n700));
  INV_X1    g514(.A(new_n525), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(new_n609), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n684), .A2(new_n321), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n699), .A2(KEYINPUT102), .A3(new_n524), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n702), .A2(new_n703), .A3(new_n581), .A4(new_n704), .ZN(new_n705));
  OR2_X1    g519(.A1(new_n698), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G122), .ZN(G24));
  INV_X1    g521(.A(KEYINPUT103), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n677), .B(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n634), .A3(new_n702), .A4(new_n704), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n589), .A2(new_n591), .A3(new_n685), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(new_n198), .ZN(G27));
  AND2_X1   g527(.A1(new_n709), .A2(KEYINPUT42), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  AOI22_X1  g529(.A1(new_n526), .A2(new_n528), .B1(new_n539), .B2(new_n544), .ZN(new_n716));
  OAI21_X1  g530(.A(new_n715), .B1(new_n716), .B2(new_n580), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n546), .A2(KEYINPUT104), .A3(new_n581), .ZN(new_n718));
  INV_X1    g532(.A(new_n187), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n481), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n413), .ZN(new_n721));
  INV_X1    g535(.A(new_n721), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n714), .A2(new_n717), .A3(new_n718), .A4(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n581), .A3(new_n546), .A4(new_n709), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT42), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NAND4_X1  g542(.A1(new_n722), .A2(new_n581), .A3(new_n546), .A4(new_n647), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G134), .ZN(G36));
  NAND2_X1  g544(.A1(new_n397), .A2(new_n401), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n404), .A2(new_n406), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT45), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n325), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n407), .A2(KEYINPUT45), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n737), .A2(KEYINPUT105), .ZN(new_n738));
  INV_X1    g552(.A(KEYINPUT105), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n735), .A2(new_n739), .A3(new_n736), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n326), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n412), .B1(new_n741), .B2(KEYINPUT46), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n743), .B(new_n326), .C1(new_n738), .C2(new_n740), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n323), .B(new_n672), .C1(new_n742), .C2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n481), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n187), .ZN(new_n748));
  INV_X1    g562(.A(new_n606), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n749), .A2(KEYINPUT43), .A3(new_n256), .ZN(new_n750));
  OAI21_X1  g564(.A(KEYINPUT43), .B1(new_n749), .B2(new_n256), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n701), .A2(new_n609), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT106), .B1(new_n753), .B2(new_n653), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT106), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n611), .A2(new_n755), .A3(new_n634), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n748), .B1(new_n757), .B2(KEYINPUT44), .ZN(new_n758));
  OR2_X1    g572(.A1(new_n757), .A2(KEYINPUT44), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n746), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G137), .ZN(G39));
  NAND4_X1  g575(.A1(new_n716), .A2(new_n580), .A3(new_n678), .A4(new_n720), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n323), .B1(new_n742), .B2(new_n744), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT47), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI211_X1 g579(.A(KEYINPUT47), .B(new_n323), .C1(new_n742), .C2(new_n744), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n762), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n196), .ZN(G42));
  NAND2_X1  g582(.A1(new_n683), .A2(new_n412), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n769), .B(KEYINPUT49), .Z(new_n770));
  INV_X1    g584(.A(new_n256), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n580), .A2(new_n719), .A3(new_n324), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(new_n771), .A3(new_n606), .A4(new_n772), .ZN(new_n773));
  OR3_X1    g587(.A1(new_n670), .A2(new_n773), .A3(new_n660), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n775));
  AND3_X1   g589(.A1(new_n589), .A2(new_n413), .A3(new_n591), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n716), .A2(new_n653), .A3(new_n646), .ZN(new_n777));
  AOI211_X1 g591(.A(new_n653), .B(new_n677), .C1(new_n529), .C2(new_n545), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n776), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n612), .A2(new_n634), .A3(new_n644), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n592), .A2(new_n666), .A3(new_n654), .A4(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n702), .A2(new_n634), .A3(new_n704), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n592), .A2(new_n685), .A3(new_n782), .A4(new_n709), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  AND3_X1   g598(.A1(new_n784), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT52), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n649), .B1(new_n648), .B2(new_n679), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n788), .A2(new_n712), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n789), .A2(KEYINPUT52), .A3(new_n781), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n784), .A2(KEYINPUT109), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n785), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n612), .A2(new_n580), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n747), .A2(new_n719), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n771), .A2(new_n313), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n321), .B1(new_n796), .B2(new_n607), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n794), .A2(new_n795), .A3(new_n753), .A4(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n639), .A2(new_n582), .A3(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n799), .B1(new_n723), .B2(new_n726), .ZN(new_n800));
  INV_X1    g614(.A(new_n233), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n313), .A2(new_n801), .A3(new_n644), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(new_n621), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n546), .A2(new_n634), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n721), .B1(new_n710), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(new_n729), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT108), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT108), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n782), .A2(new_n709), .B1(new_n695), .B2(new_n803), .ZN(new_n809));
  OAI211_X1 g623(.A(new_n729), .B(new_n808), .C1(new_n809), .C2(new_n721), .ZN(new_n810));
  AND3_X1   g624(.A1(new_n800), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n695), .A2(new_n322), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n812), .A2(new_n711), .B1(new_n698), .B2(new_n705), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n686), .B1(new_n692), .B2(new_n687), .ZN(new_n814));
  OAI21_X1  g628(.A(KEYINPUT107), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n716), .A2(new_n580), .A3(new_n684), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n816), .B(new_n592), .C1(new_n608), .C2(new_n625), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT107), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n696), .A3(new_n706), .A4(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n815), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n811), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(KEYINPUT110), .B(new_n775), .C1(new_n793), .C2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n800), .A2(new_n807), .A3(new_n810), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n815), .A2(new_n819), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT53), .A3(new_n791), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n822), .A2(new_n826), .ZN(new_n827));
  AOI22_X1  g641(.A1(new_n787), .A2(new_n790), .B1(KEYINPUT109), .B2(new_n784), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n828), .B2(new_n785), .ZN(new_n829));
  AOI21_X1  g643(.A(KEYINPUT110), .B1(new_n829), .B2(new_n775), .ZN(new_n830));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n827), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n791), .A2(new_n811), .A3(new_n820), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n775), .ZN(new_n833));
  NOR3_X1   g647(.A1(new_n813), .A2(new_n814), .A3(new_n775), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n834), .A2(new_n810), .A3(new_n800), .A4(new_n807), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n836), .B1(new_n828), .B2(new_n785), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n833), .A2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT111), .B1(new_n838), .B2(KEYINPUT54), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n769), .A2(new_n323), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n765), .A2(new_n766), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n841), .B2(KEYINPUT112), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n842), .B1(KEYINPUT112), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n752), .A2(new_n317), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n702), .A2(new_n581), .A3(new_n704), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n748), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n843), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n720), .A2(new_n318), .A3(new_n685), .ZN(new_n849));
  NOR3_X1   g663(.A1(new_n670), .A2(new_n580), .A3(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n771), .A3(new_n749), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n752), .A2(new_n849), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(new_n782), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(new_n846), .ZN(new_n855));
  NOR3_X1   g669(.A1(new_n660), .A2(new_n187), .A3(new_n684), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XOR2_X1   g671(.A(KEYINPUT113), .B(KEYINPUT50), .Z(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n855), .B(new_n856), .C1(new_n860), .C2(KEYINPUT50), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n859), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g676(.A(KEYINPUT51), .B1(new_n848), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n847), .B1(new_n841), .B2(new_n840), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n854), .A2(KEYINPUT114), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n866), .B1(new_n859), .B2(new_n861), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n851), .A2(new_n868), .A3(new_n853), .ZN(new_n869));
  AND4_X1   g683(.A1(new_n864), .A2(new_n865), .A3(new_n867), .A4(new_n869), .ZN(new_n870));
  AND2_X1   g684(.A1(new_n717), .A2(new_n718), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n852), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT48), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n850), .A2(new_n256), .A3(new_n606), .ZN(new_n874));
  OR2_X1    g688(.A1(new_n846), .A2(new_n711), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n873), .A2(new_n315), .A3(new_n874), .A4(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n863), .A2(new_n870), .A3(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(KEYINPUT53), .B1(new_n825), .B2(new_n791), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT52), .B1(new_n789), .B2(new_n781), .ZN(new_n879));
  AND4_X1   g693(.A1(KEYINPUT52), .A2(new_n779), .A3(new_n783), .A4(new_n781), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n792), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n784), .A2(KEYINPUT109), .A3(KEYINPUT52), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n835), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n878), .A2(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT111), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n884), .A2(new_n885), .A3(new_n886), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n831), .A2(new_n839), .A3(new_n877), .A4(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n774), .B1(new_n888), .B2(new_n889), .ZN(G75));
  NOR2_X1   g704(.A1(new_n470), .A2(new_n471), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT115), .Z(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT55), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(new_n467), .Z(new_n894));
  INV_X1    g708(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(G210), .A2(G902), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n897), .B1(new_n878), .B2(new_n883), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n896), .B1(new_n833), .B2(new_n837), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(KEYINPUT116), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n895), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n190), .A2(G952), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n894), .A2(KEYINPUT56), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n904), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(KEYINPUT117), .B1(new_n903), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT56), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n901), .B2(KEYINPUT116), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n898), .A2(new_n899), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n894), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT117), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n912), .A2(new_n913), .A3(new_n906), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n908), .A2(new_n914), .ZN(G51));
  XNOR2_X1  g729(.A(new_n838), .B(new_n886), .ZN(new_n916));
  XOR2_X1   g730(.A(new_n326), .B(KEYINPUT57), .Z(new_n917));
  OAI22_X1  g731(.A1(new_n916), .A2(new_n917), .B1(new_n411), .B2(new_n410), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n884), .A2(new_n188), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n919), .A2(new_n740), .A3(new_n738), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n904), .B1(new_n918), .B2(new_n920), .ZN(G54));
  NAND3_X1  g735(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n922));
  INV_X1    g736(.A(new_n249), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n904), .ZN(G60));
  INV_X1    g740(.A(new_n904), .ZN(new_n927));
  XOR2_X1   g741(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n928));
  NOR2_X1   g742(.A1(new_n257), .A2(new_n188), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n928), .B(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n600), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n927), .B1(new_n916), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n822), .A2(new_n826), .ZN(new_n934));
  INV_X1    g748(.A(new_n830), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n886), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n839), .A2(new_n887), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n931), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n600), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(G63));
  INV_X1    g754(.A(KEYINPUT61), .ZN(new_n941));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n884), .A2(new_n943), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n632), .B(KEYINPUT119), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n927), .B1(new_n944), .B2(new_n576), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OR2_X1    g763(.A1(new_n944), .A2(new_n576), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n950), .A2(KEYINPUT61), .A3(new_n927), .A4(new_n946), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(G66));
  INV_X1    g766(.A(G224), .ZN(new_n953));
  OAI21_X1  g767(.A(G953), .B1(new_n320), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT120), .Z(new_n955));
  NOR2_X1   g769(.A1(new_n824), .A2(new_n799), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n955), .B1(new_n956), .B2(G953), .ZN(new_n957));
  OAI21_X1  g771(.A(new_n892), .B1(G898), .B2(new_n190), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n957), .B(new_n958), .ZN(G69));
  INV_X1    g773(.A(new_n871), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n960), .A2(new_n745), .A3(new_n698), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n727), .A2(new_n729), .ZN(new_n962));
  NOR3_X1   g776(.A1(new_n767), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n760), .A2(new_n789), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(KEYINPUT124), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n760), .A2(new_n966), .A3(new_n789), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n965), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(KEYINPUT125), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n963), .A2(new_n965), .A3(new_n970), .A4(new_n967), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n969), .A2(new_n190), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n499), .B(KEYINPUT121), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n242), .A2(new_n243), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n973), .B(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n972), .B(new_n975), .C1(new_n643), .C2(new_n190), .ZN(new_n976));
  OAI21_X1  g790(.A(G953), .B1(new_n399), .B2(new_n643), .ZN(new_n977));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n796), .A2(new_n607), .ZN(new_n981));
  NOR3_X1   g795(.A1(new_n748), .A2(new_n981), .A3(new_n673), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n982), .A2(new_n581), .A3(new_n546), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n760), .A2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n760), .A2(KEYINPUT123), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n675), .A2(new_n789), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n767), .B1(new_n989), .B2(KEYINPUT62), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n675), .A2(new_n991), .A3(new_n789), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n988), .A2(new_n990), .A3(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n190), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n975), .B(KEYINPUT122), .Z(new_n995));
  AOI21_X1  g809(.A(new_n980), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AND3_X1   g810(.A1(new_n976), .A2(new_n979), .A3(new_n996), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n979), .B1(new_n976), .B2(new_n996), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(G72));
  INV_X1    g813(.A(new_n662), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n988), .A2(new_n990), .A3(new_n956), .A4(new_n992), .ZN(new_n1001));
  NAND2_X1  g815(.A1(G472), .A2(G902), .ZN(new_n1002));
  XOR2_X1   g816(.A(new_n1002), .B(KEYINPUT63), .Z(new_n1003));
  AOI21_X1  g817(.A(new_n1000), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT127), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n934), .A2(new_n935), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n500), .A2(new_n519), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1007), .A2(new_n1000), .A3(new_n1008), .A4(new_n1003), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n969), .A2(new_n956), .A3(new_n971), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1008), .B1(new_n1010), .B2(new_n1003), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1011), .A2(new_n904), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n1006), .A2(new_n1009), .A3(new_n1012), .ZN(G57));
endmodule


