

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796;

  INV_X1 U388 ( .A(n682), .ZN(n366) );
  NOR2_X1 U389 ( .A1(n646), .A2(n627), .ZN(n628) );
  NOR2_X1 U390 ( .A1(n608), .A2(n400), .ZN(n577) );
  AND2_X1 U391 ( .A1(n587), .A2(n419), .ZN(n589) );
  XOR2_X1 U392 ( .A(G140), .B(G122), .Z(n556) );
  BUF_X1 U393 ( .A(G143), .Z(n365) );
  XNOR2_X1 U394 ( .A(n510), .B(n511), .ZN(n782) );
  XNOR2_X1 U395 ( .A(n472), .B(n490), .ZN(n505) );
  XNOR2_X1 U396 ( .A(n543), .B(KEYINPUT4), .ZN(n510) );
  XNOR2_X1 U397 ( .A(KEYINPUT3), .B(G119), .ZN(n413) );
  INV_X1 U398 ( .A(G122), .ZN(n405) );
  INV_X1 U399 ( .A(G953), .ZN(n784) );
  INV_X2 U400 ( .A(G143), .ZN(n408) );
  XNOR2_X1 U401 ( .A(n367), .B(n366), .ZN(G51) );
  NAND2_X1 U402 ( .A1(n387), .A2(n483), .ZN(n367) );
  NAND2_X1 U403 ( .A1(n368), .A2(n462), .ZN(n460) );
  NAND2_X1 U404 ( .A1(n640), .A2(n376), .ZN(n368) );
  XNOR2_X2 U405 ( .A(n537), .B(n538), .ZN(n757) );
  XOR2_X1 U406 ( .A(KEYINPUT100), .B(KEYINPUT76), .Z(n507) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n509) );
  XNOR2_X1 U408 ( .A(G131), .B(n365), .ZN(n555) );
  XOR2_X1 U409 ( .A(KEYINPUT72), .B(G110), .Z(n534) );
  XNOR2_X1 U410 ( .A(n589), .B(n588), .ZN(n607) );
  NAND2_X1 U411 ( .A1(n607), .A2(n699), .ZN(n478) );
  BUF_X1 U412 ( .A(n652), .Z(n429) );
  XNOR2_X2 U413 ( .A(n586), .B(KEYINPUT1), .ZN(n631) );
  XNOR2_X1 U414 ( .A(n473), .B(n505), .ZN(n773) );
  AND2_X1 U415 ( .A1(n426), .A2(n425), .ZN(n587) );
  NAND2_X1 U416 ( .A1(n724), .A2(n624), .ZN(n719) );
  INV_X1 U417 ( .A(KEYINPUT16), .ZN(n418) );
  XNOR2_X1 U418 ( .A(n628), .B(KEYINPUT32), .ZN(n794) );
  XNOR2_X1 U419 ( .A(n655), .B(n404), .ZN(n704) );
  NOR2_X1 U420 ( .A1(n707), .A2(n698), .ZN(n585) );
  XNOR2_X1 U421 ( .A(n476), .B(n474), .ZN(n792) );
  NAND2_X1 U422 ( .A1(n398), .A2(n397), .ZN(n476) );
  AND2_X1 U423 ( .A1(n434), .A2(n623), .ZN(n707) );
  NOR2_X1 U424 ( .A1(n740), .A2(n738), .ZN(n593) );
  OR2_X1 U425 ( .A1(n634), .A2(n572), .ZN(n573) );
  INV_X1 U426 ( .A(n647), .ZN(n634) );
  OR2_X1 U427 ( .A1(n592), .A2(n591), .ZN(n738) );
  NAND2_X1 U428 ( .A1(n504), .A2(n503), .ZN(n395) );
  NAND2_X2 U429 ( .A1(n444), .A2(n441), .ZN(n586) );
  AND2_X1 U430 ( .A1(n446), .A2(n445), .ZN(n444) );
  OR2_X1 U431 ( .A1(n757), .A2(n442), .ZN(n441) );
  XNOR2_X1 U432 ( .A(n417), .B(n563), .ZN(n473) );
  XNOR2_X1 U433 ( .A(n369), .B(G137), .ZN(n487) );
  XNOR2_X1 U434 ( .A(n547), .B(n418), .ZN(n417) );
  NAND2_X1 U435 ( .A1(G214), .A2(n500), .ZN(n735) );
  XNOR2_X1 U436 ( .A(n413), .B(KEYINPUT71), .ZN(n472) );
  NAND2_X1 U437 ( .A1(n539), .A2(n443), .ZN(n442) );
  NOR2_X1 U438 ( .A1(n646), .A2(n647), .ZN(n648) );
  XNOR2_X2 U439 ( .A(n782), .B(G146), .ZN(n538) );
  INV_X1 U440 ( .A(G472), .ZN(n411) );
  NOR2_X1 U441 ( .A1(n795), .A2(n792), .ZN(n596) );
  XNOR2_X1 U442 ( .A(n578), .B(n436), .ZN(n647) );
  XNOR2_X1 U443 ( .A(n571), .B(KEYINPUT107), .ZN(n436) );
  NAND2_X1 U444 ( .A1(n449), .A2(n383), .ZN(n448) );
  NAND2_X1 U445 ( .A1(n704), .A2(n688), .ZN(n657) );
  NOR2_X1 U446 ( .A1(n598), .A2(n597), .ZN(n603) );
  XNOR2_X1 U447 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n558) );
  AND2_X1 U448 ( .A1(n415), .A2(n645), .ZN(n438) );
  XOR2_X1 U449 ( .A(G113), .B(G104), .Z(n563) );
  NAND2_X1 U450 ( .A1(n458), .A2(n453), .ZN(n452) );
  NAND2_X1 U451 ( .A1(n662), .A2(n667), .ZN(n453) );
  INV_X1 U452 ( .A(n735), .ZN(n406) );
  NAND2_X1 U453 ( .A1(n393), .A2(n391), .ZN(n652) );
  NAND2_X1 U454 ( .A1(n389), .A2(KEYINPUT0), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n635), .B(KEYINPUT33), .ZN(n636) );
  NOR2_X1 U456 ( .A1(n590), .A2(n420), .ZN(n419) );
  INV_X1 U457 ( .A(KEYINPUT111), .ZN(n402) );
  XNOR2_X1 U458 ( .A(n527), .B(n529), .ZN(n422) );
  XOR2_X1 U459 ( .A(n624), .B(KEYINPUT108), .Z(n725) );
  XNOR2_X1 U460 ( .A(n467), .B(n675), .ZN(n466) );
  NAND2_X1 U461 ( .A1(n763), .A2(G475), .ZN(n467) );
  XNOR2_X1 U462 ( .A(n399), .B(n465), .ZN(n537) );
  XNOR2_X1 U463 ( .A(n535), .B(n534), .ZN(n465) );
  XNOR2_X1 U464 ( .A(n779), .B(n536), .ZN(n399) );
  NAND2_X1 U465 ( .A1(n763), .A2(G210), .ZN(n388) );
  NAND2_X1 U466 ( .A1(n395), .A2(n371), .ZN(n394) );
  INV_X1 U467 ( .A(KEYINPUT17), .ZN(n491) );
  XOR2_X1 U468 ( .A(KEYINPUT18), .B(KEYINPUT95), .Z(n493) );
  XNOR2_X1 U469 ( .A(n611), .B(KEYINPUT38), .ZN(n736) );
  NOR2_X1 U470 ( .A1(G902), .A2(G237), .ZN(n497) );
  INV_X1 U471 ( .A(n394), .ZN(n390) );
  INV_X1 U472 ( .A(G113), .ZN(n424) );
  XNOR2_X1 U473 ( .A(KEYINPUT5), .B(KEYINPUT99), .ZN(n506) );
  XNOR2_X1 U474 ( .A(G131), .B(G134), .ZN(n511) );
  XNOR2_X1 U475 ( .A(n464), .B(G140), .ZN(n533) );
  INV_X1 U476 ( .A(G137), .ZN(n464) );
  NAND2_X1 U477 ( .A1(G234), .A2(G237), .ZN(n512) );
  NAND2_X1 U478 ( .A1(n736), .A2(n735), .ZN(n740) );
  INV_X1 U479 ( .A(n736), .ZN(n590) );
  INV_X1 U480 ( .A(G902), .ZN(n443) );
  NAND2_X1 U481 ( .A1(n447), .A2(G902), .ZN(n445) );
  XNOR2_X1 U482 ( .A(n565), .B(n433), .ZN(n672) );
  XNOR2_X1 U483 ( .A(n564), .B(n373), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n518), .B(n517), .ZN(n544) );
  INV_X1 U485 ( .A(KEYINPUT8), .ZN(n517) );
  XNOR2_X1 U486 ( .A(G128), .B(G119), .ZN(n521) );
  XOR2_X1 U487 ( .A(KEYINPUT23), .B(G110), .Z(n522) );
  NAND2_X1 U488 ( .A1(n454), .A2(n452), .ZN(n451) );
  NAND2_X1 U489 ( .A1(n666), .A2(n667), .ZN(n454) );
  XNOR2_X1 U490 ( .A(n533), .B(n463), .ZN(n779) );
  INV_X1 U491 ( .A(KEYINPUT97), .ZN(n463) );
  XNOR2_X1 U492 ( .A(n410), .B(n409), .ZN(n535) );
  INV_X1 U493 ( .A(G107), .ZN(n409) );
  XNOR2_X1 U494 ( .A(G101), .B(G104), .ZN(n410) );
  XNOR2_X1 U495 ( .A(n432), .B(n431), .ZN(n717) );
  INV_X1 U496 ( .A(KEYINPUT78), .ZN(n431) );
  INV_X1 U497 ( .A(n580), .ZN(n425) );
  INV_X1 U498 ( .A(KEYINPUT30), .ZN(n427) );
  XNOR2_X1 U499 ( .A(n475), .B(KEYINPUT42), .ZN(n474) );
  INV_X1 U500 ( .A(KEYINPUT112), .ZN(n475) );
  INV_X1 U501 ( .A(KEYINPUT40), .ZN(n477) );
  INV_X1 U502 ( .A(KEYINPUT35), .ZN(n459) );
  INV_X1 U503 ( .A(KEYINPUT31), .ZN(n404) );
  AND2_X1 U504 ( .A1(n622), .A2(n375), .ZN(n694) );
  AND2_X1 U505 ( .A1(n720), .A2(n470), .ZN(n469) );
  INV_X1 U506 ( .A(n725), .ZN(n470) );
  XNOR2_X1 U507 ( .A(n479), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U508 ( .A1(n480), .A2(n483), .ZN(n479) );
  XNOR2_X1 U509 ( .A(n481), .B(n382), .ZN(n480) );
  NAND2_X1 U510 ( .A1(n466), .A2(n483), .ZN(n428) );
  XNOR2_X1 U511 ( .A(n482), .B(KEYINPUT121), .ZN(G54) );
  NAND2_X1 U512 ( .A1(n484), .A2(n483), .ZN(n482) );
  XNOR2_X1 U513 ( .A(n485), .B(n381), .ZN(n484) );
  XNOR2_X1 U514 ( .A(n388), .B(n380), .ZN(n387) );
  AND2_X1 U515 ( .A1(G210), .A2(n557), .ZN(n369) );
  XOR2_X2 U516 ( .A(G146), .B(G125), .Z(n370) );
  OR2_X1 U517 ( .A1(n617), .A2(n616), .ZN(n371) );
  XOR2_X1 U518 ( .A(KEYINPUT82), .B(n669), .Z(n372) );
  XOR2_X1 U519 ( .A(n556), .B(n555), .Z(n373) );
  XOR2_X1 U520 ( .A(G134), .B(G116), .Z(n374) );
  AND2_X1 U521 ( .A1(n722), .A2(n720), .ZN(n375) );
  AND2_X1 U522 ( .A1(n642), .A2(KEYINPUT34), .ZN(n376) );
  INV_X1 U523 ( .A(n623), .ZN(n720) );
  AND2_X1 U524 ( .A1(n711), .A2(n372), .ZN(n377) );
  AND2_X1 U525 ( .A1(n642), .A2(n638), .ZN(n378) );
  INV_X1 U526 ( .A(n724), .ZN(n430) );
  XOR2_X1 U527 ( .A(n576), .B(KEYINPUT92), .Z(n379) );
  XNOR2_X1 U528 ( .A(n681), .B(n680), .ZN(n380) );
  XOR2_X1 U529 ( .A(n757), .B(n758), .Z(n381) );
  XOR2_X1 U530 ( .A(n685), .B(KEYINPUT113), .Z(n382) );
  XOR2_X1 U531 ( .A(G902), .B(KEYINPUT15), .Z(n663) );
  AND2_X1 U532 ( .A1(n458), .A2(n667), .ZN(n383) );
  XOR2_X1 U533 ( .A(n661), .B(n660), .Z(n384) );
  AND2_X1 U534 ( .A1(n663), .A2(KEYINPUT64), .ZN(n385) );
  XOR2_X1 U535 ( .A(n676), .B(KEYINPUT69), .Z(n386) );
  INV_X1 U536 ( .A(n767), .ZN(n483) );
  NAND2_X1 U537 ( .A1(n390), .A2(n396), .ZN(n389) );
  NAND2_X1 U538 ( .A1(n392), .A2(n396), .ZN(n391) );
  NOR2_X1 U539 ( .A1(n394), .A2(KEYINPUT0), .ZN(n392) );
  NAND2_X1 U540 ( .A1(n396), .A2(n395), .ZN(n618) );
  NAND2_X1 U541 ( .A1(n502), .A2(n501), .ZN(n396) );
  INV_X1 U542 ( .A(n750), .ZN(n397) );
  INV_X1 U543 ( .A(n594), .ZN(n398) );
  NAND2_X1 U544 ( .A1(n686), .A2(n658), .ZN(n468) );
  NAND2_X1 U545 ( .A1(n471), .A2(n469), .ZN(n686) );
  NOR2_X1 U546 ( .A1(n794), .A2(n694), .ZN(n644) );
  NOR2_X2 U547 ( .A1(n653), .A2(n634), .ZN(n637) );
  BUF_X1 U548 ( .A(n611), .Z(n400) );
  INV_X1 U549 ( .A(n401), .ZN(n639) );
  NOR2_X1 U550 ( .A1(n751), .A2(n429), .ZN(n401) );
  NAND2_X1 U551 ( .A1(n757), .A2(n447), .ZN(n446) );
  NAND2_X1 U552 ( .A1(n456), .A2(n385), .ZN(n455) );
  AND2_X2 U553 ( .A1(n713), .A2(n768), .ZN(n456) );
  XNOR2_X2 U554 ( .A(n403), .B(n402), .ZN(n594) );
  NAND2_X1 U555 ( .A1(n541), .A2(n540), .ZN(n403) );
  NOR2_X1 U556 ( .A1(n430), .A2(n738), .ZN(n619) );
  XNOR2_X1 U557 ( .A(n510), .B(n495), .ZN(n414) );
  XNOR2_X2 U558 ( .A(n405), .B(G107), .ZN(n547) );
  OR2_X1 U559 ( .A1(n578), .A2(n406), .ZN(n579) );
  XNOR2_X1 U560 ( .A(n505), .B(n423), .ZN(n488) );
  NAND2_X1 U561 ( .A1(n407), .A2(n659), .ZN(n440) );
  XNOR2_X1 U562 ( .A(n468), .B(KEYINPUT109), .ZN(n407) );
  XNOR2_X1 U563 ( .A(n414), .B(n496), .ZN(n416) );
  XNOR2_X2 U564 ( .A(n408), .B(G128), .ZN(n543) );
  NAND2_X1 U565 ( .A1(n793), .A2(KEYINPUT44), .ZN(n659) );
  XNOR2_X2 U566 ( .A(n460), .B(n459), .ZN(n793) );
  XNOR2_X2 U567 ( .A(n637), .B(n636), .ZN(n751) );
  XNOR2_X2 U568 ( .A(n412), .B(n411), .ZN(n578) );
  OR2_X2 U569 ( .A1(n684), .A2(G902), .ZN(n412) );
  NOR2_X2 U570 ( .A1(n572), .A2(n722), .ZN(n421) );
  XNOR2_X1 U571 ( .A(n508), .B(n424), .ZN(n423) );
  XNOR2_X1 U572 ( .A(n648), .B(KEYINPUT90), .ZN(n471) );
  XNOR2_X1 U573 ( .A(n630), .B(KEYINPUT65), .ZN(n415) );
  AND2_X1 U574 ( .A1(n670), .A2(n377), .ZN(n435) );
  XNOR2_X1 U575 ( .A(n416), .B(n773), .ZN(n677) );
  NAND2_X2 U576 ( .A1(n450), .A2(n448), .ZN(n457) );
  INV_X1 U577 ( .A(n651), .ZN(n420) );
  NOR2_X2 U578 ( .A1(n618), .A2(n594), .ZN(n542) );
  XOR2_X2 U579 ( .A(KEYINPUT81), .B(n542), .Z(n700) );
  BUF_X2 U580 ( .A(n578), .Z(n722) );
  XNOR2_X1 U581 ( .A(n421), .B(KEYINPUT28), .ZN(n541) );
  XNOR2_X2 U582 ( .A(n528), .B(n422), .ZN(n624) );
  XNOR2_X1 U583 ( .A(n593), .B(KEYINPUT41), .ZN(n750) );
  XNOR2_X1 U584 ( .A(n579), .B(n427), .ZN(n426) );
  XNOR2_X1 U585 ( .A(n428), .B(n386), .ZN(G60) );
  XNOR2_X2 U586 ( .A(n621), .B(KEYINPUT22), .ZN(n646) );
  NAND2_X1 U587 ( .A1(n435), .A2(n768), .ZN(n432) );
  XNOR2_X1 U588 ( .A(n778), .B(n489), .ZN(n523) );
  XNOR2_X1 U589 ( .A(n577), .B(n379), .ZN(n434) );
  NOR2_X2 U590 ( .A1(n604), .A2(n605), .ZN(n606) );
  XNOR2_X2 U591 ( .A(n437), .B(n384), .ZN(n768) );
  NAND2_X1 U592 ( .A1(n439), .A2(n438), .ZN(n437) );
  XNOR2_X1 U593 ( .A(n440), .B(KEYINPUT91), .ZN(n439) );
  INV_X1 U594 ( .A(n539), .ZN(n447) );
  INV_X1 U595 ( .A(n456), .ZN(n449) );
  AND2_X2 U596 ( .A1(n455), .A2(n451), .ZN(n450) );
  AND2_X4 U597 ( .A1(n457), .A2(n671), .ZN(n763) );
  INV_X1 U598 ( .A(n666), .ZN(n458) );
  NAND2_X1 U599 ( .A1(n639), .A2(n378), .ZN(n462) );
  XNOR2_X2 U600 ( .A(n478), .B(n477), .ZN(n795) );
  NAND2_X1 U601 ( .A1(n763), .A2(G472), .ZN(n481) );
  NAND2_X1 U602 ( .A1(n763), .A2(G469), .ZN(n485) );
  XNOR2_X1 U603 ( .A(n486), .B(n538), .ZN(n684) );
  XNOR2_X1 U604 ( .A(n488), .B(n487), .ZN(n486) );
  XOR2_X2 U605 ( .A(n370), .B(KEYINPUT10), .Z(n778) );
  XOR2_X1 U606 ( .A(n522), .B(n521), .Z(n489) );
  INV_X1 U607 ( .A(KEYINPUT46), .ZN(n595) );
  XNOR2_X1 U608 ( .A(n596), .B(n595), .ZN(n597) );
  XNOR2_X1 U609 ( .A(n492), .B(n491), .ZN(n494) );
  XNOR2_X1 U610 ( .A(n494), .B(n493), .ZN(n496) );
  INV_X1 U611 ( .A(KEYINPUT36), .ZN(n576) );
  XNOR2_X1 U612 ( .A(n547), .B(n374), .ZN(n548) );
  XNOR2_X1 U613 ( .A(KEYINPUT89), .B(KEYINPUT39), .ZN(n588) );
  XNOR2_X1 U614 ( .A(n523), .B(n524), .ZN(n765) );
  NOR2_X1 U615 ( .A1(G952), .A2(n784), .ZN(n767) );
  XNOR2_X1 U616 ( .A(G116), .B(G101), .ZN(n490) );
  NAND2_X1 U617 ( .A1(G224), .A2(n784), .ZN(n492) );
  XNOR2_X1 U618 ( .A(n534), .B(n370), .ZN(n495) );
  NOR2_X1 U619 ( .A1(n663), .A2(n677), .ZN(n499) );
  XNOR2_X1 U620 ( .A(n497), .B(KEYINPUT75), .ZN(n500) );
  NAND2_X1 U621 ( .A1(G210), .A2(n500), .ZN(n498) );
  XNOR2_X1 U622 ( .A(n499), .B(n498), .ZN(n575) );
  NAND2_X1 U623 ( .A1(n575), .A2(n735), .ZN(n504) );
  INV_X1 U624 ( .A(n504), .ZN(n502) );
  XOR2_X1 U625 ( .A(KEYINPUT19), .B(KEYINPUT68), .Z(n503) );
  INV_X1 U626 ( .A(n503), .ZN(n501) );
  XNOR2_X1 U627 ( .A(n507), .B(n506), .ZN(n508) );
  XOR2_X1 U628 ( .A(KEYINPUT77), .B(n509), .Z(n557) );
  XNOR2_X1 U629 ( .A(n512), .B(KEYINPUT14), .ZN(n513) );
  NAND2_X1 U630 ( .A1(G952), .A2(n513), .ZN(n749) );
  NOR2_X1 U631 ( .A1(G953), .A2(n749), .ZN(n617) );
  NAND2_X1 U632 ( .A1(G902), .A2(n513), .ZN(n514) );
  XOR2_X1 U633 ( .A(KEYINPUT96), .B(n514), .Z(n515) );
  NAND2_X1 U634 ( .A1(G953), .A2(n515), .ZN(n615) );
  NOR2_X1 U635 ( .A1(G900), .A2(n615), .ZN(n516) );
  NOR2_X1 U636 ( .A1(n617), .A2(n516), .ZN(n580) );
  XOR2_X1 U637 ( .A(n533), .B(KEYINPUT24), .Z(n520) );
  NAND2_X1 U638 ( .A1(n784), .A2(G234), .ZN(n518) );
  NAND2_X1 U639 ( .A1(G221), .A2(n544), .ZN(n519) );
  XNOR2_X1 U640 ( .A(n520), .B(n519), .ZN(n524) );
  NOR2_X1 U641 ( .A1(G902), .A2(n765), .ZN(n528) );
  INV_X1 U642 ( .A(n663), .ZN(n662) );
  NAND2_X1 U643 ( .A1(n662), .A2(G234), .ZN(n526) );
  XNOR2_X1 U644 ( .A(KEYINPUT98), .B(KEYINPUT20), .ZN(n525) );
  XNOR2_X1 U645 ( .A(n526), .B(n525), .ZN(n530) );
  NAND2_X1 U646 ( .A1(G217), .A2(n530), .ZN(n527) );
  XOR2_X1 U647 ( .A(KEYINPUT79), .B(KEYINPUT25), .Z(n529) );
  NOR2_X1 U648 ( .A1(n580), .A2(n624), .ZN(n532) );
  NAND2_X1 U649 ( .A1(n530), .A2(G221), .ZN(n531) );
  XOR2_X1 U650 ( .A(KEYINPUT21), .B(n531), .Z(n724) );
  NAND2_X1 U651 ( .A1(n532), .A2(n724), .ZN(n572) );
  AND2_X1 U652 ( .A1(G227), .A2(n784), .ZN(n536) );
  XNOR2_X1 U653 ( .A(KEYINPUT70), .B(G469), .ZN(n539) );
  INV_X1 U654 ( .A(n586), .ZN(n540) );
  XNOR2_X1 U655 ( .A(KEYINPUT9), .B(KEYINPUT106), .ZN(n551) );
  XOR2_X1 U656 ( .A(n543), .B(KEYINPUT7), .Z(n546) );
  NAND2_X1 U657 ( .A1(G217), .A2(n544), .ZN(n545) );
  XNOR2_X1 U658 ( .A(n546), .B(n545), .ZN(n549) );
  XNOR2_X1 U659 ( .A(n549), .B(n548), .ZN(n550) );
  XNOR2_X1 U660 ( .A(n551), .B(n550), .ZN(n759) );
  NOR2_X1 U661 ( .A1(G902), .A2(n759), .ZN(n552) );
  XOR2_X1 U662 ( .A(G478), .B(n552), .Z(n591) );
  INV_X1 U663 ( .A(n591), .ZN(n568) );
  XOR2_X1 U664 ( .A(KEYINPUT105), .B(KEYINPUT13), .Z(n554) );
  XNOR2_X1 U665 ( .A(KEYINPUT104), .B(G475), .ZN(n553) );
  XNOR2_X1 U666 ( .A(n554), .B(n553), .ZN(n567) );
  NAND2_X1 U667 ( .A1(G214), .A2(n557), .ZN(n561) );
  XOR2_X1 U668 ( .A(KEYINPUT12), .B(KEYINPUT103), .Z(n559) );
  XNOR2_X1 U669 ( .A(n559), .B(n558), .ZN(n560) );
  XNOR2_X1 U670 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U671 ( .A(n562), .B(KEYINPUT11), .Z(n565) );
  XNOR2_X1 U672 ( .A(n563), .B(n778), .ZN(n564) );
  NOR2_X1 U673 ( .A1(G902), .A2(n672), .ZN(n566) );
  XNOR2_X1 U674 ( .A(n567), .B(n566), .ZN(n592) );
  NAND2_X1 U675 ( .A1(n568), .A2(n592), .ZN(n702) );
  INV_X1 U676 ( .A(n702), .ZN(n699) );
  NOR2_X1 U677 ( .A1(n568), .A2(n592), .ZN(n695) );
  NOR2_X1 U678 ( .A1(n699), .A2(n695), .ZN(n741) );
  INV_X1 U679 ( .A(n741), .ZN(n599) );
  XNOR2_X1 U680 ( .A(n599), .B(KEYINPUT84), .ZN(n656) );
  AND2_X1 U681 ( .A1(n700), .A2(n656), .ZN(n569) );
  NOR2_X1 U682 ( .A1(KEYINPUT83), .A2(n569), .ZN(n570) );
  NOR2_X1 U683 ( .A1(KEYINPUT47), .A2(n570), .ZN(n605) );
  INV_X1 U684 ( .A(n631), .ZN(n623) );
  INV_X1 U685 ( .A(KEYINPUT6), .ZN(n571) );
  NOR2_X1 U686 ( .A1(n702), .A2(n573), .ZN(n574) );
  NAND2_X1 U687 ( .A1(n574), .A2(n735), .ZN(n608) );
  INV_X1 U688 ( .A(n575), .ZN(n611) );
  INV_X1 U689 ( .A(n722), .ZN(n649) );
  NAND2_X1 U690 ( .A1(n591), .A2(n592), .ZN(n641) );
  OR2_X1 U691 ( .A1(n400), .A2(n719), .ZN(n581) );
  NOR2_X1 U692 ( .A1(n641), .A2(n581), .ZN(n582) );
  NAND2_X1 U693 ( .A1(n587), .A2(n582), .ZN(n583) );
  NOR2_X1 U694 ( .A1(n586), .A2(n583), .ZN(n698) );
  NAND2_X1 U695 ( .A1(KEYINPUT83), .A2(n599), .ZN(n584) );
  NAND2_X1 U696 ( .A1(n585), .A2(n584), .ZN(n598) );
  NOR2_X1 U697 ( .A1(n586), .A2(n719), .ZN(n651) );
  OR2_X1 U698 ( .A1(KEYINPUT83), .A2(n599), .ZN(n600) );
  NAND2_X1 U699 ( .A1(n600), .A2(n700), .ZN(n601) );
  NAND2_X1 U700 ( .A1(n601), .A2(KEYINPUT47), .ZN(n602) );
  NAND2_X1 U701 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U702 ( .A(n606), .B(KEYINPUT48), .ZN(n670) );
  NAND2_X1 U703 ( .A1(n695), .A2(n607), .ZN(n668) );
  INV_X1 U704 ( .A(n668), .ZN(n710) );
  OR2_X1 U705 ( .A1(n623), .A2(n608), .ZN(n609) );
  XNOR2_X1 U706 ( .A(n609), .B(KEYINPUT110), .ZN(n610) );
  XNOR2_X1 U707 ( .A(n610), .B(KEYINPUT43), .ZN(n612) );
  NAND2_X1 U708 ( .A1(n612), .A2(n400), .ZN(n711) );
  INV_X1 U709 ( .A(n711), .ZN(n613) );
  NOR2_X1 U710 ( .A1(n710), .A2(n613), .ZN(n614) );
  AND2_X2 U711 ( .A1(n670), .A2(n614), .ZN(n713) );
  NOR2_X1 U712 ( .A1(n615), .A2(G898), .ZN(n616) );
  INV_X1 U713 ( .A(n652), .ZN(n620) );
  NAND2_X1 U714 ( .A1(n620), .A2(n619), .ZN(n621) );
  NOR2_X1 U715 ( .A1(n646), .A2(n624), .ZN(n622) );
  NAND2_X1 U716 ( .A1(n634), .A2(n725), .ZN(n625) );
  NOR2_X1 U717 ( .A1(n720), .A2(n625), .ZN(n626) );
  XOR2_X1 U718 ( .A(KEYINPUT80), .B(n626), .Z(n627) );
  INV_X1 U719 ( .A(KEYINPUT44), .ZN(n629) );
  NOR2_X1 U720 ( .A1(n644), .A2(n629), .ZN(n630) );
  NOR2_X1 U721 ( .A1(n719), .A2(n631), .ZN(n633) );
  INV_X1 U722 ( .A(KEYINPUT74), .ZN(n632) );
  XNOR2_X1 U723 ( .A(n633), .B(n632), .ZN(n653) );
  INV_X1 U724 ( .A(KEYINPUT73), .ZN(n635) );
  INV_X1 U725 ( .A(KEYINPUT34), .ZN(n638) );
  NOR2_X1 U726 ( .A1(n429), .A2(n751), .ZN(n640) );
  INV_X1 U727 ( .A(n641), .ZN(n642) );
  NOR2_X1 U728 ( .A1(n793), .A2(KEYINPUT44), .ZN(n643) );
  NAND2_X1 U729 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U730 ( .A1(n649), .A2(n429), .ZN(n650) );
  NAND2_X1 U731 ( .A1(n651), .A2(n650), .ZN(n688) );
  INV_X1 U732 ( .A(n429), .ZN(n654) );
  NOR2_X1 U733 ( .A1(n653), .A2(n722), .ZN(n731) );
  NAND2_X1 U734 ( .A1(n654), .A2(n731), .ZN(n655) );
  NAND2_X1 U735 ( .A1(n657), .A2(n656), .ZN(n658) );
  INV_X1 U736 ( .A(KEYINPUT87), .ZN(n661) );
  INV_X1 U737 ( .A(KEYINPUT45), .ZN(n660) );
  XNOR2_X1 U738 ( .A(n663), .B(KEYINPUT86), .ZN(n664) );
  NAND2_X1 U739 ( .A1(n664), .A2(KEYINPUT2), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n665), .B(KEYINPUT67), .ZN(n666) );
  INV_X1 U741 ( .A(KEYINPUT64), .ZN(n667) );
  NAND2_X1 U742 ( .A1(KEYINPUT2), .A2(n668), .ZN(n669) );
  INV_X1 U743 ( .A(n717), .ZN(n671) );
  XOR2_X1 U744 ( .A(KEYINPUT66), .B(KEYINPUT59), .Z(n674) );
  XNOR2_X1 U745 ( .A(n672), .B(KEYINPUT122), .ZN(n673) );
  XOR2_X1 U746 ( .A(n674), .B(n673), .Z(n675) );
  INV_X1 U747 ( .A(KEYINPUT60), .ZN(n676) );
  XNOR2_X1 U748 ( .A(KEYINPUT120), .B(KEYINPUT55), .ZN(n679) );
  XNOR2_X1 U749 ( .A(n677), .B(KEYINPUT94), .ZN(n678) );
  XNOR2_X1 U750 ( .A(n679), .B(n678), .ZN(n681) );
  XOR2_X1 U751 ( .A(KEYINPUT93), .B(KEYINPUT54), .Z(n680) );
  XNOR2_X1 U752 ( .A(KEYINPUT56), .B(KEYINPUT88), .ZN(n682) );
  XOR2_X1 U753 ( .A(n684), .B(KEYINPUT62), .Z(n685) );
  XNOR2_X1 U754 ( .A(G101), .B(n686), .ZN(G3) );
  NOR2_X1 U755 ( .A1(n702), .A2(n688), .ZN(n687) );
  XOR2_X1 U756 ( .A(G104), .B(n687), .Z(G6) );
  INV_X1 U757 ( .A(n695), .ZN(n705) );
  NOR2_X1 U758 ( .A1(n705), .A2(n688), .ZN(n693) );
  XOR2_X1 U759 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n690) );
  XNOR2_X1 U760 ( .A(G107), .B(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U761 ( .A(n690), .B(n689), .ZN(n691) );
  XNOR2_X1 U762 ( .A(KEYINPUT27), .B(n691), .ZN(n692) );
  XNOR2_X1 U763 ( .A(n693), .B(n692), .ZN(G9) );
  XOR2_X1 U764 ( .A(n694), .B(G110), .Z(G12) );
  XOR2_X1 U765 ( .A(G128), .B(KEYINPUT29), .Z(n697) );
  NAND2_X1 U766 ( .A1(n695), .A2(n700), .ZN(n696) );
  XNOR2_X1 U767 ( .A(n697), .B(n696), .ZN(G30) );
  XOR2_X1 U768 ( .A(n365), .B(n698), .Z(G45) );
  NAND2_X1 U769 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(G146), .ZN(G48) );
  NOR2_X1 U771 ( .A1(n702), .A2(n704), .ZN(n703) );
  XOR2_X1 U772 ( .A(G113), .B(n703), .Z(G15) );
  NOR2_X1 U773 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U774 ( .A(G116), .B(n706), .Z(G18) );
  XNOR2_X1 U775 ( .A(n707), .B(KEYINPUT116), .ZN(n708) );
  XNOR2_X1 U776 ( .A(n708), .B(KEYINPUT37), .ZN(n709) );
  XNOR2_X1 U777 ( .A(G125), .B(n709), .ZN(G27) );
  XOR2_X1 U778 ( .A(G134), .B(n710), .Z(G36) );
  XNOR2_X1 U779 ( .A(G140), .B(n711), .ZN(G42) );
  NOR2_X1 U780 ( .A1(KEYINPUT2), .A2(n768), .ZN(n712) );
  XNOR2_X1 U781 ( .A(n712), .B(KEYINPUT85), .ZN(n715) );
  OR2_X1 U782 ( .A1(n713), .A2(KEYINPUT2), .ZN(n714) );
  NAND2_X1 U783 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U785 ( .A1(G953), .A2(n718), .ZN(n755) );
  NAND2_X1 U786 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U787 ( .A(n721), .B(KEYINPUT50), .ZN(n723) );
  NAND2_X1 U788 ( .A1(n723), .A2(n722), .ZN(n728) );
  NAND2_X1 U789 ( .A1(n430), .A2(n725), .ZN(n726) );
  XNOR2_X1 U790 ( .A(KEYINPUT49), .B(n726), .ZN(n727) );
  NOR2_X1 U791 ( .A1(n728), .A2(n727), .ZN(n729) );
  XOR2_X1 U792 ( .A(KEYINPUT117), .B(n729), .Z(n730) );
  NOR2_X1 U793 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U794 ( .A(KEYINPUT51), .B(n732), .Z(n733) );
  XNOR2_X1 U795 ( .A(n733), .B(KEYINPUT118), .ZN(n734) );
  NOR2_X1 U796 ( .A1(n750), .A2(n734), .ZN(n746) );
  NOR2_X1 U797 ( .A1(n736), .A2(n735), .ZN(n737) );
  NOR2_X1 U798 ( .A1(n738), .A2(n737), .ZN(n739) );
  XOR2_X1 U799 ( .A(KEYINPUT119), .B(n739), .Z(n743) );
  NOR2_X1 U800 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U801 ( .A1(n743), .A2(n742), .ZN(n744) );
  NOR2_X1 U802 ( .A1(n751), .A2(n744), .ZN(n745) );
  NOR2_X1 U803 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U804 ( .A(n747), .B(KEYINPUT52), .ZN(n748) );
  NOR2_X1 U805 ( .A1(n749), .A2(n748), .ZN(n753) );
  NOR2_X1 U806 ( .A1(n751), .A2(n750), .ZN(n752) );
  NOR2_X1 U807 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U808 ( .A1(n755), .A2(n754), .ZN(n756) );
  XOR2_X1 U809 ( .A(KEYINPUT53), .B(n756), .Z(G75) );
  XOR2_X1 U810 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n758) );
  XOR2_X1 U811 ( .A(n759), .B(KEYINPUT123), .Z(n761) );
  NAND2_X1 U812 ( .A1(n763), .A2(G478), .ZN(n760) );
  XNOR2_X1 U813 ( .A(n761), .B(n760), .ZN(n762) );
  NOR2_X1 U814 ( .A1(n767), .A2(n762), .ZN(G63) );
  NAND2_X1 U815 ( .A1(G217), .A2(n763), .ZN(n764) );
  XNOR2_X1 U816 ( .A(n765), .B(n764), .ZN(n766) );
  NOR2_X1 U817 ( .A1(n767), .A2(n766), .ZN(G66) );
  NAND2_X1 U818 ( .A1(n784), .A2(n768), .ZN(n772) );
  NAND2_X1 U819 ( .A1(G953), .A2(G224), .ZN(n769) );
  XNOR2_X1 U820 ( .A(KEYINPUT61), .B(n769), .ZN(n770) );
  NAND2_X1 U821 ( .A1(n770), .A2(G898), .ZN(n771) );
  NAND2_X1 U822 ( .A1(n772), .A2(n771), .ZN(n777) );
  XNOR2_X1 U823 ( .A(n773), .B(G110), .ZN(n775) );
  NOR2_X1 U824 ( .A1(n784), .A2(G898), .ZN(n774) );
  NOR2_X1 U825 ( .A1(n775), .A2(n774), .ZN(n776) );
  XNOR2_X1 U826 ( .A(n777), .B(n776), .ZN(G69) );
  XOR2_X1 U827 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n781) );
  XNOR2_X1 U828 ( .A(n779), .B(n778), .ZN(n780) );
  XNOR2_X1 U829 ( .A(n781), .B(n780), .ZN(n783) );
  XOR2_X1 U830 ( .A(n783), .B(n782), .Z(n786) );
  XOR2_X1 U831 ( .A(n713), .B(n786), .Z(n785) );
  NAND2_X1 U832 ( .A1(n785), .A2(n784), .ZN(n790) );
  XNOR2_X1 U833 ( .A(G227), .B(n786), .ZN(n787) );
  NAND2_X1 U834 ( .A1(n787), .A2(G900), .ZN(n788) );
  NAND2_X1 U835 ( .A1(G953), .A2(n788), .ZN(n789) );
  NAND2_X1 U836 ( .A1(n790), .A2(n789), .ZN(n791) );
  XNOR2_X1 U837 ( .A(KEYINPUT126), .B(n791), .ZN(G72) );
  XOR2_X1 U838 ( .A(n792), .B(G137), .Z(G39) );
  XOR2_X1 U839 ( .A(n793), .B(G122), .Z(G24) );
  XOR2_X1 U840 ( .A(n794), .B(G119), .Z(G21) );
  XNOR2_X1 U841 ( .A(G131), .B(KEYINPUT127), .ZN(n796) );
  XNOR2_X1 U842 ( .A(n796), .B(n795), .ZN(G33) );
endmodule

