

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X2 U551 ( .A(n647), .ZN(n664) );
  AND2_X2 U552 ( .A1(n527), .A2(G2104), .ZN(n892) );
  NOR2_X2 U553 ( .A1(n636), .A2(n635), .ZN(n637) );
  OR2_X1 U554 ( .A1(n707), .A2(n706), .ZN(n517) );
  BUF_X1 U555 ( .A(n714), .Z(n715) );
  NOR2_X1 U556 ( .A1(n643), .A2(n642), .ZN(n646) );
  AND2_X1 U557 ( .A1(n741), .A2(n755), .ZN(n518) );
  INV_X1 U558 ( .A(KEYINPUT99), .ZN(n644) );
  XNOR2_X1 U559 ( .A(n644), .B(KEYINPUT29), .ZN(n645) );
  NAND2_X1 U560 ( .A1(n662), .A2(n661), .ZN(n672) );
  XNOR2_X1 U561 ( .A(n671), .B(KEYINPUT32), .ZN(n693) );
  INV_X1 U562 ( .A(n1001), .ZN(n689) );
  OR2_X1 U563 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U564 ( .A1(G164), .A2(G1384), .ZN(n709) );
  XNOR2_X1 U565 ( .A(n521), .B(KEYINPUT66), .ZN(n522) );
  XNOR2_X1 U566 ( .A(n523), .B(n522), .ZN(n714) );
  NOR2_X1 U567 ( .A1(n742), .A2(n518), .ZN(n743) );
  INV_X1 U568 ( .A(G651), .ZN(n541) );
  NOR2_X1 U569 ( .A1(G543), .A2(G651), .ZN(n797) );
  XNOR2_X1 U570 ( .A(KEYINPUT15), .B(n622), .ZN(n803) );
  NOR2_X1 U571 ( .A1(n577), .A2(G651), .ZN(n793) );
  NOR2_X2 U572 ( .A1(n531), .A2(n530), .ZN(G160) );
  INV_X1 U573 ( .A(G2105), .ZN(n527) );
  NAND2_X1 U574 ( .A1(G101), .A2(n892), .ZN(n519) );
  XNOR2_X1 U575 ( .A(n519), .B(KEYINPUT23), .ZN(n520) );
  XNOR2_X1 U576 ( .A(KEYINPUT65), .B(n520), .ZN(n526) );
  NOR2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  INV_X1 U578 ( .A(KEYINPUT17), .ZN(n521) );
  NAND2_X1 U579 ( .A1(n714), .A2(G137), .ZN(n524) );
  XOR2_X1 U580 ( .A(n524), .B(KEYINPUT67), .Z(n525) );
  NAND2_X1 U581 ( .A1(n526), .A2(n525), .ZN(n531) );
  AND2_X1 U582 ( .A1(G2104), .A2(G2105), .ZN(n897) );
  NAND2_X1 U583 ( .A1(G113), .A2(n897), .ZN(n529) );
  NOR2_X1 U584 ( .A1(G2104), .A2(n527), .ZN(n895) );
  NAND2_X1 U585 ( .A1(G125), .A2(n895), .ZN(n528) );
  NAND2_X1 U586 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U587 ( .A1(n892), .A2(G102), .ZN(n533) );
  NAND2_X1 U588 ( .A1(G138), .A2(n714), .ZN(n532) );
  NAND2_X1 U589 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U590 ( .A(n534), .B(KEYINPUT82), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G114), .A2(n897), .ZN(n536) );
  NAND2_X1 U592 ( .A1(G126), .A2(n895), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n538), .A2(n537), .ZN(G164) );
  NOR2_X1 U595 ( .A1(G543), .A2(n541), .ZN(n539) );
  XOR2_X1 U596 ( .A(KEYINPUT68), .B(n539), .Z(n540) );
  XNOR2_X1 U597 ( .A(KEYINPUT1), .B(n540), .ZN(n794) );
  AND2_X1 U598 ( .A1(G65), .A2(n794), .ZN(n545) );
  NAND2_X1 U599 ( .A1(G91), .A2(n797), .ZN(n543) );
  XOR2_X1 U600 ( .A(KEYINPUT0), .B(G543), .Z(n577) );
  NOR2_X1 U601 ( .A1(n577), .A2(n541), .ZN(n798) );
  NAND2_X1 U602 ( .A1(G78), .A2(n798), .ZN(n542) );
  NAND2_X1 U603 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U604 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U605 ( .A1(n793), .A2(G53), .ZN(n546) );
  NAND2_X1 U606 ( .A1(n547), .A2(n546), .ZN(G299) );
  NAND2_X1 U607 ( .A1(n793), .A2(G52), .ZN(n549) );
  NAND2_X1 U608 ( .A1(G64), .A2(n794), .ZN(n548) );
  NAND2_X1 U609 ( .A1(n549), .A2(n548), .ZN(n554) );
  NAND2_X1 U610 ( .A1(G90), .A2(n797), .ZN(n551) );
  NAND2_X1 U611 ( .A1(G77), .A2(n798), .ZN(n550) );
  NAND2_X1 U612 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U613 ( .A(KEYINPUT9), .B(n552), .Z(n553) );
  NOR2_X1 U614 ( .A1(n554), .A2(n553), .ZN(G171) );
  NAND2_X1 U615 ( .A1(n797), .A2(G89), .ZN(n555) );
  XNOR2_X1 U616 ( .A(n555), .B(KEYINPUT4), .ZN(n557) );
  NAND2_X1 U617 ( .A1(G76), .A2(n798), .ZN(n556) );
  NAND2_X1 U618 ( .A1(n557), .A2(n556), .ZN(n558) );
  XNOR2_X1 U619 ( .A(KEYINPUT5), .B(n558), .ZN(n564) );
  NAND2_X1 U620 ( .A1(n793), .A2(G51), .ZN(n560) );
  NAND2_X1 U621 ( .A1(G63), .A2(n794), .ZN(n559) );
  NAND2_X1 U622 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U623 ( .A(KEYINPUT72), .B(KEYINPUT6), .Z(n561) );
  XNOR2_X1 U624 ( .A(n562), .B(n561), .ZN(n563) );
  NAND2_X1 U625 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U626 ( .A(KEYINPUT7), .B(n565), .ZN(G168) );
  XOR2_X1 U627 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U628 ( .A1(G88), .A2(n797), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G75), .A2(n798), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n793), .A2(G50), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G62), .A2(n794), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U635 ( .A(G166), .ZN(G303) );
  NAND2_X1 U636 ( .A1(G651), .A2(G74), .ZN(n572) );
  XOR2_X1 U637 ( .A(KEYINPUT76), .B(n572), .Z(n573) );
  NOR2_X1 U638 ( .A1(n794), .A2(n573), .ZN(n575) );
  NAND2_X1 U639 ( .A1(n793), .A2(G49), .ZN(n574) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(KEYINPUT77), .ZN(n579) );
  NAND2_X1 U642 ( .A1(G87), .A2(n577), .ZN(n578) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(G288) );
  NAND2_X1 U644 ( .A1(n797), .A2(G86), .ZN(n581) );
  NAND2_X1 U645 ( .A1(G61), .A2(n794), .ZN(n580) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n584) );
  NAND2_X1 U647 ( .A1(n798), .A2(G73), .ZN(n582) );
  XOR2_X1 U648 ( .A(KEYINPUT2), .B(n582), .Z(n583) );
  NOR2_X1 U649 ( .A1(n584), .A2(n583), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n793), .A2(G48), .ZN(n585) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(G305) );
  NAND2_X1 U652 ( .A1(n797), .A2(G85), .ZN(n588) );
  NAND2_X1 U653 ( .A1(G60), .A2(n794), .ZN(n587) );
  NAND2_X1 U654 ( .A1(n588), .A2(n587), .ZN(n591) );
  NAND2_X1 U655 ( .A1(G47), .A2(n793), .ZN(n589) );
  XNOR2_X1 U656 ( .A(KEYINPUT69), .B(n589), .ZN(n590) );
  NOR2_X1 U657 ( .A1(n591), .A2(n590), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n798), .A2(G72), .ZN(n592) );
  NAND2_X1 U659 ( .A1(n593), .A2(n592), .ZN(G290) );
  XOR2_X1 U660 ( .A(KEYINPUT92), .B(KEYINPUT28), .Z(n601) );
  AND2_X1 U661 ( .A1(G160), .A2(G40), .ZN(n594) );
  NAND2_X1 U662 ( .A1(n594), .A2(n709), .ZN(n596) );
  INV_X1 U663 ( .A(KEYINPUT64), .ZN(n595) );
  XNOR2_X2 U664 ( .A(n596), .B(n595), .ZN(n647) );
  NAND2_X1 U665 ( .A1(G2072), .A2(n647), .ZN(n597) );
  XOR2_X1 U666 ( .A(KEYINPUT27), .B(n597), .Z(n599) );
  XOR2_X1 U667 ( .A(G1956), .B(KEYINPUT91), .Z(n918) );
  NAND2_X1 U668 ( .A1(n664), .A2(n918), .ZN(n598) );
  NAND2_X1 U669 ( .A1(n599), .A2(n598), .ZN(n638) );
  NAND2_X1 U670 ( .A1(n638), .A2(G299), .ZN(n600) );
  XNOR2_X1 U671 ( .A(n601), .B(n600), .ZN(n643) );
  NAND2_X1 U672 ( .A1(n664), .A2(G1341), .ZN(n603) );
  INV_X1 U673 ( .A(KEYINPUT94), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n603), .B(n602), .ZN(n614) );
  NAND2_X1 U675 ( .A1(n794), .A2(G56), .ZN(n604) );
  XOR2_X1 U676 ( .A(KEYINPUT14), .B(n604), .Z(n611) );
  NAND2_X1 U677 ( .A1(G81), .A2(n797), .ZN(n605) );
  XNOR2_X1 U678 ( .A(n605), .B(KEYINPUT70), .ZN(n606) );
  XNOR2_X1 U679 ( .A(n606), .B(KEYINPUT12), .ZN(n608) );
  NAND2_X1 U680 ( .A1(G68), .A2(n798), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n608), .A2(n607), .ZN(n609) );
  XOR2_X1 U682 ( .A(KEYINPUT13), .B(n609), .Z(n610) );
  NOR2_X1 U683 ( .A1(n611), .A2(n610), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n793), .A2(G43), .ZN(n612) );
  NAND2_X1 U685 ( .A1(n613), .A2(n612), .ZN(n998) );
  NOR2_X1 U686 ( .A1(n614), .A2(n998), .ZN(n632) );
  NAND2_X1 U687 ( .A1(n793), .A2(G54), .ZN(n621) );
  NAND2_X1 U688 ( .A1(G92), .A2(n797), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G79), .A2(n798), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n619) );
  NAND2_X1 U691 ( .A1(n794), .A2(G66), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n617), .B(KEYINPUT71), .ZN(n618) );
  NOR2_X1 U693 ( .A1(n619), .A2(n618), .ZN(n620) );
  NAND2_X1 U694 ( .A1(n621), .A2(n620), .ZN(n622) );
  XOR2_X1 U695 ( .A(KEYINPUT26), .B(KEYINPUT93), .Z(n624) );
  NAND2_X1 U696 ( .A1(G1996), .A2(n647), .ZN(n623) );
  XNOR2_X1 U697 ( .A(n624), .B(n623), .ZN(n633) );
  AND2_X1 U698 ( .A1(n803), .A2(n633), .ZN(n625) );
  AND2_X1 U699 ( .A1(n632), .A2(n625), .ZN(n630) );
  NAND2_X1 U700 ( .A1(G2067), .A2(n647), .ZN(n627) );
  NAND2_X1 U701 ( .A1(n664), .A2(G1348), .ZN(n626) );
  NAND2_X1 U702 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U703 ( .A(n628), .B(KEYINPUT95), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U705 ( .A(n631), .B(KEYINPUT96), .ZN(n636) );
  INV_X1 U706 ( .A(n803), .ZN(n1004) );
  NAND2_X1 U707 ( .A1(n633), .A2(n632), .ZN(n634) );
  AND2_X1 U708 ( .A1(n1004), .A2(n634), .ZN(n635) );
  XOR2_X1 U709 ( .A(KEYINPUT97), .B(n637), .Z(n641) );
  NOR2_X1 U710 ( .A1(G299), .A2(n638), .ZN(n639) );
  XNOR2_X1 U711 ( .A(KEYINPUT98), .B(n639), .ZN(n640) );
  NOR2_X1 U712 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U713 ( .A(n646), .B(n645), .ZN(n651) );
  XOR2_X1 U714 ( .A(G1961), .B(KEYINPUT90), .Z(n929) );
  NOR2_X1 U715 ( .A1(n929), .A2(n647), .ZN(n649) );
  XNOR2_X1 U716 ( .A(G2078), .B(KEYINPUT25), .ZN(n955) );
  NOR2_X1 U717 ( .A1(n664), .A2(n955), .ZN(n648) );
  NOR2_X1 U718 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U719 ( .A1(n652), .A2(G171), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n662) );
  NOR2_X1 U721 ( .A1(G171), .A2(n652), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT100), .ZN(n658) );
  NAND2_X1 U723 ( .A1(n664), .A2(G8), .ZN(n702) );
  NOR2_X1 U724 ( .A1(G1966), .A2(n702), .ZN(n675) );
  NOR2_X1 U725 ( .A1(n664), .A2(G2084), .ZN(n673) );
  NOR2_X1 U726 ( .A1(n675), .A2(n673), .ZN(n654) );
  NAND2_X1 U727 ( .A1(G8), .A2(n654), .ZN(n655) );
  XNOR2_X1 U728 ( .A(KEYINPUT30), .B(n655), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n656), .A2(G168), .ZN(n657) );
  NOR2_X1 U730 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U731 ( .A(KEYINPUT31), .B(n659), .ZN(n660) );
  XNOR2_X1 U732 ( .A(n660), .B(KEYINPUT101), .ZN(n661) );
  NAND2_X1 U733 ( .A1(n672), .A2(G286), .ZN(n669) );
  NOR2_X1 U734 ( .A1(G1971), .A2(n702), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT103), .B(n663), .Z(n666) );
  NOR2_X1 U736 ( .A1(n664), .A2(G2090), .ZN(n665) );
  NOR2_X1 U737 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U738 ( .A1(n667), .A2(G303), .ZN(n668) );
  NAND2_X1 U739 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U740 ( .A1(n670), .A2(G8), .ZN(n671) );
  XNOR2_X1 U741 ( .A(KEYINPUT102), .B(n672), .ZN(n677) );
  AND2_X1 U742 ( .A1(G8), .A2(n673), .ZN(n674) );
  NOR2_X1 U743 ( .A1(n675), .A2(n674), .ZN(n676) );
  NAND2_X1 U744 ( .A1(n677), .A2(n676), .ZN(n694) );
  NAND2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n1015) );
  INV_X1 U746 ( .A(n702), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n1015), .A2(n678), .ZN(n682) );
  INV_X1 U748 ( .A(n682), .ZN(n679) );
  AND2_X1 U749 ( .A1(n694), .A2(n679), .ZN(n680) );
  AND2_X1 U750 ( .A1(n693), .A2(n680), .ZN(n686) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n681) );
  NOR2_X1 U753 ( .A1(n687), .A2(n681), .ZN(n1000) );
  OR2_X1 U754 ( .A1(n682), .A2(n1000), .ZN(n684) );
  INV_X1 U755 ( .A(KEYINPUT33), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U757 ( .A1(n686), .A2(n685), .ZN(n692) );
  NAND2_X1 U758 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U759 ( .A1(n688), .A2(n702), .ZN(n690) );
  XOR2_X1 U760 ( .A(G1981), .B(G305), .Z(n1001) );
  NOR2_X1 U761 ( .A1(n692), .A2(n691), .ZN(n707) );
  NAND2_X1 U762 ( .A1(n694), .A2(n693), .ZN(n698) );
  NOR2_X1 U763 ( .A1(G2090), .A2(G303), .ZN(n695) );
  NAND2_X1 U764 ( .A1(G8), .A2(n695), .ZN(n696) );
  XNOR2_X1 U765 ( .A(n696), .B(KEYINPUT104), .ZN(n697) );
  NAND2_X1 U766 ( .A1(n698), .A2(n697), .ZN(n699) );
  NAND2_X1 U767 ( .A1(n699), .A2(n702), .ZN(n705) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XNOR2_X1 U769 ( .A(n700), .B(KEYINPUT24), .ZN(n701) );
  XNOR2_X1 U770 ( .A(n701), .B(KEYINPUT89), .ZN(n703) );
  OR2_X1 U771 ( .A1(n703), .A2(n702), .ZN(n704) );
  NAND2_X1 U772 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U773 ( .A1(G160), .A2(G40), .ZN(n708) );
  NOR2_X1 U774 ( .A1(n709), .A2(n708), .ZN(n755) );
  NAND2_X1 U775 ( .A1(n897), .A2(G117), .ZN(n710) );
  XNOR2_X1 U776 ( .A(n710), .B(KEYINPUT86), .ZN(n712) );
  NAND2_X1 U777 ( .A1(G129), .A2(n895), .ZN(n711) );
  NAND2_X1 U778 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U779 ( .A(n713), .B(KEYINPUT87), .ZN(n717) );
  NAND2_X1 U780 ( .A1(G141), .A2(n715), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U782 ( .A1(n892), .A2(G105), .ZN(n718) );
  XOR2_X1 U783 ( .A(KEYINPUT38), .B(n718), .Z(n719) );
  OR2_X1 U784 ( .A1(n720), .A2(n719), .ZN(n878) );
  NAND2_X1 U785 ( .A1(G1996), .A2(n878), .ZN(n729) );
  XNOR2_X1 U786 ( .A(KEYINPUT85), .B(G1991), .ZN(n945) );
  NAND2_X1 U787 ( .A1(G107), .A2(n897), .ZN(n722) );
  NAND2_X1 U788 ( .A1(G119), .A2(n895), .ZN(n721) );
  NAND2_X1 U789 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U790 ( .A(KEYINPUT84), .B(n723), .ZN(n727) );
  NAND2_X1 U791 ( .A1(n892), .A2(G95), .ZN(n725) );
  NAND2_X1 U792 ( .A1(G131), .A2(n715), .ZN(n724) );
  NAND2_X1 U793 ( .A1(n725), .A2(n724), .ZN(n726) );
  NOR2_X1 U794 ( .A1(n727), .A2(n726), .ZN(n875) );
  OR2_X1 U795 ( .A1(n945), .A2(n875), .ZN(n728) );
  NAND2_X1 U796 ( .A1(n729), .A2(n728), .ZN(n977) );
  NAND2_X1 U797 ( .A1(n755), .A2(n977), .ZN(n747) );
  NAND2_X1 U798 ( .A1(n892), .A2(G104), .ZN(n731) );
  NAND2_X1 U799 ( .A1(G140), .A2(n715), .ZN(n730) );
  NAND2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U801 ( .A(KEYINPUT34), .B(n732), .ZN(n737) );
  NAND2_X1 U802 ( .A1(G116), .A2(n897), .ZN(n734) );
  NAND2_X1 U803 ( .A1(G128), .A2(n895), .ZN(n733) );
  NAND2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U805 ( .A(KEYINPUT35), .B(n735), .Z(n736) );
  NOR2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U807 ( .A(KEYINPUT36), .B(n738), .ZN(n874) );
  XNOR2_X1 U808 ( .A(G2067), .B(KEYINPUT37), .ZN(n744) );
  NOR2_X1 U809 ( .A1(n874), .A2(n744), .ZN(n991) );
  NAND2_X1 U810 ( .A1(n755), .A2(n991), .ZN(n751) );
  NAND2_X1 U811 ( .A1(n747), .A2(n751), .ZN(n739) );
  XNOR2_X1 U812 ( .A(KEYINPUT88), .B(n739), .ZN(n742) );
  XOR2_X1 U813 ( .A(KEYINPUT83), .B(G1986), .Z(n740) );
  XOR2_X1 U814 ( .A(G290), .B(n740), .Z(n999) );
  INV_X1 U815 ( .A(n999), .ZN(n741) );
  NAND2_X1 U816 ( .A1(n517), .A2(n743), .ZN(n759) );
  NAND2_X1 U817 ( .A1(n874), .A2(n744), .ZN(n974) );
  OR2_X1 U818 ( .A1(n878), .A2(G1996), .ZN(n983) );
  NOR2_X1 U819 ( .A1(G1986), .A2(G290), .ZN(n745) );
  XNOR2_X1 U820 ( .A(n745), .B(KEYINPUT105), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n875), .A2(n945), .ZN(n971) );
  NAND2_X1 U822 ( .A1(n746), .A2(n971), .ZN(n748) );
  NAND2_X1 U823 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U824 ( .A1(n983), .A2(n749), .ZN(n750) );
  XOR2_X1 U825 ( .A(KEYINPUT39), .B(n750), .Z(n752) );
  NAND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  NAND2_X1 U827 ( .A1(n974), .A2(n753), .ZN(n754) );
  XNOR2_X1 U828 ( .A(KEYINPUT106), .B(n754), .ZN(n756) );
  NAND2_X1 U829 ( .A1(n756), .A2(n755), .ZN(n757) );
  XOR2_X1 U830 ( .A(KEYINPUT107), .B(n757), .Z(n758) );
  NAND2_X1 U831 ( .A1(n759), .A2(n758), .ZN(n760) );
  XNOR2_X1 U832 ( .A(n760), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U833 ( .A(G2443), .B(G2446), .Z(n762) );
  XNOR2_X1 U834 ( .A(G2427), .B(G2451), .ZN(n761) );
  XNOR2_X1 U835 ( .A(n762), .B(n761), .ZN(n768) );
  XOR2_X1 U836 ( .A(G2430), .B(G2454), .Z(n764) );
  XNOR2_X1 U837 ( .A(G1341), .B(G1348), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n764), .B(n763), .ZN(n766) );
  XOR2_X1 U839 ( .A(G2435), .B(G2438), .Z(n765) );
  XNOR2_X1 U840 ( .A(n766), .B(n765), .ZN(n767) );
  XOR2_X1 U841 ( .A(n768), .B(n767), .Z(n769) );
  AND2_X1 U842 ( .A1(G14), .A2(n769), .ZN(G401) );
  INV_X1 U843 ( .A(G171), .ZN(G301) );
  AND2_X1 U844 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U845 ( .A1(n897), .A2(G111), .ZN(n771) );
  NAND2_X1 U846 ( .A1(G135), .A2(n715), .ZN(n770) );
  NAND2_X1 U847 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U848 ( .A1(n895), .A2(G123), .ZN(n772) );
  XOR2_X1 U849 ( .A(KEYINPUT18), .B(n772), .Z(n773) );
  NOR2_X1 U850 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U851 ( .A1(n892), .A2(G99), .ZN(n775) );
  NAND2_X1 U852 ( .A1(n776), .A2(n775), .ZN(n970) );
  XNOR2_X1 U853 ( .A(G2096), .B(n970), .ZN(n777) );
  OR2_X1 U854 ( .A1(G2100), .A2(n777), .ZN(G156) );
  INV_X1 U855 ( .A(G57), .ZN(G237) );
  NAND2_X1 U856 ( .A1(G7), .A2(G661), .ZN(n778) );
  XOR2_X1 U857 ( .A(n778), .B(KEYINPUT10), .Z(n833) );
  NAND2_X1 U858 ( .A1(n833), .A2(G567), .ZN(n779) );
  XOR2_X1 U859 ( .A(KEYINPUT11), .B(n779), .Z(G234) );
  INV_X1 U860 ( .A(G860), .ZN(n786) );
  OR2_X1 U861 ( .A1(n998), .A2(n786), .ZN(G153) );
  NAND2_X1 U862 ( .A1(G868), .A2(G301), .ZN(n781) );
  INV_X1 U863 ( .A(G868), .ZN(n782) );
  NAND2_X1 U864 ( .A1(n1004), .A2(n782), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(G284) );
  NOR2_X1 U866 ( .A1(G286), .A2(n782), .ZN(n784) );
  NOR2_X1 U867 ( .A1(G868), .A2(G299), .ZN(n783) );
  NOR2_X1 U868 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U869 ( .A(KEYINPUT73), .B(n785), .Z(G297) );
  NAND2_X1 U870 ( .A1(G559), .A2(n786), .ZN(n787) );
  XNOR2_X1 U871 ( .A(KEYINPUT74), .B(n787), .ZN(n788) );
  NAND2_X1 U872 ( .A1(n788), .A2(n803), .ZN(n789) );
  XNOR2_X1 U873 ( .A(KEYINPUT16), .B(n789), .ZN(G148) );
  NOR2_X1 U874 ( .A1(G868), .A2(n998), .ZN(n792) );
  NAND2_X1 U875 ( .A1(n803), .A2(G868), .ZN(n790) );
  NOR2_X1 U876 ( .A1(G559), .A2(n790), .ZN(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(G282) );
  NAND2_X1 U878 ( .A1(n793), .A2(G55), .ZN(n796) );
  NAND2_X1 U879 ( .A1(G67), .A2(n794), .ZN(n795) );
  NAND2_X1 U880 ( .A1(n796), .A2(n795), .ZN(n802) );
  NAND2_X1 U881 ( .A1(G93), .A2(n797), .ZN(n800) );
  NAND2_X1 U882 ( .A1(G80), .A2(n798), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U884 ( .A1(n802), .A2(n801), .ZN(n810) );
  NAND2_X1 U885 ( .A1(G559), .A2(n803), .ZN(n804) );
  XNOR2_X1 U886 ( .A(n804), .B(n998), .ZN(n814) );
  NOR2_X1 U887 ( .A1(G860), .A2(n814), .ZN(n805) );
  XOR2_X1 U888 ( .A(KEYINPUT75), .B(n805), .Z(n806) );
  XNOR2_X1 U889 ( .A(n810), .B(n806), .ZN(G145) );
  NOR2_X1 U890 ( .A1(G868), .A2(n810), .ZN(n807) );
  XOR2_X1 U891 ( .A(n807), .B(KEYINPUT78), .Z(n817) );
  XOR2_X1 U892 ( .A(G303), .B(KEYINPUT19), .Z(n813) );
  XOR2_X1 U893 ( .A(G305), .B(G288), .Z(n808) );
  XNOR2_X1 U894 ( .A(G290), .B(n808), .ZN(n809) );
  XNOR2_X1 U895 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U896 ( .A(n811), .B(G299), .ZN(n812) );
  XNOR2_X1 U897 ( .A(n813), .B(n812), .ZN(n839) );
  XNOR2_X1 U898 ( .A(n839), .B(n814), .ZN(n815) );
  NAND2_X1 U899 ( .A1(G868), .A2(n815), .ZN(n816) );
  NAND2_X1 U900 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U901 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XOR2_X1 U902 ( .A(KEYINPUT20), .B(n818), .Z(n819) );
  NAND2_X1 U903 ( .A1(G2090), .A2(n819), .ZN(n820) );
  XNOR2_X1 U904 ( .A(KEYINPUT21), .B(n820), .ZN(n821) );
  NAND2_X1 U905 ( .A1(n821), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U906 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U907 ( .A1(G120), .A2(G69), .ZN(n822) );
  NOR2_X1 U908 ( .A1(G237), .A2(n822), .ZN(n823) );
  XNOR2_X1 U909 ( .A(KEYINPUT80), .B(n823), .ZN(n824) );
  NAND2_X1 U910 ( .A1(n824), .A2(G108), .ZN(n837) );
  NAND2_X1 U911 ( .A1(n837), .A2(G567), .ZN(n830) );
  XOR2_X1 U912 ( .A(KEYINPUT79), .B(KEYINPUT22), .Z(n826) );
  NAND2_X1 U913 ( .A1(G132), .A2(G82), .ZN(n825) );
  XNOR2_X1 U914 ( .A(n826), .B(n825), .ZN(n827) );
  NOR2_X1 U915 ( .A1(n827), .A2(G218), .ZN(n828) );
  NAND2_X1 U916 ( .A1(G96), .A2(n828), .ZN(n838) );
  NAND2_X1 U917 ( .A1(n838), .A2(G2106), .ZN(n829) );
  NAND2_X1 U918 ( .A1(n830), .A2(n829), .ZN(n916) );
  NAND2_X1 U919 ( .A1(G483), .A2(G661), .ZN(n831) );
  NOR2_X1 U920 ( .A1(n916), .A2(n831), .ZN(n832) );
  XOR2_X1 U921 ( .A(KEYINPUT81), .B(n832), .Z(n836) );
  NAND2_X1 U922 ( .A1(n836), .A2(G36), .ZN(G176) );
  NAND2_X1 U923 ( .A1(G2106), .A2(n833), .ZN(G217) );
  INV_X1 U924 ( .A(n833), .ZN(G223) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n834) );
  NAND2_X1 U926 ( .A1(G661), .A2(n834), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n835) );
  NAND2_X1 U928 ( .A1(n836), .A2(n835), .ZN(G188) );
  INV_X1 U930 ( .A(G132), .ZN(G219) );
  INV_X1 U931 ( .A(G120), .ZN(G236) );
  INV_X1 U932 ( .A(G108), .ZN(G238) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G82), .ZN(G220) );
  INV_X1 U935 ( .A(G69), .ZN(G235) );
  NOR2_X1 U936 ( .A1(n838), .A2(n837), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(n1004), .B(n998), .Z(n840) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(n841), .B(KEYINPUT118), .Z(n843) );
  XOR2_X1 U941 ( .A(G301), .B(G286), .Z(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  NOR2_X1 U943 ( .A1(G37), .A2(n844), .ZN(G397) );
  XOR2_X1 U944 ( .A(G1991), .B(G1986), .Z(n846) );
  XNOR2_X1 U945 ( .A(G1996), .B(G1976), .ZN(n845) );
  XNOR2_X1 U946 ( .A(n846), .B(n845), .ZN(n856) );
  XOR2_X1 U947 ( .A(G2474), .B(KEYINPUT111), .Z(n848) );
  XNOR2_X1 U948 ( .A(G1956), .B(KEYINPUT41), .ZN(n847) );
  XNOR2_X1 U949 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U950 ( .A(G1981), .B(G1971), .Z(n850) );
  XNOR2_X1 U951 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U952 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U953 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U954 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U955 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U956 ( .A(n856), .B(n855), .Z(G229) );
  XOR2_X1 U957 ( .A(G2096), .B(KEYINPUT43), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2067), .B(KEYINPUT108), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U960 ( .A(n859), .B(G2678), .Z(n861) );
  XNOR2_X1 U961 ( .A(G2072), .B(G2090), .ZN(n860) );
  XNOR2_X1 U962 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U963 ( .A(KEYINPUT42), .B(G2100), .Z(n863) );
  XNOR2_X1 U964 ( .A(G2084), .B(G2078), .ZN(n862) );
  XNOR2_X1 U965 ( .A(n863), .B(n862), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(G227) );
  NAND2_X1 U967 ( .A1(G124), .A2(n895), .ZN(n866) );
  XNOR2_X1 U968 ( .A(n866), .B(KEYINPUT44), .ZN(n869) );
  NAND2_X1 U969 ( .A1(n715), .A2(G136), .ZN(n867) );
  XNOR2_X1 U970 ( .A(n867), .B(KEYINPUT112), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n873) );
  NAND2_X1 U972 ( .A1(G100), .A2(n892), .ZN(n871) );
  NAND2_X1 U973 ( .A1(G112), .A2(n897), .ZN(n870) );
  NAND2_X1 U974 ( .A1(n871), .A2(n870), .ZN(n872) );
  NOR2_X1 U975 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U976 ( .A(n874), .B(G162), .ZN(n877) );
  XNOR2_X1 U977 ( .A(G164), .B(n875), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n879) );
  XNOR2_X1 U979 ( .A(n879), .B(n878), .ZN(n891) );
  NAND2_X1 U980 ( .A1(G118), .A2(n897), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n880), .B(KEYINPUT114), .ZN(n889) );
  NAND2_X1 U982 ( .A1(n895), .A2(G130), .ZN(n881) );
  XNOR2_X1 U983 ( .A(KEYINPUT113), .B(n881), .ZN(n887) );
  NAND2_X1 U984 ( .A1(n892), .A2(G106), .ZN(n883) );
  NAND2_X1 U985 ( .A1(G142), .A2(n715), .ZN(n882) );
  NAND2_X1 U986 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U987 ( .A(KEYINPUT45), .B(n884), .ZN(n885) );
  XNOR2_X1 U988 ( .A(KEYINPUT115), .B(n885), .ZN(n886) );
  NOR2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n908) );
  XOR2_X1 U992 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n905) );
  NAND2_X1 U993 ( .A1(n892), .A2(G103), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G139), .A2(n715), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U996 ( .A1(n895), .A2(G127), .ZN(n896) );
  XNOR2_X1 U997 ( .A(n896), .B(KEYINPUT116), .ZN(n899) );
  NAND2_X1 U998 ( .A1(G115), .A2(n897), .ZN(n898) );
  NAND2_X1 U999 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n900), .Z(n901) );
  NOR2_X1 U1001 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1002 ( .A(KEYINPUT117), .B(n903), .Z(n978) );
  XNOR2_X1 U1003 ( .A(G160), .B(n978), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(n905), .B(n904), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n970), .B(n906), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n909), .ZN(G395) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n910) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n911), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n916), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT119), .B(n912), .ZN(n913) );
  NOR2_X1 U1013 ( .A1(G395), .A2(n913), .ZN(n914) );
  NAND2_X1 U1014 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n916), .ZN(G319) );
  XNOR2_X1 U1017 ( .A(KEYINPUT125), .B(G1966), .ZN(n917) );
  XNOR2_X1 U1018 ( .A(n917), .B(G21), .ZN(n941) );
  XNOR2_X1 U1019 ( .A(n918), .B(G20), .ZN(n922) );
  XNOR2_X1 U1020 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n919) );
  XNOR2_X1 U1021 ( .A(n919), .B(G4), .ZN(n920) );
  XNOR2_X1 U1022 ( .A(n920), .B(G1348), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n926) );
  XNOR2_X1 U1024 ( .A(G1341), .B(G19), .ZN(n924) );
  XNOR2_X1 U1025 ( .A(G6), .B(G1981), .ZN(n923) );
  NOR2_X1 U1026 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1028 ( .A(n927), .B(KEYINPUT124), .ZN(n928) );
  XOR2_X1 U1029 ( .A(KEYINPUT60), .B(n928), .Z(n931) );
  XNOR2_X1 U1030 ( .A(n929), .B(G5), .ZN(n930) );
  NAND2_X1 U1031 ( .A1(n931), .A2(n930), .ZN(n939) );
  XNOR2_X1 U1032 ( .A(G1976), .B(G23), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(G1986), .B(G24), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n936) );
  XOR2_X1 U1035 ( .A(G1971), .B(KEYINPUT126), .Z(n934) );
  XNOR2_X1 U1036 ( .A(G22), .B(n934), .ZN(n935) );
  NAND2_X1 U1037 ( .A1(n936), .A2(n935), .ZN(n937) );
  XNOR2_X1 U1038 ( .A(KEYINPUT58), .B(n937), .ZN(n938) );
  NOR2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(n942), .B(KEYINPUT61), .Z(n943) );
  XNOR2_X1 U1042 ( .A(KEYINPUT127), .B(n943), .ZN(n944) );
  NOR2_X1 U1043 ( .A1(G16), .A2(n944), .ZN(n969) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n960) );
  XOR2_X1 U1045 ( .A(KEYINPUT121), .B(n945), .Z(n946) );
  XNOR2_X1 U1046 ( .A(n946), .B(G25), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G2072), .B(G33), .ZN(n948) );
  XNOR2_X1 U1048 ( .A(G2067), .B(G26), .ZN(n947) );
  NOR2_X1 U1049 ( .A1(n948), .A2(n947), .ZN(n949) );
  NAND2_X1 U1050 ( .A1(G28), .A2(n949), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(G32), .B(G1996), .ZN(n950) );
  XNOR2_X1 U1052 ( .A(KEYINPUT122), .B(n950), .ZN(n951) );
  NOR2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1054 ( .A1(n954), .A2(n953), .ZN(n957) );
  XOR2_X1 U1055 ( .A(G27), .B(n955), .Z(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n958) );
  XNOR2_X1 U1057 ( .A(KEYINPUT53), .B(n958), .ZN(n959) );
  NOR2_X1 U1058 ( .A1(n960), .A2(n959), .ZN(n963) );
  XOR2_X1 U1059 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1060 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1061 ( .A1(n963), .A2(n962), .ZN(n964) );
  XOR2_X1 U1062 ( .A(KEYINPUT55), .B(n964), .Z(n966) );
  INV_X1 U1063 ( .A(G29), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n967), .ZN(n968) );
  NOR2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n997) );
  NAND2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n973) );
  XOR2_X1 U1068 ( .A(G160), .B(G2084), .Z(n972) );
  NOR2_X1 U1069 ( .A1(n973), .A2(n972), .ZN(n975) );
  NAND2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n989) );
  XNOR2_X1 U1072 ( .A(G164), .B(G2078), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G2072), .B(n978), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(n979), .B(KEYINPUT120), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(n982), .B(KEYINPUT50), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(G162), .B(G2090), .ZN(n984) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n985) );
  XOR2_X1 U1079 ( .A(KEYINPUT51), .B(n985), .Z(n986) );
  NOR2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n990) );
  NOR2_X1 U1082 ( .A1(n991), .A2(n990), .ZN(n992) );
  XNOR2_X1 U1083 ( .A(KEYINPUT52), .B(n992), .ZN(n994) );
  INV_X1 U1084 ( .A(KEYINPUT55), .ZN(n993) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n995), .A2(G29), .ZN(n996) );
  NAND2_X1 U1087 ( .A1(n997), .A2(n996), .ZN(n1022) );
  XOR2_X1 U1088 ( .A(KEYINPUT56), .B(G16), .Z(n1020) );
  XNOR2_X1 U1089 ( .A(G1341), .B(n998), .ZN(n1018) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1014) );
  XNOR2_X1 U1091 ( .A(G1966), .B(G168), .ZN(n1002) );
  NAND2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT57), .ZN(n1012) );
  XOR2_X1 U1094 ( .A(n1004), .B(G1348), .Z(n1006) );
  NAND2_X1 U1095 ( .A1(G1971), .A2(G303), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(G299), .B(G1956), .Z(n1008) );
  XOR2_X1 U1098 ( .A(G301), .B(G1961), .Z(n1007) );
  NAND2_X1 U1099 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1101 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NOR2_X1 U1102 ( .A1(n1014), .A2(n1013), .ZN(n1016) );
  NAND2_X1 U1103 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NOR2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XOR2_X1 U1107 ( .A(n1023), .B(KEYINPUT62), .Z(G150) );
  INV_X1 U1108 ( .A(G150), .ZN(G311) );
endmodule

