//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 0 1 0 0 1 1 0 1 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 1 1 0 1 0 0 0 1 1 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:32 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  INV_X1    g001(.A(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT11), .B(G169gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  AND2_X1   g006(.A1(G43gat), .A2(G50gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(G43gat), .A2(G50gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT15), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(G43gat), .ZN(new_n211));
  INV_X1    g010(.A(G50gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT15), .ZN(new_n214));
  NAND2_X1  g013(.A1(G43gat), .A2(G50gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n210), .A2(new_n216), .A3(KEYINPUT91), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT91), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n213), .A2(new_n218), .A3(new_n214), .A4(new_n215), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G29gat), .A2(G36gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT14), .B1(new_n221), .B2(KEYINPUT90), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT90), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n223), .A2(G29gat), .A3(G36gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT14), .ZN(new_n226));
  OAI211_X1 g025(.A(new_n223), .B(new_n226), .C1(G29gat), .C2(G36gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G29gat), .A2(G36gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n225), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT92), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n220), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n228), .B(new_n227), .C1(new_n222), .C2(new_n224), .ZN(new_n233));
  INV_X1    g032(.A(new_n210), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT92), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n233), .B1(new_n217), .B2(new_n219), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n239), .A2(KEYINPUT94), .ZN(new_n240));
  XNOR2_X1  g039(.A(G15gat), .B(G22gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G22gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G15gat), .ZN(new_n245));
  INV_X1    g044(.A(G15gat), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n246), .A2(G22gat), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT93), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n245), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(G1gat), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n241), .A2(new_n248), .A3(G1gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n243), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(KEYINPUT94), .A3(new_n239), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n239), .A2(KEYINPUT94), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n243), .A2(new_n251), .A3(new_n252), .A4(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n238), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n220), .A2(new_n230), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n231), .B1(new_n233), .B2(new_n234), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n261), .A2(new_n232), .A3(new_n256), .A4(new_n254), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n258), .A2(new_n262), .A3(KEYINPUT95), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  XOR2_X1   g063(.A(new_n264), .B(KEYINPUT13), .Z(new_n265));
  INV_X1    g064(.A(KEYINPUT95), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n238), .A2(new_n266), .A3(new_n257), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n263), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT96), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT96), .ZN(new_n270));
  NAND4_X1  g069(.A1(new_n263), .A2(new_n270), .A3(new_n265), .A4(new_n267), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g071(.A(KEYINPUT17), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n232), .B(new_n273), .C1(new_n236), .C2(new_n237), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n257), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n273), .B1(new_n261), .B2(new_n232), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n264), .B(new_n262), .C1(new_n275), .C2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT18), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n238), .A2(KEYINPUT17), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n257), .A3(new_n274), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT18), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n280), .A2(new_n281), .A3(new_n264), .A4(new_n262), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n278), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(new_n207), .B1(new_n272), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT97), .ZN(new_n286));
  AND4_X1   g085(.A1(new_n286), .A2(new_n272), .A3(new_n207), .A4(new_n283), .ZN(new_n287));
  AOI22_X1  g086(.A1(new_n269), .A2(new_n271), .B1(new_n278), .B2(new_n282), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n286), .B1(new_n288), .B2(new_n207), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n285), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G15gat), .B(G43gat), .Z(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(G169gat), .A2(G176gat), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT25), .B1(new_n302), .B2(KEYINPUT65), .ZN(new_n303));
  NAND2_X1  g102(.A1(G183gat), .A2(G190gat), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT24), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  OR2_X1    g105(.A1(new_n306), .A2(KEYINPUT64), .ZN(new_n307));
  NAND3_X1  g106(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n308), .B1(G183gat), .B2(G190gat), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n309), .B1(KEYINPUT64), .B2(new_n306), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n300), .A2(new_n301), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT65), .ZN(new_n312));
  AOI22_X1  g111(.A1(new_n307), .A2(new_n310), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(new_n301), .B(KEYINPUT66), .Z(new_n314));
  XNOR2_X1  g113(.A(KEYINPUT67), .B(G190gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n306), .A2(new_n308), .ZN(new_n317));
  OAI211_X1 g116(.A(new_n314), .B(new_n300), .C1(new_n316), .C2(new_n317), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n303), .A2(new_n313), .B1(KEYINPUT25), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(new_n315), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT27), .B(G183gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g121(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n323));
  OR2_X1    g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT26), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n301), .B1(new_n296), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n327));
  OR2_X1    g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n326), .A2(new_n327), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n296), .A2(new_n325), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n322), .A2(new_n323), .ZN(new_n332));
  NAND4_X1  g131(.A1(new_n324), .A2(new_n331), .A3(new_n332), .A4(new_n304), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n319), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT1), .ZN(new_n335));
  AND2_X1   g134(.A1(G127gat), .A2(G134gat), .ZN(new_n336));
  NOR2_X1   g135(.A1(G127gat), .A2(G134gat), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n335), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  XOR2_X1   g137(.A(KEYINPUT71), .B(G120gat), .Z(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(G113gat), .ZN(new_n340));
  INV_X1    g139(.A(G113gat), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(G120gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n338), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n340), .A2(KEYINPUT72), .A3(new_n342), .ZN(new_n346));
  XNOR2_X1  g145(.A(KEYINPUT70), .B(G134gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G127gat), .ZN(new_n348));
  INV_X1    g147(.A(G120gat), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(G113gat), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n342), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n337), .B1(new_n351), .B2(new_n335), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n345), .A2(new_n346), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n334), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n345), .A2(new_n346), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n348), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n357), .A2(new_n333), .A3(new_n319), .ZN(new_n358));
  INV_X1    g157(.A(G227gat), .ZN(new_n359));
  INV_X1    g158(.A(G233gat), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n358), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n295), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT34), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n354), .A2(new_n358), .ZN(new_n366));
  INV_X1    g165(.A(new_n361), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  AOI211_X1 g167(.A(KEYINPUT34), .B(new_n361), .C1(new_n354), .C2(new_n358), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n364), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n364), .A2(new_n368), .A3(new_n369), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n362), .A2(KEYINPUT32), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n373), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n368), .A2(new_n369), .ZN(new_n376));
  INV_X1    g175(.A(new_n364), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n375), .B1(new_n378), .B2(new_n370), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n374), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G197gat), .B(G204gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT22), .ZN(new_n383));
  INV_X1    g182(.A(G211gat), .ZN(new_n384));
  INV_X1    g183(.A(G218gat), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n382), .A2(new_n386), .ZN(new_n387));
  XNOR2_X1  g186(.A(G211gat), .B(G218gat), .ZN(new_n388));
  XNOR2_X1  g187(.A(new_n387), .B(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(KEYINPUT29), .B1(new_n319), .B2(new_n333), .ZN(new_n391));
  INV_X1    g190(.A(G226gat), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n392), .A2(new_n360), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI211_X1 g193(.A(new_n392), .B(new_n360), .C1(new_n319), .C2(new_n333), .ZN(new_n395));
  OAI21_X1  g194(.A(KEYINPUT73), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n395), .A2(KEYINPUT73), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n390), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n334), .A2(new_n393), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n399), .B1(new_n393), .B2(new_n391), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n400), .A2(new_n389), .ZN(new_n401));
  XNOR2_X1  g200(.A(G8gat), .B(G36gat), .ZN(new_n402));
  XNOR2_X1  g201(.A(G64gat), .B(G92gat), .ZN(new_n403));
  XOR2_X1   g202(.A(new_n402), .B(new_n403), .Z(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n398), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  OAI21_X1  g205(.A(KEYINPUT75), .B1(new_n406), .B2(KEYINPUT30), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n396), .A2(new_n397), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n389), .ZN(new_n409));
  INV_X1    g208(.A(new_n401), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n409), .A2(new_n410), .A3(new_n404), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT75), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT30), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n407), .A2(new_n414), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n409), .A2(KEYINPUT30), .A3(new_n410), .A4(new_n404), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT74), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n398), .A2(new_n401), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT74), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n418), .A2(new_n419), .A3(KEYINPUT30), .A4(new_n404), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n405), .B1(new_n398), .B2(new_n401), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n415), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT84), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n388), .A2(new_n382), .A3(KEYINPUT80), .A4(new_n386), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT29), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n425), .B(new_n426), .C1(new_n390), .C2(KEYINPUT80), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(G141gat), .B(G148gat), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT2), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n431), .B1(G155gat), .B2(G162gat), .ZN(new_n432));
  INV_X1    g231(.A(G155gat), .ZN(new_n433));
  INV_X1    g232(.A(G162gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n430), .A2(new_n432), .B1(KEYINPUT76), .B2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G155gat), .B(G162gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n436), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n429), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n426), .B1(new_n438), .B2(KEYINPUT3), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n389), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n439), .A2(new_n441), .B1(G228gat), .B2(G233gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(G228gat), .A2(G233gat), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n428), .B1(new_n389), .B2(KEYINPUT29), .ZN(new_n444));
  AOI21_X1  g243(.A(new_n443), .B1(new_n444), .B2(new_n438), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT81), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(new_n446), .A3(new_n389), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n446), .B1(new_n440), .B2(new_n389), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n445), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT82), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OAI211_X1 g251(.A(KEYINPUT82), .B(new_n445), .C1(new_n448), .C2(new_n449), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n442), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT83), .B1(new_n454), .B2(new_n244), .ZN(new_n455));
  XNOR2_X1  g254(.A(G78gat), .B(G106gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT79), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(KEYINPUT31), .ZN(new_n458));
  XNOR2_X1  g257(.A(new_n458), .B(new_n212), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n424), .B1(new_n455), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n452), .A2(new_n453), .ZN(new_n462));
  INV_X1    g261(.A(new_n442), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(G22gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n454), .A2(new_n244), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n455), .A2(new_n424), .A3(new_n459), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n461), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n469), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n467), .B1(new_n471), .B2(new_n460), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n381), .B(new_n423), .C1(new_n470), .C2(new_n472), .ZN(new_n473));
  XOR2_X1   g272(.A(new_n436), .B(new_n437), .Z(new_n474));
  NAND3_X1  g273(.A1(new_n355), .A2(new_n356), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT77), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT4), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n353), .A2(KEYINPUT77), .A3(new_n474), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(G225gat), .A2(G233gat), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n438), .B(new_n428), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n357), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n474), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n480), .A2(new_n481), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT5), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n357), .A2(new_n438), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n477), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(new_n481), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n486), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n486), .A3(new_n481), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n475), .A2(new_n478), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n494), .B1(new_n495), .B2(KEYINPUT4), .ZN(new_n496));
  AOI22_X1  g295(.A1(new_n485), .A2(new_n490), .B1(new_n492), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g296(.A(G1gat), .B(G29gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(new_n498), .B(KEYINPUT0), .ZN(new_n499));
  XNOR2_X1  g298(.A(G57gat), .B(G85gat), .ZN(new_n500));
  XOR2_X1   g299(.A(new_n499), .B(new_n500), .Z(new_n501));
  AOI21_X1  g300(.A(KEYINPUT6), .B1(new_n497), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n490), .A2(new_n485), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n492), .A2(new_n496), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g304(.A(new_n501), .B(KEYINPUT85), .Z(new_n506));
  NAND2_X1  g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n501), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n505), .A2(KEYINPUT6), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT35), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n473), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n472), .A2(new_n470), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n380), .ZN(new_n514));
  INV_X1    g313(.A(new_n423), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT78), .B1(new_n497), .B2(new_n501), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT78), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n505), .A2(new_n517), .A3(new_n509), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n502), .A3(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n519), .A2(new_n510), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n515), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT35), .B1(new_n514), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n512), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(KEYINPUT39), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n478), .B1(new_n477), .B2(new_n479), .ZN(new_n526));
  INV_X1    g325(.A(new_n483), .ZN(new_n527));
  NOR3_X1   g326(.A1(new_n526), .A2(new_n527), .A3(new_n494), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n528), .A2(KEYINPUT86), .A3(new_n481), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT86), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n531), .A2(new_n483), .A3(new_n493), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n532), .B2(new_n489), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n525), .B1(new_n529), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT86), .B1(new_n528), .B2(new_n481), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n532), .A2(new_n530), .A3(new_n489), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n488), .A2(new_n489), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n535), .A2(new_n536), .A3(KEYINPUT39), .A4(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT87), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT40), .ZN(new_n540));
  AOI21_X1  g339(.A(new_n506), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n534), .A2(new_n538), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  AND2_X1   g342(.A1(new_n543), .A2(new_n507), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n534), .A2(new_n538), .A3(new_n541), .ZN(new_n545));
  OAI21_X1  g344(.A(new_n545), .B1(new_n539), .B2(new_n540), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(new_n423), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT37), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n404), .A2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n395), .A2(KEYINPUT73), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n550), .B1(new_n400), .B2(KEYINPUT73), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n410), .B1(new_n551), .B2(new_n390), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n549), .B1(new_n552), .B2(new_n405), .ZN(new_n553));
  INV_X1    g352(.A(new_n400), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n548), .B1(new_n554), .B2(new_n389), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n555), .B1(new_n551), .B2(new_n389), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT38), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(KEYINPUT88), .B1(new_n553), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n549), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n422), .A2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT88), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n561), .A2(new_n562), .A3(new_n557), .A4(new_n556), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n508), .A2(new_n510), .A3(new_n411), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n418), .A2(new_n548), .ZN(new_n566));
  OAI211_X1 g365(.A(KEYINPUT89), .B(KEYINPUT38), .C1(new_n553), .C2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT89), .ZN(new_n568));
  AOI22_X1  g367(.A1(new_n422), .A2(new_n560), .B1(new_n552), .B2(KEYINPUT37), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n569), .B2(new_n557), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n565), .A3(new_n567), .A4(new_n570), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n547), .A2(new_n571), .A3(new_n513), .ZN(new_n572));
  OAI211_X1 g371(.A(new_n472), .B(new_n470), .C1(new_n423), .C2(new_n520), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT36), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(new_n374), .B2(new_n379), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n373), .B1(new_n371), .B2(new_n372), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n378), .A2(new_n375), .A3(new_n370), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n576), .A2(KEYINPUT36), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n572), .A2(new_n573), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n291), .B1(new_n524), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(G64gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  INV_X1    g383(.A(G71gat), .ZN(new_n585));
  INV_X1    g384(.A(G78gat), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT9), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n584), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n587), .A2(new_n584), .ZN(new_n590));
  OR2_X1    g389(.A1(G57gat), .A2(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G57gat), .A2(G64gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n591), .A2(KEYINPUT9), .A3(new_n592), .ZN(new_n593));
  AOI22_X1  g392(.A1(new_n583), .A2(new_n589), .B1(new_n590), .B2(new_n593), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n594), .A2(KEYINPUT21), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n597), .B(G127gat), .ZN(new_n598));
  OR2_X1    g397(.A1(new_n594), .A2(KEYINPUT99), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n594), .A2(KEYINPUT99), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(KEYINPUT21), .A3(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n257), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n598), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(G183gat), .B(G211gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT100), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(new_n433), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n605), .B(new_n607), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n603), .B(new_n608), .Z(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  AND3_X1   g409(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT101), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n612), .A2(KEYINPUT7), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT7), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(KEYINPUT101), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n613), .A2(new_n615), .A3(G85gat), .A4(G92gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(G85gat), .A2(G92gat), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n618), .A2(KEYINPUT101), .A3(new_n614), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT8), .ZN(new_n621));
  OR2_X1    g420(.A1(G85gat), .A2(G92gat), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(G99gat), .ZN(new_n624));
  INV_X1    g423(.A(G106gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT102), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n620), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n627), .B1(new_n626), .B2(new_n620), .ZN(new_n630));
  OAI22_X1  g429(.A1(new_n617), .A2(new_n623), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AND3_X1   g430(.A1(new_n619), .A2(new_n621), .A3(new_n622), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n620), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT102), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n632), .A2(new_n634), .A3(new_n628), .A4(new_n616), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n631), .A2(new_n635), .A3(KEYINPUT103), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT103), .B1(new_n631), .B2(new_n635), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n238), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n611), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT103), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n616), .A2(new_n621), .A3(new_n619), .A4(new_n622), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n634), .A2(new_n628), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AOI22_X1  g444(.A1(new_n632), .A2(new_n616), .B1(new_n634), .B2(new_n628), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n647), .A2(new_n636), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n279), .A2(new_n274), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n641), .A2(new_n649), .ZN(new_n650));
  XOR2_X1   g449(.A(G190gat), .B(G218gat), .Z(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n641), .A2(new_n649), .A3(new_n651), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT104), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n650), .A2(KEYINPUT104), .A3(new_n651), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n652), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n658), .B1(new_n656), .B2(new_n655), .ZN(new_n659));
  XNOR2_X1  g458(.A(G134gat), .B(G162gat), .ZN(new_n660));
  AOI21_X1  g459(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n657), .A2(new_n659), .A3(new_n663), .ZN(new_n664));
  AOI221_X4 g463(.A(new_n652), .B1(new_n658), .B2(new_n662), .C1(new_n655), .C2(new_n656), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT10), .ZN(new_n667));
  AND3_X1   g466(.A1(new_n631), .A2(new_n635), .A3(new_n594), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n594), .B1(new_n631), .B2(new_n635), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n667), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n594), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n673), .B1(new_n645), .B2(new_n646), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n631), .A2(new_n635), .A3(new_n594), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g475(.A(KEYINPUT106), .B1(new_n676), .B2(new_n667), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n599), .A2(KEYINPUT10), .A3(new_n600), .ZN(new_n678));
  OAI22_X1  g477(.A1(new_n672), .A2(new_n677), .B1(new_n648), .B2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(G230gat), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n680), .A2(new_n360), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n679), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g482(.A1(new_n674), .A2(new_n681), .A3(new_n675), .ZN(new_n684));
  XNOR2_X1  g483(.A(G120gat), .B(G148gat), .ZN(new_n685));
  XNOR2_X1  g484(.A(G176gat), .B(G204gat), .ZN(new_n686));
  XOR2_X1   g485(.A(new_n685), .B(new_n686), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n683), .A2(new_n684), .A3(new_n687), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n683), .B2(new_n684), .ZN(new_n690));
  NOR2_X1   g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g491(.A1(new_n610), .A2(new_n666), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n581), .A2(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n521), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n250), .ZN(G1324gat));
  INV_X1    g495(.A(KEYINPUT42), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n694), .A2(new_n515), .ZN(new_n698));
  XOR2_X1   g497(.A(KEYINPUT16), .B(G8gat), .Z(new_n699));
  AOI21_X1  g498(.A(new_n697), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G8gat), .B1(new_n694), .B2(new_n515), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT107), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n699), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n697), .A2(KEYINPUT107), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n699), .B2(new_n704), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n700), .A2(new_n701), .B1(new_n698), .B2(new_n705), .ZN(G1325gat));
  INV_X1    g505(.A(new_n694), .ZN(new_n707));
  AOI21_X1  g506(.A(G15gat), .B1(new_n707), .B2(new_n380), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709));
  AND3_X1   g508(.A1(new_n575), .A2(new_n578), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n709), .B1(new_n575), .B2(new_n578), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n246), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT109), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n708), .B1(new_n707), .B2(new_n714), .ZN(G1326gat));
  NOR2_X1   g514(.A1(new_n694), .A2(new_n513), .ZN(new_n716));
  XOR2_X1   g515(.A(KEYINPUT43), .B(G22gat), .Z(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  NAND2_X1  g517(.A1(new_n610), .A2(new_n691), .ZN(new_n719));
  INV_X1    g518(.A(new_n666), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n521), .A2(G29gat), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n581), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(KEYINPUT110), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(KEYINPUT45), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT44), .ZN(new_n728));
  AND3_X1   g527(.A1(new_n547), .A2(new_n571), .A3(new_n513), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n712), .A2(new_n573), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT112), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT112), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n572), .A2(new_n732), .A3(new_n573), .A4(new_n712), .ZN(new_n733));
  AOI22_X1  g532(.A1(new_n731), .A2(new_n733), .B1(new_n523), .B2(new_n512), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n728), .B1(new_n734), .B2(new_n720), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n524), .A2(new_n580), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n736), .A2(KEYINPUT44), .A3(new_n666), .ZN(new_n737));
  AND2_X1   g536(.A1(new_n735), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT111), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n272), .A2(new_n207), .A3(new_n283), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT97), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n288), .A2(new_n286), .A3(new_n207), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n739), .B1(new_n743), .B2(new_n285), .ZN(new_n744));
  AOI211_X1 g543(.A(KEYINPUT111), .B(new_n284), .C1(new_n741), .C2(new_n742), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n747), .A2(new_n719), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n738), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g548(.A(G29gat), .B1(new_n749), .B2(new_n521), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n724), .A2(KEYINPUT45), .A3(new_n725), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n727), .A2(new_n750), .A3(new_n751), .ZN(G1328gat));
  NAND4_X1  g551(.A1(new_n735), .A2(new_n423), .A3(new_n737), .A4(new_n748), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(G36gat), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n515), .A2(G36gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n581), .A2(new_n721), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n757));
  OR2_X1    g556(.A1(new_n756), .A2(KEYINPUT46), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(new_n757), .A3(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1329gat));
  INV_X1    g560(.A(new_n712), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n735), .A2(new_n762), .A3(new_n737), .A4(new_n748), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G43gat), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n581), .A2(new_n721), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n765), .A2(G43gat), .A3(new_n381), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT47), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n764), .A2(new_n769), .ZN(new_n770));
  OR2_X1    g569(.A1(new_n767), .A2(KEYINPUT114), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1330gat));
  OAI21_X1  g571(.A(new_n212), .B1(new_n765), .B2(new_n513), .ZN(new_n773));
  INV_X1    g572(.A(new_n513), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(G50gat), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n749), .B2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n776), .A2(KEYINPUT48), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n778), .B(new_n773), .C1(new_n749), .C2(new_n775), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1331gat));
  NAND4_X1  g579(.A1(new_n747), .A2(new_n720), .A3(new_n609), .A4(new_n692), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n734), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(new_n520), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n783), .B(G57gat), .ZN(G1332gat));
  INV_X1    g583(.A(KEYINPUT49), .ZN(new_n785));
  INV_X1    g584(.A(G64gat), .ZN(new_n786));
  OAI211_X1 g585(.A(new_n782), .B(new_n423), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(KEYINPUT115), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n787), .A2(KEYINPUT115), .ZN(new_n790));
  OAI22_X1  g589(.A1(new_n789), .A2(new_n790), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n787), .A2(KEYINPUT115), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n792), .A2(new_n785), .A3(new_n786), .A4(new_n788), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(G1333gat));
  NAND3_X1  g593(.A1(new_n782), .A2(new_n585), .A3(new_n380), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n734), .A2(new_n712), .A3(new_n781), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n796), .B2(new_n585), .ZN(new_n797));
  XOR2_X1   g596(.A(new_n797), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n774), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g599(.A1(new_n746), .A2(new_n609), .ZN(new_n801));
  INV_X1    g600(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n691), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n738), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n520), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(G85gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n731), .A2(new_n733), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n720), .B1(new_n807), .B2(new_n524), .ZN(new_n808));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n808), .B2(new_n801), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT51), .ZN(new_n810));
  NOR4_X1   g609(.A1(new_n734), .A2(new_n810), .A3(new_n720), .A4(new_n802), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n521), .A2(G85gat), .A3(new_n691), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n806), .A2(new_n814), .ZN(G1336gat));
  NAND4_X1  g614(.A1(new_n735), .A2(new_n423), .A3(new_n737), .A4(new_n803), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G92gat), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n515), .A2(G92gat), .A3(new_n691), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n818), .B1(new_n809), .B2(new_n811), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g619(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n820), .B(new_n821), .ZN(G1337gat));
  NAND4_X1  g621(.A1(new_n812), .A2(new_n624), .A3(new_n380), .A4(new_n692), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n804), .A2(new_n762), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n624), .ZN(G1338gat));
  NOR2_X1   g624(.A1(new_n513), .A2(new_n691), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n826), .B1(new_n809), .B2(new_n811), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n625), .ZN(new_n828));
  NAND2_X1  g627(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n513), .A2(new_n625), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n735), .A2(new_n737), .A3(new_n803), .A4(new_n830), .ZN(new_n831));
  OR2_X1    g630(.A1(KEYINPUT117), .A2(KEYINPUT53), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND3_X1   g632(.A1(new_n828), .A2(new_n829), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n829), .B1(new_n828), .B2(new_n833), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n834), .A2(new_n835), .ZN(G1339gat));
  NAND2_X1  g635(.A1(new_n747), .A2(new_n693), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT54), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n679), .A2(new_n839), .A3(new_n682), .ZN(new_n840));
  INV_X1    g639(.A(new_n687), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n648), .A2(new_n678), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n670), .A2(new_n671), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n676), .A2(KEYINPUT106), .A3(new_n667), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(KEYINPUT54), .B1(new_n845), .B2(new_n681), .ZN(new_n846));
  AOI211_X1 g645(.A(new_n682), .B(new_n842), .C1(new_n843), .C2(new_n844), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n840), .B(new_n841), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT55), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n688), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n845), .A2(new_n681), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n687), .B1(new_n851), .B2(new_n839), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n845), .A2(new_n681), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n683), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT55), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n265), .B1(new_n263), .B2(new_n267), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n264), .B1(new_n280), .B2(new_n262), .ZN(new_n858));
  OR2_X1    g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g658(.A1(new_n741), .A2(new_n742), .B1(new_n206), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n666), .A2(new_n856), .A3(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n692), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n863), .B1(new_n746), .B2(new_n856), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n861), .B1(new_n864), .B2(new_n666), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n838), .B1(new_n865), .B2(new_n610), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n521), .ZN(new_n867));
  AND2_X1   g666(.A1(new_n867), .A2(new_n473), .ZN(new_n868));
  AOI21_X1  g667(.A(G113gat), .B1(new_n868), .B2(new_n746), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n290), .A2(KEYINPUT111), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n743), .A2(new_n739), .A3(new_n285), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(new_n871), .A3(new_n856), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n666), .B1(new_n872), .B2(new_n862), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n666), .A2(new_n856), .A3(new_n860), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n610), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(new_n837), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n513), .ZN(new_n877));
  XNOR2_X1  g676(.A(new_n877), .B(KEYINPUT118), .ZN(new_n878));
  AND4_X1   g677(.A1(new_n520), .A2(new_n878), .A3(new_n515), .A4(new_n380), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n291), .A2(new_n341), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(G1340gat));
  NAND3_X1  g680(.A1(new_n868), .A2(new_n339), .A3(new_n692), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n879), .A2(new_n692), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n882), .B1(new_n884), .B2(new_n349), .ZN(G1341gat));
  INV_X1    g684(.A(G127gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n868), .A2(new_n886), .A3(new_n609), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n879), .A2(new_n609), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n886), .ZN(G1342gat));
  NAND2_X1  g689(.A1(new_n879), .A2(new_n666), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(G134gat), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n347), .B1(KEYINPUT119), .B2(KEYINPUT56), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n666), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g693(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n894), .B(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n892), .A2(new_n896), .ZN(G1343gat));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  OAI211_X1 g697(.A(KEYINPUT120), .B(new_n898), .C1(new_n866), .C2(new_n513), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n513), .B1(new_n875), .B2(new_n837), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n900), .B1(new_n901), .B2(KEYINPUT57), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n290), .A2(new_n856), .B1(new_n860), .B2(new_n692), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n861), .B1(new_n903), .B2(new_n666), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n837), .B1(new_n905), .B2(new_n609), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n906), .A2(KEYINPUT57), .A3(new_n774), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n899), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n762), .A2(new_n521), .A3(new_n423), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G141gat), .B1(new_n910), .B2(new_n291), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n762), .A2(new_n513), .ZN(new_n912));
  INV_X1    g711(.A(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(new_n423), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n867), .A2(new_n914), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(G141gat), .A3(new_n291), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n916), .A2(KEYINPUT58), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(new_n910), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n746), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n916), .B1(new_n920), .B2(G141gat), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT58), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n921), .B2(new_n922), .ZN(G1344gat));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n692), .A3(new_n909), .ZN(new_n924));
  INV_X1    g723(.A(G148gat), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n925), .A2(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n924), .A2(new_n926), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT122), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n774), .A2(new_n898), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n856), .A2(new_n290), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n666), .B1(new_n930), .B2(new_n862), .ZN(new_n931));
  OAI21_X1  g730(.A(KEYINPUT121), .B1(new_n931), .B2(new_n874), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT121), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n861), .B(new_n933), .C1(new_n903), .C2(new_n666), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(new_n610), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n693), .A2(new_n291), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n876), .A2(new_n774), .ZN(new_n938));
  AOI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(KEYINPUT57), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n909), .A2(new_n692), .ZN(new_n940));
  INV_X1    g739(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n925), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(KEYINPUT59), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n928), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n609), .B1(new_n904), .B2(KEYINPUT121), .ZN(new_n945));
  AOI22_X1  g744(.A1(new_n945), .A2(new_n934), .B1(new_n291), .B2(new_n693), .ZN(new_n946));
  OAI22_X1  g745(.A1(new_n901), .A2(new_n898), .B1(new_n946), .B2(new_n929), .ZN(new_n947));
  OAI21_X1  g746(.A(G148gat), .B1(new_n947), .B2(new_n940), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n948), .A2(KEYINPUT122), .A3(KEYINPUT59), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n927), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n915), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n925), .A3(new_n692), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT123), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n950), .A2(new_n955), .A3(new_n952), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n954), .A2(new_n956), .ZN(G1345gat));
  OAI21_X1  g756(.A(G155gat), .B1(new_n910), .B2(new_n610), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n951), .A2(new_n433), .A3(new_n609), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(G1346gat));
  AOI21_X1  g759(.A(G162gat), .B1(new_n951), .B2(new_n666), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n720), .A2(new_n434), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n919), .B2(new_n962), .ZN(G1347gat));
  NAND2_X1  g762(.A1(new_n876), .A2(new_n521), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT124), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n514), .A2(new_n515), .ZN(new_n966));
  AND2_X1   g765(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n746), .ZN(new_n968));
  NOR3_X1   g767(.A1(new_n515), .A2(new_n520), .A3(new_n381), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n878), .A2(new_n969), .ZN(new_n970));
  INV_X1    g769(.A(new_n970), .ZN(new_n971));
  AND2_X1   g770(.A1(new_n290), .A2(G169gat), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(G1348gat));
  NAND3_X1  g772(.A1(new_n971), .A2(G176gat), .A3(new_n692), .ZN(new_n974));
  INV_X1    g773(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g774(.A(G176gat), .B1(new_n967), .B2(new_n692), .ZN(new_n976));
  OR2_X1    g775(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(KEYINPUT125), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n975), .B1(new_n977), .B2(new_n978), .ZN(G1349gat));
  OAI21_X1  g778(.A(G183gat), .B1(new_n970), .B2(new_n610), .ZN(new_n980));
  INV_X1    g779(.A(new_n967), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n609), .A2(new_n321), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n980), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(KEYINPUT60), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT60), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n980), .B(new_n985), .C1(new_n981), .C2(new_n982), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n984), .A2(new_n986), .ZN(G1350gat));
  NAND3_X1  g786(.A1(new_n967), .A2(new_n320), .A3(new_n666), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n971), .A2(new_n666), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n989), .A2(new_n990), .A3(G190gat), .ZN(new_n991));
  AOI21_X1  g790(.A(new_n990), .B1(new_n989), .B2(G190gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1351gat));
  NOR2_X1   g792(.A1(new_n515), .A2(new_n520), .ZN(new_n994));
  NAND3_X1  g793(.A1(new_n939), .A2(new_n712), .A3(new_n994), .ZN(new_n995));
  NOR3_X1   g794(.A1(new_n995), .A2(new_n203), .A3(new_n291), .ZN(new_n996));
  NOR2_X1   g795(.A1(new_n913), .A2(new_n515), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n965), .A2(new_n997), .ZN(new_n998));
  OR2_X1    g797(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n1000));
  NAND3_X1  g799(.A1(new_n999), .A2(new_n746), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g800(.A(new_n996), .B1(new_n1001), .B2(new_n203), .ZN(G1352gat));
  OR3_X1    g801(.A1(new_n998), .A2(G204gat), .A3(new_n691), .ZN(new_n1003));
  OR2_X1    g802(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1004));
  OAI21_X1  g803(.A(G204gat), .B1(new_n995), .B2(new_n691), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1003), .A2(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .ZN(G1353gat));
  OAI21_X1  g806(.A(G211gat), .B1(new_n995), .B2(new_n610), .ZN(new_n1008));
  XOR2_X1   g807(.A(new_n1008), .B(KEYINPUT63), .Z(new_n1009));
  NAND2_X1  g808(.A1(new_n999), .A2(new_n1000), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n609), .A2(new_n384), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1009), .B1(new_n1010), .B2(new_n1011), .ZN(G1354gat));
  OAI21_X1  g811(.A(G218gat), .B1(new_n995), .B2(new_n720), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n666), .A2(new_n385), .ZN(new_n1014));
  OAI21_X1  g813(.A(new_n1013), .B1(new_n1010), .B2(new_n1014), .ZN(G1355gat));
endmodule


