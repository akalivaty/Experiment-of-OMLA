//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 0 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n831,
    new_n832, new_n833, new_n834, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n886, new_n887, new_n888, new_n889, new_n891, new_n892,
    new_n893, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n950, new_n951, new_n952, new_n954,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  INV_X1    g001(.A(G36gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  INV_X1    g005(.A(G43gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n207), .A2(G50gat), .ZN(new_n208));
  AND3_X1   g007(.A1(new_n206), .A2(new_n208), .A3(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT14), .ZN(new_n210));
  NAND3_X1  g009(.A1(new_n210), .A2(new_n202), .A3(new_n203), .ZN(new_n211));
  OAI21_X1  g010(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  AOI211_X1 g011(.A(new_n204), .B(new_n209), .C1(new_n211), .C2(new_n212), .ZN(new_n213));
  XNOR2_X1  g012(.A(new_n208), .B(KEYINPUT92), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n206), .B(KEYINPUT91), .ZN(new_n215));
  AND2_X1   g014(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n213), .B1(KEYINPUT15), .B2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n212), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT90), .ZN(new_n219));
  MUX2_X1   g018(.A(KEYINPUT90), .B(new_n219), .S(new_n211), .Z(new_n220));
  OAI21_X1  g019(.A(new_n209), .B1(new_n220), .B2(new_n204), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT93), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT93), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n222), .A2(new_n226), .A3(new_n223), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g027(.A(G15gat), .B(G22gat), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n229), .A2(KEYINPUT94), .ZN(new_n230));
  NOR2_X1   g029(.A1(new_n229), .A2(KEYINPUT94), .ZN(new_n231));
  OR3_X1    g030(.A1(new_n230), .A2(new_n231), .A3(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT96), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT16), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT95), .B(G1gat), .ZN(new_n235));
  OAI22_X1  g034(.A1(new_n230), .A2(new_n231), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n233), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(G8gat), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n232), .A2(new_n233), .A3(new_n239), .A4(new_n236), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT97), .ZN(new_n242));
  NOR2_X1   g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n217), .A2(KEYINPUT17), .A3(new_n221), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n242), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n228), .A2(new_n244), .A3(new_n245), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G229gat), .A2(G233gat), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n248), .B(KEYINPUT98), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n241), .A2(new_n222), .ZN(new_n251));
  NAND3_X1  g050(.A1(new_n247), .A2(new_n250), .A3(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n247), .A2(KEYINPUT18), .A3(new_n250), .A4(new_n251), .ZN(new_n255));
  XNOR2_X1  g054(.A(new_n241), .B(new_n222), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n249), .B(KEYINPUT13), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  XNOR2_X1  g057(.A(G113gat), .B(G141gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT11), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n260), .B(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT89), .B(G197gat), .ZN(new_n263));
  XNOR2_X1  g062(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT12), .ZN(new_n265));
  NAND4_X1  g064(.A1(new_n254), .A2(new_n255), .A3(new_n258), .A4(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT99), .ZN(new_n267));
  INV_X1    g066(.A(new_n265), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n246), .A2(new_n245), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n269), .A2(new_n243), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n270), .A2(new_n228), .B1(new_n222), .B2(new_n241), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT18), .B1(new_n271), .B2(new_n250), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n258), .ZN(new_n273));
  OAI211_X1 g072(.A(new_n267), .B(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n254), .A2(new_n255), .A3(new_n258), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n267), .B1(new_n276), .B2(new_n268), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n266), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  XNOR2_X1  g078(.A(G211gat), .B(G218gat), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G197gat), .B(G204gat), .ZN(new_n282));
  INV_X1    g081(.A(G218gat), .ZN(new_n283));
  INV_X1    g082(.A(G211gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(G211gat), .ZN(new_n287));
  AOI21_X1  g086(.A(new_n283), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  OAI211_X1 g087(.A(KEYINPUT74), .B(new_n282), .C1(new_n288), .C2(KEYINPUT22), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT22), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT73), .B(G211gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(new_n283), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT74), .B1(new_n293), .B2(new_n282), .ZN(new_n294));
  OAI211_X1 g093(.A(KEYINPUT75), .B(new_n281), .C1(new_n290), .C2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n282), .B1(new_n288), .B2(KEYINPUT22), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  AOI21_X1  g097(.A(new_n280), .B1(new_n298), .B2(new_n289), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT75), .ZN(new_n300));
  XOR2_X1   g099(.A(G197gat), .B(G204gat), .Z(new_n301));
  NOR2_X1   g100(.A1(new_n286), .A2(G211gat), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n284), .A2(KEYINPUT73), .ZN(new_n303));
  OAI21_X1  g102(.A(G218gat), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n301), .B1(new_n304), .B2(new_n291), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n300), .B1(new_n305), .B2(new_n280), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n295), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT29), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT3), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G148gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT79), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT79), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G148gat), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(new_n313), .A3(G141gat), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(G148gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NOR2_X1   g116(.A1(G155gat), .A2(G162gat), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT2), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n320), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n310), .A2(G141gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n316), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n325), .A2(new_n319), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n321), .A2(new_n318), .ZN(new_n327));
  AOI22_X1  g126(.A1(new_n317), .A2(new_n323), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT83), .B1(new_n309), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT84), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT83), .ZN(new_n331));
  XNOR2_X1  g130(.A(G141gat), .B(G148gat), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n327), .B1(new_n332), .B2(KEYINPUT2), .ZN(new_n333));
  INV_X1    g132(.A(new_n316), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT79), .B(G148gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n335), .B2(G141gat), .ZN(new_n336));
  AOI21_X1  g135(.A(new_n321), .B1(new_n319), .B2(new_n318), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n333), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n281), .B1(new_n290), .B2(new_n294), .ZN(new_n339));
  INV_X1    g138(.A(new_n306), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT29), .B1(new_n341), .B2(new_n295), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n331), .B(new_n338), .C1(new_n342), .C2(KEYINPUT3), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT3), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(new_n333), .C1(new_n336), .C2(new_n337), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(new_n308), .ZN(new_n346));
  INV_X1    g145(.A(new_n346), .ZN(new_n347));
  OAI211_X1 g146(.A(G228gat), .B(G233gat), .C1(new_n307), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n329), .A2(new_n330), .A3(new_n343), .A4(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n305), .A2(new_n280), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n296), .A2(new_n281), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n338), .B1(new_n353), .B2(KEYINPUT3), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n354), .B1(new_n307), .B2(new_n347), .ZN(new_n355));
  INV_X1    g154(.A(G228gat), .ZN(new_n356));
  INV_X1    g155(.A(G233gat), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n355), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n350), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n298), .A2(new_n289), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n306), .B1(new_n360), .B2(new_n281), .ZN(new_n361));
  AOI211_X1 g160(.A(new_n300), .B(new_n280), .C1(new_n298), .C2(new_n289), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n308), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n328), .B1(new_n363), .B2(new_n344), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n348), .B1(new_n364), .B2(new_n331), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n330), .B1(new_n365), .B2(new_n329), .ZN(new_n366));
  OAI21_X1  g165(.A(G22gat), .B1(new_n359), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT85), .ZN(new_n368));
  INV_X1    g167(.A(new_n329), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n343), .A2(new_n349), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT84), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(G22gat), .ZN(new_n372));
  NAND4_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n350), .A4(new_n358), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n367), .A2(new_n373), .ZN(new_n374));
  XNOR2_X1  g173(.A(G78gat), .B(G106gat), .ZN(new_n375));
  XNOR2_X1  g174(.A(KEYINPUT31), .B(G50gat), .ZN(new_n376));
  XNOR2_X1  g175(.A(new_n375), .B(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n368), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  OAI211_X1 g178(.A(new_n367), .B(new_n373), .C1(KEYINPUT85), .C2(new_n377), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G1gat), .B(G29gat), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n382), .B(KEYINPUT0), .ZN(new_n383));
  XNOR2_X1  g182(.A(G57gat), .B(G85gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  AOI22_X1  g185(.A1(new_n314), .A2(new_n316), .B1(new_n322), .B2(new_n320), .ZN(new_n387));
  XNOR2_X1  g186(.A(G155gat), .B(G162gat), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n388), .B1(new_n319), .B2(new_n325), .ZN(new_n389));
  OAI21_X1  g188(.A(KEYINPUT3), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G127gat), .B(G134gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n392));
  INV_X1    g191(.A(G113gat), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n393), .A2(G120gat), .ZN(new_n394));
  INV_X1    g193(.A(G120gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n395), .A2(G113gat), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n391), .B(new_n392), .C1(new_n394), .C2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G113gat), .B(G120gat), .ZN(new_n398));
  INV_X1    g197(.A(G127gat), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n399), .A2(G134gat), .ZN(new_n400));
  NOR2_X1   g199(.A1(new_n399), .A2(G134gat), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n398), .A2(KEYINPUT1), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n397), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n390), .A2(new_n345), .A3(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n397), .A2(new_n402), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(new_n328), .A3(KEYINPUT4), .ZN(new_n406));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n407));
  OAI21_X1  g206(.A(new_n407), .B1(new_n338), .B2(new_n403), .ZN(new_n408));
  NAND2_X1  g207(.A1(G225gat), .A2(G233gat), .ZN(new_n409));
  NAND4_X1  g208(.A1(new_n404), .A2(new_n406), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n386), .B1(new_n410), .B2(KEYINPUT5), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n338), .A2(new_n403), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n317), .A2(new_n323), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n413), .A2(new_n333), .A3(new_n402), .A4(new_n397), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n409), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT5), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n409), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n338), .A2(new_n403), .ZN(new_n419));
  AOI22_X1  g218(.A1(new_n413), .A2(new_n333), .B1(new_n402), .B2(new_n397), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n416), .B(new_n418), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n411), .B1(new_n423), .B2(new_n410), .ZN(new_n424));
  AND4_X1   g223(.A1(new_n409), .A2(new_n404), .A3(new_n408), .A4(new_n406), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT5), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT81), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n419), .B2(new_n420), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(KEYINPUT80), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n429), .A2(KEYINPUT5), .A3(new_n410), .A4(new_n421), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n427), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n385), .B1(new_n424), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n423), .A2(new_n410), .A3(new_n411), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n430), .ZN(new_n435));
  INV_X1    g234(.A(new_n385), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n432), .A2(new_n433), .A3(new_n437), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT6), .A4(new_n436), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT88), .ZN(new_n441));
  INV_X1    g240(.A(G226gat), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n442), .A2(new_n357), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT23), .ZN(new_n445));
  OAI211_X1 g244(.A(new_n445), .B(KEYINPUT65), .C1(G169gat), .C2(G176gat), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n447), .A2(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(G183gat), .A2(G190gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT24), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT24), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(G183gat), .A3(G190gat), .ZN(new_n452));
  AND2_X1   g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NOR2_X1   g252(.A1(G183gat), .A2(G190gat), .ZN(new_n454));
  OAI211_X1 g253(.A(new_n446), .B(new_n448), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  XOR2_X1   g254(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n456));
  AND2_X1   g255(.A1(new_n448), .A2(new_n446), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT25), .ZN(new_n458));
  INV_X1    g257(.A(G190gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT66), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT66), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G190gat), .ZN(new_n462));
  INV_X1    g261(.A(G183gat), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n460), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n450), .A2(new_n452), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n458), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n455), .A2(new_n456), .B1(new_n457), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT69), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n460), .A2(new_n462), .A3(KEYINPUT28), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT27), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(G183gat), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n463), .A2(KEYINPUT27), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  XNOR2_X1  g273(.A(KEYINPUT66), .B(G190gat), .ZN(new_n475));
  OAI21_X1  g274(.A(KEYINPUT67), .B1(new_n463), .B2(KEYINPUT27), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT27), .B(G183gat), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n475), .B(new_n476), .C1(new_n477), .C2(KEYINPUT67), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT28), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n474), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT26), .ZN(new_n481));
  INV_X1    g280(.A(G176gat), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n481), .A2(new_n261), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G169gat), .A2(G176gat), .ZN(new_n484));
  OAI211_X1 g283(.A(KEYINPUT68), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT68), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n449), .B1(new_n486), .B2(new_n490), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n468), .B1(new_n480), .B2(new_n491), .ZN(new_n492));
  AND3_X1   g291(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n493));
  AOI22_X1  g292(.A1(new_n493), .A2(new_n489), .B1(G183gat), .B2(G190gat), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n476), .A2(new_n460), .A3(new_n462), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT67), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n473), .A2(new_n496), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT28), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n494), .B(KEYINPUT69), .C1(new_n498), .C2(new_n474), .ZN(new_n499));
  AOI211_X1 g298(.A(new_n444), .B(new_n467), .C1(new_n492), .C2(new_n499), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n443), .A2(KEYINPUT29), .ZN(new_n501));
  INV_X1    g300(.A(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n467), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n494), .B1(new_n498), .B2(new_n474), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n502), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n307), .B1(new_n500), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g305(.A1(new_n361), .A2(new_n362), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n503), .A2(new_n504), .A3(new_n443), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n467), .B1(new_n492), .B2(new_n499), .ZN(new_n509));
  OAI211_X1 g308(.A(new_n507), .B(new_n508), .C1(new_n509), .C2(new_n502), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G8gat), .B(G36gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(G64gat), .B(G92gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT76), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(new_n514), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n506), .A2(new_n510), .A3(KEYINPUT30), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n506), .A2(new_n510), .A3(new_n517), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT30), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT78), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n520), .A2(KEYINPUT78), .A3(new_n521), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n519), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  AND3_X1   g325(.A1(new_n440), .A2(new_n441), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n441), .B1(new_n440), .B2(new_n526), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT34), .ZN(new_n530));
  NAND2_X1  g329(.A1(G227gat), .A2(G233gat), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT71), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n492), .A2(new_n499), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(new_n503), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n536), .A2(new_n405), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n509), .A2(new_n403), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n534), .B1(new_n539), .B2(new_n531), .ZN(new_n540));
  INV_X1    g339(.A(new_n531), .ZN(new_n541));
  AOI211_X1 g340(.A(new_n541), .B(new_n533), .C1(new_n537), .C2(new_n538), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(new_n541), .A3(new_n538), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT32), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT33), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(G15gat), .B(G43gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n548), .B(KEYINPUT70), .ZN(new_n549));
  XOR2_X1   g348(.A(G71gat), .B(G99gat), .Z(new_n550));
  XOR2_X1   g349(.A(new_n549), .B(new_n550), .Z(new_n551));
  NAND3_X1  g350(.A1(new_n545), .A2(new_n547), .A3(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n544), .B(KEYINPUT32), .C1(new_n546), .C2(new_n553), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n543), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n542), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n531), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n533), .ZN(new_n558));
  AOI22_X1  g357(.A1(new_n552), .A2(new_n554), .B1(new_n556), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n381), .A2(new_n529), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT35), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n552), .A2(new_n554), .ZN(new_n563));
  INV_X1    g362(.A(new_n543), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n543), .A2(new_n552), .A3(new_n554), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT72), .B(KEYINPUT36), .Z(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(KEYINPUT72), .A2(KEYINPUT36), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n568), .B1(new_n560), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n404), .A2(new_n408), .A3(new_n406), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(new_n418), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT39), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n419), .A2(new_n420), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n409), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n436), .B1(new_n572), .B2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n571), .A2(new_n573), .A3(new_n418), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT40), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n437), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT86), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n581), .B1(new_n578), .B2(new_n579), .ZN(new_n582));
  AOI211_X1 g381(.A(KEYINPUT86), .B(KEYINPUT40), .C1(new_n576), .C2(new_n577), .ZN(new_n583));
  OR4_X1    g382(.A1(new_n526), .A2(new_n580), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n517), .B1(new_n511), .B2(KEYINPUT37), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT87), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n511), .A2(KEYINPUT37), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n585), .A2(KEYINPUT87), .ZN(new_n589));
  OAI21_X1  g388(.A(KEYINPUT38), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n440), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT38), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n507), .B1(new_n500), .B2(new_n505), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n307), .B(new_n508), .C1(new_n509), .C2(new_n502), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(KEYINPUT37), .A3(new_n594), .ZN(new_n595));
  NAND4_X1  g394(.A1(new_n587), .A2(new_n592), .A3(new_n515), .A4(new_n595), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n590), .A2(new_n591), .A3(new_n520), .A4(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n570), .B1(new_n584), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g397(.A1(new_n561), .A2(new_n562), .B1(new_n598), .B2(new_n381), .ZN(new_n599));
  OR2_X1    g398(.A1(new_n519), .A2(KEYINPUT77), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n524), .A2(new_n525), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n519), .A2(KEYINPUT77), .ZN(new_n602));
  NAND4_X1  g401(.A1(new_n440), .A2(new_n600), .A3(new_n601), .A4(new_n602), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT82), .ZN(new_n604));
  OR2_X1    g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  AND2_X1   g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n565), .A2(new_n566), .ZN(new_n608));
  AOI211_X1 g407(.A(new_n562), .B(new_n608), .C1(new_n379), .C2(new_n380), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n381), .A2(new_n570), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  AOI21_X1  g410(.A(new_n279), .B1(new_n599), .B2(new_n611), .ZN(new_n612));
  XOR2_X1   g411(.A(G183gat), .B(G211gat), .Z(new_n613));
  INV_X1    g412(.A(KEYINPUT9), .ZN(new_n614));
  INV_X1    g413(.A(G64gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(G57gat), .ZN(new_n616));
  INV_X1    g415(.A(G57gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(G64gat), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n614), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g418(.A(KEYINPUT100), .B1(G71gat), .B2(G78gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(G71gat), .A2(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NOR3_X1   g421(.A1(KEYINPUT100), .A2(G71gat), .A3(G78gat), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n619), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  OR3_X1    g423(.A1(new_n617), .A2(KEYINPUT101), .A3(G64gat), .ZN(new_n625));
  OAI21_X1  g424(.A(G64gat), .B1(new_n617), .B2(KEYINPUT101), .ZN(new_n626));
  INV_X1    g425(.A(G71gat), .ZN(new_n627));
  INV_X1    g426(.A(G78gat), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n627), .A2(new_n628), .A3(KEYINPUT9), .ZN(new_n629));
  AOI22_X1  g428(.A1(new_n625), .A2(new_n626), .B1(new_n621), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n624), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n631), .A2(KEYINPUT21), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT102), .ZN(new_n633));
  NAND2_X1  g432(.A1(G231gat), .A2(G233gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G127gat), .B(G155gat), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g436(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n636), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n635), .B(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n638), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n241), .B1(KEYINPUT21), .B2(new_n631), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n639), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n645), .B1(new_n639), .B2(new_n643), .ZN(new_n648));
  OAI21_X1  g447(.A(new_n613), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n639), .A2(new_n643), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n644), .ZN(new_n651));
  INV_X1    g450(.A(new_n613), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n651), .A2(new_n646), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n649), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(G232gat), .A2(G233gat), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(KEYINPUT41), .ZN(new_n656));
  NOR2_X1   g455(.A1(KEYINPUT103), .A2(KEYINPUT7), .ZN(new_n657));
  NAND2_X1  g456(.A1(G85gat), .A2(G92gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI211_X1 g458(.A(G85gat), .B(G92gat), .C1(KEYINPUT103), .C2(KEYINPUT7), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n659), .A2(new_n660), .B1(KEYINPUT103), .B2(KEYINPUT7), .ZN(new_n661));
  NAND2_X1  g460(.A1(G99gat), .A2(G106gat), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT8), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n663), .B1(G85gat), .B2(G92gat), .ZN(new_n664));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g464(.A(G99gat), .B(G106gat), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n667), .B1(KEYINPUT104), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n668), .A2(KEYINPUT104), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n228), .A2(new_n245), .A3(new_n672), .ZN(new_n673));
  AOI22_X1  g472(.A1(new_n671), .A2(new_n222), .B1(KEYINPUT41), .B2(new_n655), .ZN(new_n674));
  XNOR2_X1  g473(.A(G190gat), .B(G218gat), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n673), .A2(new_n674), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n676), .B1(new_n673), .B2(new_n674), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n656), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n679), .ZN(new_n681));
  INV_X1    g480(.A(new_n656), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n681), .A2(new_n682), .A3(new_n677), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g483(.A(G134gat), .B(G162gat), .Z(new_n685));
  NAND2_X1  g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n685), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n680), .A2(new_n683), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n654), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(G230gat), .A2(G233gat), .ZN(new_n691));
  INV_X1    g490(.A(new_n631), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n692), .B1(new_n669), .B2(new_n670), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT10), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n667), .A2(new_n631), .A3(new_n668), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n693), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n671), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(KEYINPUT105), .ZN(new_n699));
  INV_X1    g498(.A(KEYINPUT105), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n700), .B1(new_n696), .B2(new_n697), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n691), .B1(new_n699), .B2(new_n701), .ZN(new_n702));
  AOI21_X1  g501(.A(new_n691), .B1(new_n693), .B2(new_n695), .ZN(new_n703));
  XOR2_X1   g502(.A(G120gat), .B(G148gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(KEYINPUT106), .ZN(new_n705));
  XOR2_X1   g504(.A(G176gat), .B(G204gat), .Z(new_n706));
  XNOR2_X1  g505(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n702), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n698), .A2(new_n691), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n707), .B1(new_n711), .B2(new_n703), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n709), .A2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n612), .A2(new_n690), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n715), .A2(new_n591), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(G1gat), .ZN(G1324gat));
  INV_X1    g516(.A(new_n526), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT42), .B1(new_n720), .B2(new_n239), .ZN(new_n721));
  XOR2_X1   g520(.A(KEYINPUT16), .B(G8gat), .Z(new_n722));
  NAND2_X1  g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  MUX2_X1   g522(.A(KEYINPUT42), .B(new_n721), .S(new_n723), .Z(G1325gat));
  INV_X1    g523(.A(G15gat), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n715), .A2(new_n725), .A3(new_n560), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n715), .A2(new_n570), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n726), .B1(new_n727), .B2(new_n725), .ZN(G1326gat));
  INV_X1    g527(.A(new_n381), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n715), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT43), .B(G22gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n730), .B(new_n731), .ZN(G1327gat));
  AND4_X1   g531(.A1(new_n612), .A2(new_n654), .A3(new_n689), .A4(new_n714), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n733), .A2(new_n202), .A3(new_n591), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(KEYINPUT45), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n561), .A2(new_n562), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n598), .A2(new_n381), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n605), .A2(new_n606), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n381), .A2(KEYINPUT35), .A3(new_n560), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n608), .A2(KEYINPUT72), .A3(KEYINPUT36), .ZN(new_n741));
  NAND4_X1  g540(.A1(new_n379), .A2(new_n741), .A3(new_n380), .A4(new_n568), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n739), .B1(new_n740), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n689), .B1(new_n738), .B2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n599), .A2(new_n611), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n747), .A2(KEYINPUT44), .A3(new_n689), .ZN(new_n748));
  AND2_X1   g547(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n654), .B(KEYINPUT107), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n750), .A2(new_n279), .A3(new_n713), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  OAI21_X1  g551(.A(G29gat), .B1(new_n752), .B2(new_n440), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n753), .ZN(G1328gat));
  OAI21_X1  g553(.A(G36gat), .B1(new_n752), .B2(new_n526), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n733), .A2(new_n203), .A3(new_n718), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT108), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT46), .ZN(new_n758));
  AND2_X1   g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n755), .B1(new_n759), .B2(new_n760), .ZN(G1329gat));
  NAND3_X1  g560(.A1(new_n749), .A2(new_n570), .A3(new_n751), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G43gat), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT47), .B1(new_n763), .B2(KEYINPUT109), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n733), .A2(new_n207), .A3(new_n560), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n764), .B(new_n766), .ZN(G1330gat));
  OAI21_X1  g566(.A(G50gat), .B1(new_n752), .B2(new_n381), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n733), .A2(new_n205), .A3(new_n729), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI21_X1  g569(.A(KEYINPUT48), .B1(new_n769), .B2(KEYINPUT110), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n770), .B(new_n771), .ZN(G1331gat));
  AND4_X1   g571(.A1(new_n279), .A2(new_n747), .A3(new_n690), .A4(new_n713), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(new_n591), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n774), .B(G57gat), .ZN(G1332gat));
  INV_X1    g574(.A(KEYINPUT49), .ZN(new_n776));
  OAI211_X1 g575(.A(new_n773), .B(new_n718), .C1(new_n776), .C2(new_n615), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n615), .ZN(new_n778));
  XNOR2_X1  g577(.A(new_n777), .B(new_n778), .ZN(G1333gat));
  AOI21_X1  g578(.A(G71gat), .B1(new_n773), .B2(new_n560), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n627), .B1(new_n741), .B2(new_n568), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n773), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g582(.A1(new_n773), .A2(new_n729), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT111), .B(G78gat), .Z(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1335gat));
  NAND2_X1  g585(.A1(new_n279), .A2(new_n654), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n714), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n749), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G85gat), .B1(new_n789), .B2(new_n440), .ZN(new_n790));
  INV_X1    g589(.A(new_n787), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n689), .B(new_n791), .C1(new_n738), .C2(new_n743), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n689), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n599), .B2(new_n611), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT51), .B1(new_n796), .B2(new_n791), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n714), .A2(G85gat), .A3(new_n440), .ZN(new_n799));
  XOR2_X1   g598(.A(new_n799), .B(KEYINPUT112), .Z(new_n800));
  OAI21_X1  g599(.A(new_n790), .B1(new_n798), .B2(new_n800), .ZN(G1336gat));
  INV_X1    g600(.A(KEYINPUT115), .ZN(new_n802));
  XOR2_X1   g601(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n803));
  NAND2_X1  g602(.A1(new_n792), .A2(new_n793), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n796), .A2(KEYINPUT51), .A3(new_n791), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n714), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n526), .A2(G92gat), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n803), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g607(.A1(new_n746), .A2(new_n718), .A3(new_n748), .A4(new_n788), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G92gat), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n802), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  OAI211_X1 g610(.A(new_n713), .B(new_n807), .C1(new_n794), .C2(new_n797), .ZN(new_n812));
  INV_X1    g611(.A(new_n803), .ZN(new_n813));
  AND4_X1   g612(.A1(new_n802), .A2(new_n810), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n811), .A2(new_n814), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT52), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n812), .A2(KEYINPUT113), .B1(G92gat), .B2(new_n809), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n806), .A2(new_n818), .A3(new_n807), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n816), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(KEYINPUT116), .B1(new_n815), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n808), .A2(new_n810), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n802), .A3(new_n810), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT116), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n817), .A2(new_n819), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT52), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n825), .A2(new_n826), .A3(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n821), .A2(new_n829), .ZN(G1337gat));
  INV_X1    g629(.A(new_n789), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(G99gat), .A3(new_n570), .ZN(new_n832));
  AND2_X1   g631(.A1(new_n806), .A2(new_n560), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n832), .B1(G99gat), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT117), .ZN(G1338gat));
  NAND3_X1  g634(.A1(new_n831), .A2(G106gat), .A3(new_n729), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n806), .A2(new_n729), .ZN(new_n837));
  OAI21_X1  g636(.A(new_n836), .B1(G106gat), .B2(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT53), .ZN(new_n839));
  XNOR2_X1  g638(.A(new_n838), .B(new_n839), .ZN(G1339gat));
  NOR2_X1   g639(.A1(new_n271), .A2(new_n250), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n256), .A2(new_n257), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n264), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n266), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n686), .B2(new_n688), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT118), .ZN(new_n846));
  INV_X1    g645(.A(new_n691), .ZN(new_n847));
  AOI211_X1 g646(.A(KEYINPUT54), .B(new_n847), .C1(new_n696), .C2(new_n697), .ZN(new_n848));
  INV_X1    g647(.A(new_n707), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT118), .B(new_n707), .C1(new_n710), .C2(KEYINPUT54), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n696), .A2(new_n847), .A3(new_n697), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n702), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT55), .ZN(new_n856));
  AND3_X1   g655(.A1(new_n852), .A2(new_n855), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n852), .B2(new_n855), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n709), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT119), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT119), .ZN(new_n861));
  OAI211_X1 g660(.A(new_n709), .B(new_n861), .C1(new_n857), .C2(new_n858), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n845), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT120), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n845), .A2(new_n860), .A3(KEYINPUT120), .A4(new_n862), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n860), .A2(new_n278), .A3(new_n862), .ZN(new_n868));
  INV_X1    g667(.A(new_n844), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n869), .A2(new_n713), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n795), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n750), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n690), .A2(new_n279), .A3(new_n714), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n718), .A2(new_n440), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n729), .A2(new_n608), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n279), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(new_n393), .ZN(G1340gat));
  NOR2_X1   g682(.A1(new_n881), .A2(new_n714), .ZN(new_n884));
  XNOR2_X1  g683(.A(new_n884), .B(new_n395), .ZN(G1341gat));
  INV_X1    g684(.A(new_n750), .ZN(new_n886));
  OAI21_X1  g685(.A(G127gat), .B1(new_n881), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n654), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n399), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n881), .B2(new_n889), .ZN(G1342gat));
  NAND2_X1  g689(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n891));
  NAND4_X1  g690(.A1(new_n879), .A2(new_n880), .A3(new_n689), .A4(new_n891), .ZN(new_n892));
  NOR2_X1   g691(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n893));
  XOR2_X1   g692(.A(new_n892), .B(new_n893), .Z(G1343gat));
  AND2_X1   g693(.A1(new_n865), .A2(new_n866), .ZN(new_n895));
  INV_X1    g694(.A(new_n859), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n278), .A2(new_n896), .B1(new_n713), .B2(new_n869), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n897), .A2(new_n689), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n654), .B1(new_n895), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(new_n874), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n900), .A2(KEYINPUT57), .A3(new_n729), .ZN(new_n901));
  XNOR2_X1  g700(.A(KEYINPUT121), .B(KEYINPUT57), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n902), .B1(new_n876), .B2(new_n381), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n878), .A2(new_n570), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(G141gat), .B1(new_n906), .B2(new_n279), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT58), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n879), .A2(new_n610), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n909), .A2(G141gat), .A3(new_n279), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n907), .A2(new_n908), .A3(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(new_n905), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n913), .B1(new_n901), .B2(new_n903), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n315), .B1(new_n914), .B2(new_n278), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT58), .B1(new_n915), .B2(new_n910), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n912), .A2(new_n916), .ZN(G1344gat));
  NAND4_X1  g716(.A1(new_n879), .A2(new_n335), .A3(new_n610), .A4(new_n713), .ZN(new_n918));
  AOI211_X1 g717(.A(KEYINPUT59), .B(new_n335), .C1(new_n914), .C2(new_n713), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT59), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n867), .A2(new_n872), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n874), .B1(new_n921), .B2(new_n750), .ZN(new_n922));
  INV_X1    g721(.A(new_n902), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n922), .A2(new_n729), .A3(new_n923), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n845), .A2(new_n896), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n926), .B1(new_n897), .B2(new_n689), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n875), .B1(new_n927), .B2(new_n654), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n925), .B1(new_n928), .B2(new_n381), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n924), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n930), .A2(new_n713), .A3(new_n905), .ZN(new_n931));
  AOI21_X1  g730(.A(new_n920), .B1(new_n931), .B2(G148gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n918), .B1(new_n919), .B2(new_n932), .ZN(G1345gat));
  NOR3_X1   g732(.A1(new_n909), .A2(KEYINPUT122), .A3(new_n654), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(G155gat), .ZN(new_n935));
  OAI21_X1  g734(.A(KEYINPUT122), .B1(new_n909), .B2(new_n654), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n750), .A2(G155gat), .ZN(new_n937));
  AOI22_X1  g736(.A1(new_n935), .A2(new_n936), .B1(new_n914), .B2(new_n937), .ZN(G1346gat));
  OAI21_X1  g737(.A(G162gat), .B1(new_n906), .B2(new_n795), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n742), .A2(G162gat), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n922), .A2(new_n689), .A3(new_n877), .A4(new_n940), .ZN(new_n941));
  XNOR2_X1  g740(.A(new_n941), .B(KEYINPUT123), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n939), .A2(new_n943), .A3(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(G162gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n914), .B2(new_n689), .ZN(new_n947));
  OAI21_X1  g746(.A(KEYINPUT124), .B1(new_n947), .B2(new_n942), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n945), .A2(new_n948), .ZN(G1347gat));
  NOR2_X1   g748(.A1(new_n591), .A2(new_n526), .ZN(new_n950));
  OAI211_X1 g749(.A(new_n880), .B(new_n950), .C1(new_n873), .C2(new_n875), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n279), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(new_n261), .ZN(G1348gat));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n714), .ZN(new_n954));
  XNOR2_X1  g753(.A(new_n954), .B(new_n482), .ZN(G1349gat));
  OAI21_X1  g754(.A(G183gat), .B1(new_n951), .B2(new_n886), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n888), .A2(new_n477), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n951), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g758(.A(G190gat), .B1(new_n951), .B2(new_n795), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n960), .A2(KEYINPUT125), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  OAI211_X1 g762(.A(new_n963), .B(G190gat), .C1(new_n951), .C2(new_n795), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n961), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n961), .A2(new_n967), .A3(new_n962), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n961), .A2(new_n964), .ZN(new_n969));
  NAND2_X1  g768(.A1(new_n969), .A2(KEYINPUT61), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n966), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  INV_X1    g770(.A(new_n950), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n876), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n973), .A2(new_n475), .A3(new_n880), .A4(new_n689), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n971), .A2(new_n974), .ZN(G1351gat));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n610), .ZN(new_n976));
  INV_X1    g775(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g776(.A(G197gat), .B1(new_n977), .B2(new_n278), .ZN(new_n978));
  NOR2_X1   g777(.A1(new_n972), .A2(new_n570), .ZN(new_n979));
  INV_X1    g778(.A(new_n979), .ZN(new_n980));
  AOI21_X1  g779(.A(new_n980), .B1(new_n924), .B2(new_n929), .ZN(new_n981));
  AND2_X1   g780(.A1(new_n278), .A2(G197gat), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n978), .B1(new_n981), .B2(new_n982), .ZN(G1352gat));
  OR2_X1    g782(.A1(new_n714), .A2(G204gat), .ZN(new_n984));
  OAI21_X1  g783(.A(KEYINPUT62), .B1(new_n976), .B2(new_n984), .ZN(new_n985));
  INV_X1    g784(.A(KEYINPUT127), .ZN(new_n986));
  XNOR2_X1  g785(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NOR3_X1   g786(.A1(new_n976), .A2(KEYINPUT62), .A3(new_n984), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n930), .A2(new_n713), .A3(new_n979), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n988), .B1(G204gat), .B2(new_n989), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n987), .A2(new_n990), .ZN(G1353gat));
  NAND3_X1  g790(.A1(new_n977), .A2(new_n292), .A3(new_n888), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n981), .A2(new_n888), .ZN(new_n993));
  AND3_X1   g792(.A1(new_n993), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n994));
  AOI21_X1  g793(.A(KEYINPUT63), .B1(new_n993), .B2(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(G1354gat));
  NAND3_X1  g795(.A1(new_n977), .A2(new_n283), .A3(new_n689), .ZN(new_n997));
  AND2_X1   g796(.A1(new_n981), .A2(new_n689), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n997), .B1(new_n998), .B2(new_n283), .ZN(G1355gat));
endmodule


