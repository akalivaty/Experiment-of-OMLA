

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U553 ( .A1(n839), .A2(n764), .ZN(n783) );
  XNOR2_X1 U554 ( .A(n551), .B(n571), .ZN(n763) );
  XNOR2_X2 U555 ( .A(n827), .B(n826), .ZN(n593) );
  AND2_X2 U556 ( .A1(n556), .A2(n574), .ZN(n558) );
  INV_X1 U557 ( .A(n1039), .ZN(n541) );
  AND2_X1 U558 ( .A1(n532), .A2(n531), .ZN(n799) );
  NAND2_X1 U559 ( .A1(n538), .A2(n785), .ZN(n795) );
  NOR2_X2 U560 ( .A1(n676), .A2(n675), .ZN(n1028) );
  XNOR2_X1 U561 ( .A(n561), .B(KEYINPUT17), .ZN(n698) );
  NOR2_X2 U562 ( .A1(n734), .A2(n613), .ZN(n722) );
  INV_X1 U563 ( .A(G2105), .ZN(n562) );
  NAND2_X1 U564 ( .A1(n788), .A2(G1956), .ZN(n542) );
  NOR2_X1 U565 ( .A1(n783), .A2(n979), .ZN(n782) );
  INV_X1 U566 ( .A(G8), .ZN(n765) );
  INV_X1 U567 ( .A(KEYINPUT101), .ZN(n603) );
  INV_X1 U568 ( .A(n833), .ZN(n590) );
  NAND2_X1 U569 ( .A1(n833), .A2(n586), .ZN(n585) );
  NAND2_X1 U570 ( .A1(n587), .A2(n589), .ZN(n586) );
  INV_X1 U571 ( .A(n1024), .ZN(n587) );
  NOR2_X1 U572 ( .A1(n572), .A2(n520), .ZN(n552) );
  AND2_X1 U573 ( .A1(n698), .A2(G138), .ZN(n572) );
  INV_X1 U574 ( .A(n795), .ZN(n537) );
  INV_X1 U575 ( .A(G168), .ZN(n568) );
  NOR2_X1 U576 ( .A1(n773), .A2(n772), .ZN(n775) );
  XNOR2_X1 U577 ( .A(n801), .B(KEYINPUT28), .ZN(n549) );
  INV_X1 U578 ( .A(KEYINPUT29), .ZN(n548) );
  NOR2_X1 U579 ( .A1(n604), .A2(n603), .ZN(n602) );
  NAND2_X1 U580 ( .A1(n600), .A2(n599), .ZN(n598) );
  NAND2_X1 U581 ( .A1(n601), .A2(n603), .ZN(n600) );
  NAND2_X1 U582 ( .A1(n821), .A2(n522), .ZN(n599) );
  INV_X1 U583 ( .A(n821), .ZN(n601) );
  AND2_X1 U584 ( .A1(n1024), .A2(KEYINPUT103), .ZN(n592) );
  NAND2_X1 U585 ( .A1(n832), .A2(n836), .ZN(n833) );
  INV_X1 U586 ( .A(KEYINPUT103), .ZN(n589) );
  AND2_X1 U587 ( .A1(n578), .A2(n869), .ZN(n577) );
  NAND2_X1 U588 ( .A1(n579), .A2(n868), .ZN(n578) );
  INV_X1 U589 ( .A(n525), .ZN(n579) );
  INV_X1 U590 ( .A(KEYINPUT106), .ZN(n573) );
  NAND2_X1 U591 ( .A1(n563), .A2(n562), .ZN(n561) );
  INV_X1 U592 ( .A(G2104), .ZN(n563) );
  XNOR2_X1 U593 ( .A(n629), .B(n628), .ZN(n631) );
  INV_X1 U594 ( .A(KEYINPUT64), .ZN(n627) );
  NAND2_X1 U595 ( .A1(G2067), .A2(n784), .ZN(n785) );
  INV_X1 U596 ( .A(G299), .ZN(n539) );
  NOR2_X1 U597 ( .A1(n794), .A2(n793), .ZN(n797) );
  AND2_X1 U598 ( .A1(n783), .A2(n769), .ZN(n770) );
  NAND2_X1 U599 ( .A1(n570), .A2(n567), .ZN(n566) );
  AND2_X1 U600 ( .A1(n565), .A2(G8), .ZN(n564) );
  INV_X1 U601 ( .A(G1966), .ZN(n565) );
  XNOR2_X1 U602 ( .A(n535), .B(n548), .ZN(n534) );
  NAND2_X1 U603 ( .A1(n596), .A2(n523), .ZN(n595) );
  AND2_X1 U604 ( .A1(n591), .A2(n584), .ZN(n583) );
  NAND2_X1 U605 ( .A1(n582), .A2(n524), .ZN(n581) );
  NAND2_X1 U606 ( .A1(n776), .A2(G8), .ZN(n836) );
  NAND2_X1 U607 ( .A1(n533), .A2(n668), .ZN(n670) );
  NAND2_X1 U608 ( .A1(n519), .A2(n555), .ZN(n557) );
  NAND2_X1 U609 ( .A1(n576), .A2(n868), .ZN(n555) );
  XNOR2_X1 U610 ( .A(n684), .B(KEYINPUT15), .ZN(n1039) );
  INV_X1 U611 ( .A(KEYINPUT86), .ZN(n571) );
  NOR2_X1 U612 ( .A1(n637), .A2(n636), .ZN(G160) );
  XNOR2_X1 U613 ( .A(n566), .B(n527), .ZN(n809) );
  AND2_X1 U614 ( .A1(n575), .A2(n529), .ZN(n519) );
  AND2_X1 U615 ( .A1(G102), .A2(n939), .ZN(n520) );
  BUF_X1 U616 ( .A(n783), .Z(n776) );
  INV_X1 U617 ( .A(G2105), .ZN(n632) );
  BUF_X2 U618 ( .A(n783), .Z(n788) );
  AND2_X1 U619 ( .A1(n542), .A2(n539), .ZN(n521) );
  OR2_X1 U620 ( .A1(n817), .A2(KEYINPUT101), .ZN(n522) );
  AND2_X1 U621 ( .A1(n821), .A2(n603), .ZN(n523) );
  AND2_X1 U622 ( .A1(n776), .A2(n564), .ZN(n813) );
  AND2_X1 U623 ( .A1(n833), .A2(n589), .ZN(n524) );
  AND2_X1 U624 ( .A1(n877), .A2(n870), .ZN(n525) );
  XOR2_X1 U625 ( .A(KEYINPUT96), .B(KEYINPUT30), .Z(n526) );
  XOR2_X1 U626 ( .A(KEYINPUT31), .B(KEYINPUT97), .Z(n527) );
  AND2_X1 U627 ( .A1(n525), .A2(KEYINPUT105), .ZN(n528) );
  AND2_X1 U628 ( .A1(n577), .A2(n573), .ZN(n529) );
  INV_X1 U629 ( .A(KEYINPUT105), .ZN(n868) );
  AND2_X1 U630 ( .A1(n868), .A2(KEYINPUT106), .ZN(n530) );
  NAND2_X1 U631 ( .A1(n537), .A2(n541), .ZN(n531) );
  NAND2_X1 U632 ( .A1(n521), .A2(n540), .ZN(n532) );
  XNOR2_X1 U633 ( .A(n547), .B(KEYINPUT32), .ZN(n544) );
  XNOR2_X1 U634 ( .A(n666), .B(n667), .ZN(n533) );
  NOR2_X2 U635 ( .A1(G543), .A2(G651), .ZN(n719) );
  NAND2_X1 U636 ( .A1(n534), .A2(n803), .ZN(n810) );
  NAND2_X1 U637 ( .A1(n536), .A2(n549), .ZN(n535) );
  XNOR2_X1 U638 ( .A(n800), .B(n550), .ZN(n536) );
  XNOR2_X1 U639 ( .A(n782), .B(n781), .ZN(n540) );
  NAND2_X1 U640 ( .A1(n788), .A2(G1348), .ZN(n538) );
  NAND2_X1 U641 ( .A1(n540), .A2(n542), .ZN(n560) );
  XNOR2_X2 U642 ( .A(n543), .B(KEYINPUT100), .ZN(n829) );
  NAND2_X1 U643 ( .A1(n545), .A2(n544), .ZN(n543) );
  NAND2_X1 U644 ( .A1(n546), .A2(n605), .ZN(n545) );
  XNOR2_X1 U645 ( .A(n811), .B(KEYINPUT98), .ZN(n546) );
  NAND2_X1 U646 ( .A1(n808), .A2(n607), .ZN(n547) );
  INV_X1 U647 ( .A(KEYINPUT95), .ZN(n550) );
  NAND2_X1 U648 ( .A1(n553), .A2(n552), .ZN(n551) );
  XNOR2_X1 U649 ( .A(n554), .B(KEYINPUT85), .ZN(n553) );
  NAND2_X1 U650 ( .A1(n655), .A2(n654), .ZN(n554) );
  NAND2_X1 U651 ( .A1(n575), .A2(n577), .ZN(n559) );
  NAND2_X1 U652 ( .A1(n559), .A2(KEYINPUT106), .ZN(n556) );
  NAND2_X1 U653 ( .A1(n558), .A2(n557), .ZN(n883) );
  NAND2_X1 U654 ( .A1(n560), .A2(G299), .ZN(n801) );
  NAND2_X1 U655 ( .A1(n569), .A2(n568), .ZN(n567) );
  XNOR2_X1 U656 ( .A(n768), .B(n526), .ZN(n569) );
  OR2_X2 U657 ( .A1(n802), .A2(G171), .ZN(n570) );
  XNOR2_X1 U658 ( .A(n775), .B(n774), .ZN(n802) );
  NAND2_X1 U659 ( .A1(n576), .A2(n530), .ZN(n574) );
  NAND2_X1 U660 ( .A1(n580), .A2(n528), .ZN(n575) );
  INV_X1 U661 ( .A(n580), .ZN(n576) );
  NAND2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n588), .A2(n585), .ZN(n584) );
  XNOR2_X2 U664 ( .A(n838), .B(KEYINPUT104), .ZN(n580) );
  NAND2_X1 U665 ( .A1(n583), .A2(n581), .ZN(n837) );
  INV_X1 U666 ( .A(n593), .ZN(n582) );
  NAND2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n591) );
  AND2_X1 U668 ( .A1(n594), .A2(n598), .ZN(n597) );
  NAND2_X1 U669 ( .A1(n829), .A2(n602), .ZN(n594) );
  NAND2_X1 U670 ( .A1(n597), .A2(n595), .ZN(n825) );
  INV_X1 U671 ( .A(n829), .ZN(n596) );
  INV_X1 U672 ( .A(n817), .ZN(n604) );
  AND2_X1 U673 ( .A1(n815), .A2(n814), .ZN(n605) );
  OR2_X1 U674 ( .A1(n836), .A2(n835), .ZN(n606) );
  AND2_X1 U675 ( .A1(n807), .A2(G8), .ZN(n607) );
  AND2_X1 U676 ( .A1(n789), .A2(G1996), .ZN(n790) );
  NAND2_X1 U677 ( .A1(n784), .A2(n790), .ZN(n791) );
  INV_X1 U678 ( .A(KEYINPUT102), .ZN(n826) );
  XNOR2_X1 U679 ( .A(KEYINPUT13), .B(KEYINPUT70), .ZN(n669) );
  XNOR2_X1 U680 ( .A(n670), .B(n669), .ZN(n673) );
  XNOR2_X1 U681 ( .A(n627), .B(KEYINPUT23), .ZN(n628) );
  OR2_X1 U682 ( .A1(n626), .A2(n625), .ZN(G299) );
  NAND2_X1 U683 ( .A1(n719), .A2(G89), .ZN(n608) );
  XNOR2_X1 U684 ( .A(KEYINPUT4), .B(n608), .ZN(n611) );
  XOR2_X1 U685 ( .A(G543), .B(KEYINPUT0), .Z(n734) );
  INV_X1 U686 ( .A(G651), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n722), .A2(G76), .ZN(n609) );
  XOR2_X1 U688 ( .A(KEYINPUT75), .B(n609), .Z(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n612) );
  XNOR2_X1 U690 ( .A(n612), .B(KEYINPUT5), .ZN(n619) );
  NOR2_X1 U691 ( .A1(G543), .A2(n613), .ZN(n614) );
  XOR2_X2 U692 ( .A(KEYINPUT1), .B(n614), .Z(n733) );
  NAND2_X1 U693 ( .A1(G63), .A2(n733), .ZN(n616) );
  NOR2_X2 U694 ( .A1(G651), .A2(n734), .ZN(n729) );
  NAND2_X1 U695 ( .A1(G51), .A2(n729), .ZN(n615) );
  NAND2_X1 U696 ( .A1(n616), .A2(n615), .ZN(n617) );
  XOR2_X1 U697 ( .A(KEYINPUT6), .B(n617), .Z(n618) );
  NAND2_X1 U698 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U699 ( .A(n620), .B(KEYINPUT7), .ZN(G168) );
  NAND2_X1 U700 ( .A1(G65), .A2(n733), .ZN(n622) );
  NAND2_X1 U701 ( .A1(G53), .A2(n729), .ZN(n621) );
  NAND2_X1 U702 ( .A1(n622), .A2(n621), .ZN(n626) );
  NAND2_X1 U703 ( .A1(G78), .A2(n722), .ZN(n624) );
  NAND2_X1 U704 ( .A1(G91), .A2(n719), .ZN(n623) );
  NAND2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n625) );
  AND2_X4 U706 ( .A1(n562), .A2(G2104), .ZN(n939) );
  NAND2_X1 U707 ( .A1(G101), .A2(n939), .ZN(n629) );
  NAND2_X1 U708 ( .A1(G137), .A2(n698), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n637) );
  NOR2_X2 U710 ( .A1(n632), .A2(G2104), .ZN(n651) );
  BUF_X1 U711 ( .A(n651), .Z(n942) );
  NAND2_X1 U712 ( .A1(G125), .A2(n942), .ZN(n635) );
  NAND2_X1 U713 ( .A1(G2105), .A2(G2104), .ZN(n633) );
  XNOR2_X1 U714 ( .A(n633), .B(KEYINPUT65), .ZN(n653) );
  BUF_X1 U715 ( .A(n653), .Z(n943) );
  NAND2_X1 U716 ( .A1(G113), .A2(n943), .ZN(n634) );
  NAND2_X1 U717 ( .A1(n635), .A2(n634), .ZN(n636) );
  NAND2_X1 U718 ( .A1(G64), .A2(n733), .ZN(n639) );
  NAND2_X1 U719 ( .A1(G52), .A2(n729), .ZN(n638) );
  NAND2_X1 U720 ( .A1(n639), .A2(n638), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G77), .A2(n722), .ZN(n641) );
  NAND2_X1 U722 ( .A1(G90), .A2(n719), .ZN(n640) );
  NAND2_X1 U723 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U724 ( .A(KEYINPUT9), .B(n642), .Z(n643) );
  NOR2_X1 U725 ( .A1(n644), .A2(n643), .ZN(G171) );
  NAND2_X1 U726 ( .A1(G60), .A2(n733), .ZN(n646) );
  NAND2_X1 U727 ( .A1(G47), .A2(n729), .ZN(n645) );
  NAND2_X1 U728 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U729 ( .A1(G72), .A2(n722), .ZN(n648) );
  NAND2_X1 U730 ( .A1(G85), .A2(n719), .ZN(n647) );
  NAND2_X1 U731 ( .A1(n648), .A2(n647), .ZN(n649) );
  OR2_X1 U732 ( .A1(n650), .A2(n649), .ZN(G290) );
  NAND2_X1 U733 ( .A1(n651), .A2(G126), .ZN(n652) );
  XNOR2_X1 U734 ( .A(n652), .B(KEYINPUT84), .ZN(n655) );
  NAND2_X1 U735 ( .A1(G114), .A2(n653), .ZN(n654) );
  BUF_X1 U736 ( .A(n763), .Z(G164) );
  AND2_X1 U737 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U738 ( .A(G132), .ZN(G219) );
  INV_X1 U739 ( .A(G108), .ZN(G238) );
  NAND2_X1 U740 ( .A1(G75), .A2(n722), .ZN(n656) );
  XNOR2_X1 U741 ( .A(n656), .B(KEYINPUT80), .ZN(n658) );
  NAND2_X1 U742 ( .A1(n729), .A2(G50), .ZN(n657) );
  NAND2_X1 U743 ( .A1(n658), .A2(n657), .ZN(n662) );
  NAND2_X1 U744 ( .A1(G62), .A2(n733), .ZN(n660) );
  NAND2_X1 U745 ( .A1(G88), .A2(n719), .ZN(n659) );
  NAND2_X1 U746 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U747 ( .A1(n662), .A2(n661), .ZN(G166) );
  XOR2_X1 U748 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U749 ( .A(KEYINPUT10), .B(KEYINPUT67), .Z(n664) );
  NAND2_X1 U750 ( .A1(G7), .A2(G661), .ZN(n663) );
  XNOR2_X1 U751 ( .A(n664), .B(n663), .ZN(G223) );
  XOR2_X1 U752 ( .A(G223), .B(KEYINPUT68), .Z(n885) );
  NAND2_X1 U753 ( .A1(n885), .A2(G567), .ZN(n665) );
  XOR2_X1 U754 ( .A(KEYINPUT11), .B(n665), .Z(G234) );
  NAND2_X1 U755 ( .A1(G68), .A2(n722), .ZN(n668) );
  XOR2_X1 U756 ( .A(KEYINPUT69), .B(KEYINPUT12), .Z(n667) );
  NAND2_X1 U757 ( .A1(G81), .A2(n719), .ZN(n666) );
  NAND2_X1 U758 ( .A1(G43), .A2(n729), .ZN(n671) );
  XOR2_X1 U759 ( .A(KEYINPUT71), .B(n671), .Z(n672) );
  NAND2_X1 U760 ( .A1(n673), .A2(n672), .ZN(n676) );
  NAND2_X1 U761 ( .A1(n733), .A2(G56), .ZN(n674) );
  XOR2_X1 U762 ( .A(KEYINPUT14), .B(n674), .Z(n675) );
  NAND2_X1 U763 ( .A1(G860), .A2(n1028), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n677), .B(KEYINPUT72), .ZN(G153) );
  NAND2_X1 U765 ( .A1(G79), .A2(n722), .ZN(n679) );
  NAND2_X1 U766 ( .A1(G92), .A2(n719), .ZN(n678) );
  NAND2_X1 U767 ( .A1(n679), .A2(n678), .ZN(n683) );
  NAND2_X1 U768 ( .A1(G66), .A2(n733), .ZN(n681) );
  NAND2_X1 U769 ( .A1(G54), .A2(n729), .ZN(n680) );
  NAND2_X1 U770 ( .A1(n681), .A2(n680), .ZN(n682) );
  NOR2_X1 U771 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U772 ( .A1(n541), .A2(G868), .ZN(n685) );
  XOR2_X1 U773 ( .A(KEYINPUT74), .B(n685), .Z(n688) );
  INV_X1 U774 ( .A(G868), .ZN(n695) );
  NOR2_X1 U775 ( .A1(G171), .A2(n695), .ZN(n686) );
  XNOR2_X1 U776 ( .A(KEYINPUT73), .B(n686), .ZN(n687) );
  NAND2_X1 U777 ( .A1(n688), .A2(n687), .ZN(G284) );
  NOR2_X1 U778 ( .A1(G286), .A2(n695), .ZN(n690) );
  NOR2_X1 U779 ( .A1(G868), .A2(G299), .ZN(n689) );
  NOR2_X1 U780 ( .A1(n690), .A2(n689), .ZN(G297) );
  INV_X1 U781 ( .A(G860), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n691), .A2(G559), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n692), .A2(n541), .ZN(n693) );
  XNOR2_X1 U784 ( .A(n693), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U785 ( .A1(n541), .A2(G868), .ZN(n694) );
  NOR2_X1 U786 ( .A1(G559), .A2(n694), .ZN(n697) );
  AND2_X1 U787 ( .A1(n695), .A2(n1028), .ZN(n696) );
  NOR2_X1 U788 ( .A1(n697), .A2(n696), .ZN(G282) );
  BUF_X1 U789 ( .A(n698), .Z(n938) );
  NAND2_X1 U790 ( .A1(G135), .A2(n938), .ZN(n699) );
  XNOR2_X1 U791 ( .A(n699), .B(KEYINPUT76), .ZN(n702) );
  NAND2_X1 U792 ( .A1(G123), .A2(n942), .ZN(n700) );
  XNOR2_X1 U793 ( .A(n700), .B(KEYINPUT18), .ZN(n701) );
  NAND2_X1 U794 ( .A1(n702), .A2(n701), .ZN(n706) );
  NAND2_X1 U795 ( .A1(G111), .A2(n943), .ZN(n704) );
  NAND2_X1 U796 ( .A1(G99), .A2(n939), .ZN(n703) );
  NAND2_X1 U797 ( .A1(n704), .A2(n703), .ZN(n705) );
  NOR2_X1 U798 ( .A1(n706), .A2(n705), .ZN(n1002) );
  XNOR2_X1 U799 ( .A(G2096), .B(n1002), .ZN(n708) );
  INV_X1 U800 ( .A(G2100), .ZN(n707) );
  NAND2_X1 U801 ( .A1(n708), .A2(n707), .ZN(G156) );
  NAND2_X1 U802 ( .A1(G55), .A2(n729), .ZN(n709) );
  XNOR2_X1 U803 ( .A(n709), .B(KEYINPUT78), .ZN(n712) );
  NAND2_X1 U804 ( .A1(G93), .A2(n719), .ZN(n710) );
  XOR2_X1 U805 ( .A(KEYINPUT77), .B(n710), .Z(n711) );
  NAND2_X1 U806 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U807 ( .A1(G67), .A2(n733), .ZN(n714) );
  NAND2_X1 U808 ( .A1(G80), .A2(n722), .ZN(n713) );
  NAND2_X1 U809 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U810 ( .A1(n716), .A2(n715), .ZN(n746) );
  NAND2_X1 U811 ( .A1(n541), .A2(G559), .ZN(n744) );
  XOR2_X1 U812 ( .A(n1028), .B(n744), .Z(n717) );
  NOR2_X1 U813 ( .A1(G860), .A2(n717), .ZN(n718) );
  XNOR2_X1 U814 ( .A(n746), .B(n718), .ZN(G145) );
  NAND2_X1 U815 ( .A1(G61), .A2(n733), .ZN(n721) );
  NAND2_X1 U816 ( .A1(G86), .A2(n719), .ZN(n720) );
  NAND2_X1 U817 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U818 ( .A1(n722), .A2(G73), .ZN(n723) );
  XOR2_X1 U819 ( .A(KEYINPUT2), .B(n723), .Z(n724) );
  NOR2_X1 U820 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U821 ( .A(KEYINPUT79), .B(n726), .Z(n728) );
  NAND2_X1 U822 ( .A1(n729), .A2(G48), .ZN(n727) );
  NAND2_X1 U823 ( .A1(n728), .A2(n727), .ZN(G305) );
  NAND2_X1 U824 ( .A1(G49), .A2(n729), .ZN(n731) );
  NAND2_X1 U825 ( .A1(G74), .A2(G651), .ZN(n730) );
  NAND2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  NOR2_X1 U827 ( .A1(n733), .A2(n732), .ZN(n736) );
  NAND2_X1 U828 ( .A1(n734), .A2(G87), .ZN(n735) );
  NAND2_X1 U829 ( .A1(n736), .A2(n735), .ZN(G288) );
  XNOR2_X1 U830 ( .A(n1028), .B(n746), .ZN(n738) );
  XNOR2_X1 U831 ( .A(G305), .B(G166), .ZN(n737) );
  XNOR2_X1 U832 ( .A(n738), .B(n737), .ZN(n741) );
  XOR2_X1 U833 ( .A(G290), .B(G299), .Z(n739) );
  XNOR2_X1 U834 ( .A(G288), .B(n739), .ZN(n740) );
  XOR2_X1 U835 ( .A(n741), .B(n740), .Z(n743) );
  XNOR2_X1 U836 ( .A(KEYINPUT81), .B(KEYINPUT19), .ZN(n742) );
  XNOR2_X1 U837 ( .A(n743), .B(n742), .ZN(n952) );
  XOR2_X1 U838 ( .A(n952), .B(n744), .Z(n745) );
  NAND2_X1 U839 ( .A1(G868), .A2(n745), .ZN(n748) );
  OR2_X1 U840 ( .A1(n746), .A2(G868), .ZN(n747) );
  NAND2_X1 U841 ( .A1(n748), .A2(n747), .ZN(G295) );
  NAND2_X1 U842 ( .A1(G2084), .A2(G2078), .ZN(n749) );
  XOR2_X1 U843 ( .A(KEYINPUT20), .B(n749), .Z(n750) );
  NAND2_X1 U844 ( .A1(G2090), .A2(n750), .ZN(n751) );
  XNOR2_X1 U845 ( .A(KEYINPUT21), .B(n751), .ZN(n752) );
  NAND2_X1 U846 ( .A1(n752), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U847 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U848 ( .A(KEYINPUT66), .B(G82), .Z(G220) );
  NAND2_X1 U849 ( .A1(G69), .A2(G120), .ZN(n753) );
  XNOR2_X1 U850 ( .A(KEYINPUT82), .B(n753), .ZN(n754) );
  NOR2_X1 U851 ( .A1(G238), .A2(n754), .ZN(n755) );
  NAND2_X1 U852 ( .A1(G57), .A2(n755), .ZN(n891) );
  NAND2_X1 U853 ( .A1(n891), .A2(G567), .ZN(n760) );
  NOR2_X1 U854 ( .A1(G220), .A2(G219), .ZN(n756) );
  XOR2_X1 U855 ( .A(KEYINPUT22), .B(n756), .Z(n757) );
  NOR2_X1 U856 ( .A1(G218), .A2(n757), .ZN(n758) );
  NAND2_X1 U857 ( .A1(G96), .A2(n758), .ZN(n890) );
  NAND2_X1 U858 ( .A1(n890), .A2(G2106), .ZN(n759) );
  NAND2_X1 U859 ( .A1(n760), .A2(n759), .ZN(n893) );
  NAND2_X1 U860 ( .A1(G483), .A2(G661), .ZN(n761) );
  NOR2_X1 U861 ( .A1(n893), .A2(n761), .ZN(n887) );
  NAND2_X1 U862 ( .A1(n887), .A2(G36), .ZN(n762) );
  XOR2_X1 U863 ( .A(KEYINPUT83), .B(n762), .Z(G176) );
  INV_X1 U864 ( .A(G166), .ZN(G303) );
  NOR2_X2 U865 ( .A1(n763), .A2(G1384), .ZN(n839) );
  NAND2_X1 U866 ( .A1(G160), .A2(G40), .ZN(n840) );
  INV_X1 U867 ( .A(n840), .ZN(n764) );
  NOR2_X1 U868 ( .A1(n813), .A2(n765), .ZN(n767) );
  NOR2_X1 U869 ( .A1(G2084), .A2(n788), .ZN(n812) );
  INV_X1 U870 ( .A(n812), .ZN(n766) );
  NAND2_X1 U871 ( .A1(n767), .A2(n766), .ZN(n768) );
  INV_X1 U872 ( .A(G1961), .ZN(n769) );
  XNOR2_X1 U873 ( .A(n770), .B(KEYINPUT90), .ZN(n773) );
  XNOR2_X1 U874 ( .A(G2078), .B(KEYINPUT25), .ZN(n771) );
  XNOR2_X1 U875 ( .A(n771), .B(KEYINPUT91), .ZN(n974) );
  NOR2_X1 U876 ( .A1(n788), .A2(n974), .ZN(n772) );
  INV_X1 U877 ( .A(KEYINPUT92), .ZN(n774) );
  NOR2_X1 U878 ( .A1(G2090), .A2(n776), .ZN(n777) );
  XNOR2_X1 U879 ( .A(KEYINPUT99), .B(n777), .ZN(n780) );
  NOR2_X1 U880 ( .A1(G1971), .A2(n836), .ZN(n778) );
  NOR2_X1 U881 ( .A1(G166), .A2(n778), .ZN(n779) );
  NAND2_X1 U882 ( .A1(n780), .A2(n779), .ZN(n805) );
  AND2_X1 U883 ( .A1(n809), .A2(n805), .ZN(n804) );
  INV_X1 U884 ( .A(G2072), .ZN(n979) );
  XOR2_X1 U885 ( .A(KEYINPUT93), .B(KEYINPUT27), .Z(n781) );
  INV_X1 U886 ( .A(n783), .ZN(n784) );
  XNOR2_X1 U887 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n789) );
  OR2_X1 U888 ( .A1(n789), .A2(G1996), .ZN(n786) );
  NAND2_X1 U889 ( .A1(n1028), .A2(n786), .ZN(n794) );
  INV_X1 U890 ( .A(G1341), .ZN(n1060) );
  NAND2_X1 U891 ( .A1(n1060), .A2(n789), .ZN(n787) );
  NAND2_X1 U892 ( .A1(n787), .A2(n788), .ZN(n792) );
  INV_X1 U893 ( .A(G1996), .ZN(n973) );
  NAND2_X1 U894 ( .A1(n792), .A2(n791), .ZN(n793) );
  NAND2_X1 U895 ( .A1(n795), .A2(n1039), .ZN(n796) );
  NAND2_X1 U896 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U897 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n802), .A2(G171), .ZN(n803) );
  NAND2_X1 U899 ( .A1(n804), .A2(n810), .ZN(n808) );
  INV_X1 U900 ( .A(n805), .ZN(n806) );
  OR2_X1 U901 ( .A1(n806), .A2(G286), .ZN(n807) );
  NAND2_X1 U902 ( .A1(n810), .A2(n809), .ZN(n811) );
  NAND2_X1 U903 ( .A1(G8), .A2(n812), .ZN(n815) );
  INV_X1 U904 ( .A(n813), .ZN(n814) );
  NOR2_X1 U905 ( .A1(G1976), .A2(G288), .ZN(n822) );
  NOR2_X1 U906 ( .A1(G1971), .A2(G303), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n822), .A2(n816), .ZN(n1036) );
  INV_X1 U908 ( .A(KEYINPUT33), .ZN(n820) );
  AND2_X1 U909 ( .A1(n1036), .A2(n820), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G1976), .A2(G288), .ZN(n1035) );
  INV_X1 U911 ( .A(n836), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n1035), .A2(n818), .ZN(n819) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(KEYINPUT33), .ZN(n823) );
  OR2_X1 U915 ( .A1(n836), .A2(n823), .ZN(n824) );
  NAND2_X1 U916 ( .A1(n825), .A2(n824), .ZN(n827) );
  XOR2_X1 U917 ( .A(G1981), .B(G305), .Z(n1024) );
  NOR2_X1 U918 ( .A1(G2090), .A2(G303), .ZN(n828) );
  NAND2_X1 U919 ( .A1(G8), .A2(n828), .ZN(n831) );
  BUF_X1 U920 ( .A(n829), .Z(n830) );
  NAND2_X1 U921 ( .A1(n831), .A2(n830), .ZN(n832) );
  NOR2_X1 U922 ( .A1(G1981), .A2(G305), .ZN(n834) );
  XOR2_X1 U923 ( .A(n834), .B(KEYINPUT24), .Z(n835) );
  NAND2_X1 U924 ( .A1(n837), .A2(n606), .ZN(n838) );
  NOR2_X1 U925 ( .A1(n839), .A2(n840), .ZN(n880) );
  XNOR2_X1 U926 ( .A(KEYINPUT37), .B(G2067), .ZN(n878) );
  NAND2_X1 U927 ( .A1(n938), .A2(G140), .ZN(n841) );
  XOR2_X1 U928 ( .A(KEYINPUT87), .B(n841), .Z(n843) );
  NAND2_X1 U929 ( .A1(n939), .A2(G104), .ZN(n842) );
  NAND2_X1 U930 ( .A1(n843), .A2(n842), .ZN(n844) );
  XNOR2_X1 U931 ( .A(KEYINPUT34), .B(n844), .ZN(n849) );
  NAND2_X1 U932 ( .A1(G128), .A2(n942), .ZN(n846) );
  NAND2_X1 U933 ( .A1(G116), .A2(n943), .ZN(n845) );
  NAND2_X1 U934 ( .A1(n846), .A2(n845), .ZN(n847) );
  XOR2_X1 U935 ( .A(KEYINPUT35), .B(n847), .Z(n848) );
  NOR2_X1 U936 ( .A1(n849), .A2(n848), .ZN(n850) );
  XNOR2_X1 U937 ( .A(KEYINPUT36), .B(n850), .ZN(n932) );
  NOR2_X1 U938 ( .A1(n878), .A2(n932), .ZN(n1015) );
  NAND2_X1 U939 ( .A1(n880), .A2(n1015), .ZN(n877) );
  NAND2_X1 U940 ( .A1(G119), .A2(n942), .ZN(n852) );
  NAND2_X1 U941 ( .A1(G131), .A2(n938), .ZN(n851) );
  NAND2_X1 U942 ( .A1(n852), .A2(n851), .ZN(n856) );
  NAND2_X1 U943 ( .A1(G107), .A2(n943), .ZN(n854) );
  NAND2_X1 U944 ( .A1(G95), .A2(n939), .ZN(n853) );
  NAND2_X1 U945 ( .A1(n854), .A2(n853), .ZN(n855) );
  OR2_X1 U946 ( .A1(n856), .A2(n855), .ZN(n929) );
  NAND2_X1 U947 ( .A1(G1991), .A2(n929), .ZN(n867) );
  NAND2_X1 U948 ( .A1(G129), .A2(n942), .ZN(n858) );
  NAND2_X1 U949 ( .A1(G141), .A2(n938), .ZN(n857) );
  NAND2_X1 U950 ( .A1(n858), .A2(n857), .ZN(n863) );
  XOR2_X1 U951 ( .A(KEYINPUT38), .B(KEYINPUT89), .Z(n860) );
  NAND2_X1 U952 ( .A1(G105), .A2(n939), .ZN(n859) );
  XNOR2_X1 U953 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U954 ( .A(KEYINPUT88), .B(n861), .Z(n862) );
  NOR2_X1 U955 ( .A1(n863), .A2(n862), .ZN(n865) );
  NAND2_X1 U956 ( .A1(n943), .A2(G117), .ZN(n864) );
  NAND2_X1 U957 ( .A1(n865), .A2(n864), .ZN(n934) );
  NAND2_X1 U958 ( .A1(G1996), .A2(n934), .ZN(n866) );
  NAND2_X1 U959 ( .A1(n867), .A2(n866), .ZN(n1003) );
  NAND2_X1 U960 ( .A1(n880), .A2(n1003), .ZN(n870) );
  XNOR2_X1 U961 ( .A(G1986), .B(G290), .ZN(n1032) );
  NAND2_X1 U962 ( .A1(n880), .A2(n1032), .ZN(n869) );
  NOR2_X1 U963 ( .A1(G1996), .A2(n934), .ZN(n1008) );
  INV_X1 U964 ( .A(n870), .ZN(n873) );
  NOR2_X1 U965 ( .A1(G1986), .A2(G290), .ZN(n871) );
  NOR2_X1 U966 ( .A1(G1991), .A2(n929), .ZN(n1004) );
  NOR2_X1 U967 ( .A1(n871), .A2(n1004), .ZN(n872) );
  NOR2_X1 U968 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U969 ( .A1(n1008), .A2(n874), .ZN(n875) );
  XNOR2_X1 U970 ( .A(KEYINPUT39), .B(n875), .ZN(n876) );
  NAND2_X1 U971 ( .A1(n877), .A2(n876), .ZN(n879) );
  NAND2_X1 U972 ( .A1(n878), .A2(n932), .ZN(n1012) );
  NAND2_X1 U973 ( .A1(n879), .A2(n1012), .ZN(n881) );
  NAND2_X1 U974 ( .A1(n881), .A2(n880), .ZN(n882) );
  NAND2_X1 U975 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U976 ( .A(n884), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U977 ( .A1(G2106), .A2(n885), .ZN(G217) );
  AND2_X1 U978 ( .A1(G15), .A2(G2), .ZN(n886) );
  NAND2_X1 U979 ( .A1(G661), .A2(n886), .ZN(G259) );
  NAND2_X1 U980 ( .A1(G3), .A2(G1), .ZN(n888) );
  NAND2_X1 U981 ( .A1(n888), .A2(n887), .ZN(n889) );
  XOR2_X1 U982 ( .A(KEYINPUT107), .B(n889), .Z(G188) );
  XOR2_X1 U983 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U985 ( .A(G96), .ZN(G221) );
  INV_X1 U986 ( .A(G69), .ZN(G235) );
  NOR2_X1 U987 ( .A1(n891), .A2(n890), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n892), .B(KEYINPUT109), .ZN(G261) );
  INV_X1 U989 ( .A(G261), .ZN(G325) );
  INV_X1 U990 ( .A(n893), .ZN(G319) );
  XOR2_X1 U991 ( .A(G2096), .B(KEYINPUT43), .Z(n895) );
  XNOR2_X1 U992 ( .A(G2072), .B(G2678), .ZN(n894) );
  XNOR2_X1 U993 ( .A(n895), .B(n894), .ZN(n896) );
  XOR2_X1 U994 ( .A(n896), .B(KEYINPUT110), .Z(n898) );
  XNOR2_X1 U995 ( .A(G2067), .B(G2090), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n902) );
  XOR2_X1 U997 ( .A(KEYINPUT42), .B(G2100), .Z(n900) );
  XNOR2_X1 U998 ( .A(G2084), .B(G2078), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(G227) );
  XOR2_X1 U1001 ( .A(G1971), .B(G1961), .Z(n904) );
  XNOR2_X1 U1002 ( .A(G1986), .B(G1966), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n905) );
  XOR2_X1 U1004 ( .A(n905), .B(G2474), .Z(n907) );
  XNOR2_X1 U1005 ( .A(G1981), .B(G1956), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n911) );
  XOR2_X1 U1007 ( .A(KEYINPUT41), .B(G1976), .Z(n909) );
  XNOR2_X1 U1008 ( .A(G1996), .B(G1991), .ZN(n908) );
  XNOR2_X1 U1009 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(G229) );
  NAND2_X1 U1011 ( .A1(n942), .A2(G124), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n912), .B(KEYINPUT44), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(G112), .A2(n943), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n918) );
  NAND2_X1 U1015 ( .A1(G136), .A2(n938), .ZN(n916) );
  NAND2_X1 U1016 ( .A1(G100), .A2(n939), .ZN(n915) );
  NAND2_X1 U1017 ( .A1(n916), .A2(n915), .ZN(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(G162) );
  NAND2_X1 U1019 ( .A1(G130), .A2(n942), .ZN(n920) );
  NAND2_X1 U1020 ( .A1(G118), .A2(n943), .ZN(n919) );
  NAND2_X1 U1021 ( .A1(n920), .A2(n919), .ZN(n925) );
  NAND2_X1 U1022 ( .A1(G142), .A2(n938), .ZN(n922) );
  NAND2_X1 U1023 ( .A1(G106), .A2(n939), .ZN(n921) );
  NAND2_X1 U1024 ( .A1(n922), .A2(n921), .ZN(n923) );
  XOR2_X1 U1025 ( .A(KEYINPUT45), .B(n923), .Z(n924) );
  NOR2_X1 U1026 ( .A1(n925), .A2(n924), .ZN(n937) );
  XOR2_X1 U1027 ( .A(KEYINPUT48), .B(KEYINPUT111), .Z(n927) );
  XNOR2_X1 U1028 ( .A(G160), .B(KEYINPUT46), .ZN(n926) );
  XNOR2_X1 U1029 ( .A(n927), .B(n926), .ZN(n928) );
  XNOR2_X1 U1030 ( .A(n1002), .B(n928), .ZN(n931) );
  XNOR2_X1 U1031 ( .A(n929), .B(G162), .ZN(n930) );
  XNOR2_X1 U1032 ( .A(n931), .B(n930), .ZN(n933) );
  XNOR2_X1 U1033 ( .A(n933), .B(n932), .ZN(n935) );
  XNOR2_X1 U1034 ( .A(n935), .B(n934), .ZN(n936) );
  XNOR2_X1 U1035 ( .A(n937), .B(n936), .ZN(n950) );
  NAND2_X1 U1036 ( .A1(G139), .A2(n938), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(G103), .A2(n939), .ZN(n940) );
  NAND2_X1 U1038 ( .A1(n941), .A2(n940), .ZN(n948) );
  NAND2_X1 U1039 ( .A1(G127), .A2(n942), .ZN(n945) );
  NAND2_X1 U1040 ( .A1(G115), .A2(n943), .ZN(n944) );
  NAND2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1042 ( .A(KEYINPUT47), .B(n946), .Z(n947) );
  NOR2_X1 U1043 ( .A1(n948), .A2(n947), .ZN(n997) );
  XNOR2_X1 U1044 ( .A(G164), .B(n997), .ZN(n949) );
  XNOR2_X1 U1045 ( .A(n950), .B(n949), .ZN(n951) );
  NOR2_X1 U1046 ( .A1(G37), .A2(n951), .ZN(G395) );
  INV_X1 U1047 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U1048 ( .A(n952), .B(KEYINPUT112), .ZN(n954) );
  XNOR2_X1 U1049 ( .A(n1039), .B(G286), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(n954), .B(n953), .ZN(n955) );
  XNOR2_X1 U1051 ( .A(n955), .B(G301), .ZN(n956) );
  NOR2_X1 U1052 ( .A1(G37), .A2(n956), .ZN(G397) );
  XOR2_X1 U1053 ( .A(G2451), .B(G2430), .Z(n958) );
  XNOR2_X1 U1054 ( .A(G2438), .B(G2443), .ZN(n957) );
  XNOR2_X1 U1055 ( .A(n958), .B(n957), .ZN(n964) );
  XOR2_X1 U1056 ( .A(G2435), .B(G2454), .Z(n960) );
  XNOR2_X1 U1057 ( .A(G1348), .B(G1341), .ZN(n959) );
  XNOR2_X1 U1058 ( .A(n960), .B(n959), .ZN(n962) );
  XOR2_X1 U1059 ( .A(G2446), .B(G2427), .Z(n961) );
  XNOR2_X1 U1060 ( .A(n962), .B(n961), .ZN(n963) );
  XOR2_X1 U1061 ( .A(n964), .B(n963), .Z(n965) );
  NAND2_X1 U1062 ( .A1(G14), .A2(n965), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(G319), .A2(n972), .ZN(n969) );
  NOR2_X1 U1064 ( .A1(G227), .A2(G229), .ZN(n966) );
  XOR2_X1 U1065 ( .A(KEYINPUT113), .B(n966), .Z(n967) );
  XNOR2_X1 U1066 ( .A(n967), .B(KEYINPUT49), .ZN(n968) );
  NOR2_X1 U1067 ( .A1(n969), .A2(n968), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(G395), .A2(G397), .ZN(n970) );
  NAND2_X1 U1069 ( .A1(n971), .A2(n970), .ZN(G225) );
  INV_X1 U1070 ( .A(G225), .ZN(G308) );
  INV_X1 U1071 ( .A(G57), .ZN(G237) );
  INV_X1 U1072 ( .A(n972), .ZN(G401) );
  XOR2_X1 U1073 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n988) );
  XNOR2_X1 U1074 ( .A(G1991), .B(G25), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(G32), .B(n973), .ZN(n978) );
  XNOR2_X1 U1076 ( .A(G2067), .B(G26), .ZN(n976) );
  XNOR2_X1 U1077 ( .A(n974), .B(G27), .ZN(n975) );
  NOR2_X1 U1078 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1079 ( .A1(n978), .A2(n977), .ZN(n982) );
  XOR2_X1 U1080 ( .A(KEYINPUT116), .B(n979), .Z(n980) );
  XNOR2_X1 U1081 ( .A(G33), .B(n980), .ZN(n981) );
  NOR2_X1 U1082 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1083 ( .A(KEYINPUT117), .B(n983), .ZN(n984) );
  NOR2_X1 U1084 ( .A1(n985), .A2(n984), .ZN(n986) );
  NAND2_X1 U1085 ( .A1(n986), .A2(G28), .ZN(n987) );
  XNOR2_X1 U1086 ( .A(n988), .B(n987), .ZN(n990) );
  XNOR2_X1 U1087 ( .A(G35), .B(G2090), .ZN(n989) );
  NOR2_X1 U1088 ( .A1(n990), .A2(n989), .ZN(n993) );
  XOR2_X1 U1089 ( .A(G2084), .B(KEYINPUT54), .Z(n991) );
  XNOR2_X1 U1090 ( .A(G34), .B(n991), .ZN(n992) );
  NAND2_X1 U1091 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1092 ( .A(KEYINPUT119), .B(n994), .ZN(n995) );
  NOR2_X1 U1093 ( .A1(G29), .A2(n995), .ZN(n996) );
  XNOR2_X1 U1094 ( .A(n996), .B(KEYINPUT55), .ZN(n1023) );
  XOR2_X1 U1095 ( .A(G2072), .B(n997), .Z(n999) );
  XOR2_X1 U1096 ( .A(G164), .B(G2078), .Z(n998) );
  NOR2_X1 U1097 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1000), .Z(n1018) );
  XOR2_X1 U1099 ( .A(G160), .B(G2084), .Z(n1001) );
  NOR2_X1 U1100 ( .A1(n1002), .A2(n1001), .ZN(n1006) );
  NOR2_X1 U1101 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1102 ( .A1(n1006), .A2(n1005), .ZN(n1011) );
  XOR2_X1 U1103 ( .A(G2090), .B(G162), .Z(n1007) );
  NOR2_X1 U1104 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1105 ( .A(n1009), .B(KEYINPUT51), .ZN(n1010) );
  NOR2_X1 U1106 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  NAND2_X1 U1107 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NOR2_X1 U1108 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1109 ( .A(KEYINPUT114), .B(n1016), .Z(n1017) );
  NOR2_X1 U1110 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1111 ( .A(n1019), .B(KEYINPUT52), .ZN(n1020) );
  XNOR2_X1 U1112 ( .A(n1020), .B(KEYINPUT115), .ZN(n1021) );
  NAND2_X1 U1113 ( .A1(G29), .A2(n1021), .ZN(n1022) );
  NAND2_X1 U1114 ( .A1(n1023), .A2(n1022), .ZN(n1080) );
  XOR2_X1 U1115 ( .A(G16), .B(KEYINPUT56), .Z(n1048) );
  XNOR2_X1 U1116 ( .A(G1966), .B(G168), .ZN(n1025) );
  NAND2_X1 U1117 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  XNOR2_X1 U1118 ( .A(n1026), .B(KEYINPUT120), .ZN(n1027) );
  XNOR2_X1 U1119 ( .A(KEYINPUT57), .B(n1027), .ZN(n1034) );
  XNOR2_X1 U1120 ( .A(n1028), .B(G1341), .ZN(n1030) );
  NAND2_X1 U1121 ( .A1(G1971), .A2(G303), .ZN(n1029) );
  NAND2_X1 U1122 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  NOR2_X1 U1123 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NAND2_X1 U1124 ( .A1(n1034), .A2(n1033), .ZN(n1046) );
  NAND2_X1 U1125 ( .A1(n1036), .A2(n1035), .ZN(n1038) );
  XNOR2_X1 U1126 ( .A(G1956), .B(G299), .ZN(n1037) );
  NOR2_X1 U1127 ( .A1(n1038), .A2(n1037), .ZN(n1044) );
  XNOR2_X1 U1128 ( .A(G301), .B(G1961), .ZN(n1041) );
  XNOR2_X1 U1129 ( .A(n1039), .B(G1348), .ZN(n1040) );
  NOR2_X1 U1130 ( .A1(n1041), .A2(n1040), .ZN(n1042) );
  XOR2_X1 U1131 ( .A(KEYINPUT121), .B(n1042), .Z(n1043) );
  NAND2_X1 U1132 ( .A1(n1044), .A2(n1043), .ZN(n1045) );
  NOR2_X1 U1133 ( .A1(n1046), .A2(n1045), .ZN(n1047) );
  NOR2_X1 U1134 ( .A1(n1048), .A2(n1047), .ZN(n1077) );
  XOR2_X1 U1135 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n1055) );
  XNOR2_X1 U1136 ( .A(G1971), .B(G22), .ZN(n1050) );
  XNOR2_X1 U1137 ( .A(G23), .B(G1976), .ZN(n1049) );
  NOR2_X1 U1138 ( .A1(n1050), .A2(n1049), .ZN(n1053) );
  XNOR2_X1 U1139 ( .A(G1986), .B(KEYINPUT125), .ZN(n1051) );
  XNOR2_X1 U1140 ( .A(n1051), .B(G24), .ZN(n1052) );
  NAND2_X1 U1141 ( .A1(n1053), .A2(n1052), .ZN(n1054) );
  XNOR2_X1 U1142 ( .A(n1055), .B(n1054), .ZN(n1059) );
  XNOR2_X1 U1143 ( .A(G1966), .B(G21), .ZN(n1057) );
  XNOR2_X1 U1144 ( .A(G5), .B(G1961), .ZN(n1056) );
  NOR2_X1 U1145 ( .A1(n1057), .A2(n1056), .ZN(n1058) );
  NAND2_X1 U1146 ( .A1(n1059), .A2(n1058), .ZN(n1073) );
  XOR2_X1 U1147 ( .A(G1956), .B(G20), .Z(n1062) );
  XNOR2_X1 U1148 ( .A(n1060), .B(G19), .ZN(n1061) );
  NAND2_X1 U1149 ( .A1(n1062), .A2(n1061), .ZN(n1064) );
  XNOR2_X1 U1150 ( .A(G6), .B(G1981), .ZN(n1063) );
  NOR2_X1 U1151 ( .A1(n1064), .A2(n1063), .ZN(n1065) );
  XNOR2_X1 U1152 ( .A(KEYINPUT122), .B(n1065), .ZN(n1069) );
  XOR2_X1 U1153 ( .A(KEYINPUT123), .B(G4), .Z(n1067) );
  XNOR2_X1 U1154 ( .A(G1348), .B(KEYINPUT59), .ZN(n1066) );
  XNOR2_X1 U1155 ( .A(n1067), .B(n1066), .ZN(n1068) );
  NAND2_X1 U1156 ( .A1(n1069), .A2(n1068), .ZN(n1070) );
  XNOR2_X1 U1157 ( .A(n1070), .B(KEYINPUT124), .ZN(n1071) );
  XNOR2_X1 U1158 ( .A(n1071), .B(KEYINPUT60), .ZN(n1072) );
  NOR2_X1 U1159 ( .A1(n1073), .A2(n1072), .ZN(n1074) );
  XOR2_X1 U1160 ( .A(KEYINPUT61), .B(n1074), .Z(n1075) );
  NOR2_X1 U1161 ( .A1(G16), .A2(n1075), .ZN(n1076) );
  NOR2_X1 U1162 ( .A1(n1077), .A2(n1076), .ZN(n1078) );
  XNOR2_X1 U1163 ( .A(KEYINPUT127), .B(n1078), .ZN(n1079) );
  NOR2_X1 U1164 ( .A1(n1080), .A2(n1079), .ZN(n1081) );
  NAND2_X1 U1165 ( .A1(n1081), .A2(G11), .ZN(n1082) );
  XOR2_X1 U1166 ( .A(KEYINPUT62), .B(n1082), .Z(G311) );
  INV_X1 U1167 ( .A(G311), .ZN(G150) );
endmodule

