//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n242, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n258, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1034, new_n1035,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1074, new_n1075, new_n1076, new_n1077, new_n1078,
    new_n1079, new_n1080, new_n1081, new_n1082, new_n1083, new_n1084,
    new_n1085, new_n1086, new_n1087, new_n1088, new_n1089, new_n1090,
    new_n1091, new_n1092, new_n1093, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1118, new_n1119, new_n1120, new_n1121,
    new_n1122, new_n1123, new_n1124, new_n1125, new_n1126, new_n1127,
    new_n1128, new_n1129, new_n1130, new_n1131, new_n1132, new_n1133,
    new_n1134, new_n1135, new_n1136, new_n1137, new_n1138, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1201, new_n1202;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0008(.A(KEYINPUT65), .ZN(new_n209));
  INV_X1    g0009(.A(G1), .ZN(new_n210));
  INV_X1    g0010(.A(G20), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  OAI21_X1  g0013(.A(new_n209), .B1(new_n213), .B2(G13), .ZN(new_n214));
  INV_X1    g0014(.A(G13), .ZN(new_n215));
  NAND3_X1  g0015(.A1(new_n212), .A2(KEYINPUT65), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT66), .B(KEYINPUT0), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n218), .B(new_n219), .ZN(new_n220));
  XOR2_X1   g0020(.A(KEYINPUT68), .B(G244), .Z(new_n221));
  AOI22_X1  g0021(.A1(new_n221), .A2(G77), .B1(G116), .B2(G270), .ZN(new_n222));
  INV_X1    g0022(.A(G50), .ZN(new_n223));
  INV_X1    g0023(.A(G226), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G87), .ZN(new_n228));
  INV_X1    g0028(.A(G250), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n202), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g0032(.A1(G68), .A2(G238), .ZN(new_n233));
  NOR4_X1   g0033(.A1(new_n227), .A2(new_n230), .A3(new_n232), .A4(new_n233), .ZN(new_n234));
  NAND2_X1  g0034(.A1(G97), .A2(G257), .ZN(new_n235));
  AOI21_X1  g0035(.A(new_n212), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(KEYINPUT1), .ZN(new_n237));
  AND2_X1   g0037(.A1(G1), .A2(G13), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n238), .A2(G20), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n206), .A2(G50), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(new_n241));
  OAI22_X1  g0041(.A1(new_n236), .A2(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  AOI211_X1 g0042(.A(new_n220), .B(new_n242), .C1(new_n237), .C2(new_n236), .ZN(G361));
  XNOR2_X1  g0043(.A(G238), .B(G244), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(new_n231), .ZN(new_n245));
  XOR2_X1   g0045(.A(KEYINPUT2), .B(G226), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G250), .B(G257), .Z(new_n248));
  XNOR2_X1  g0048(.A(G264), .B(G270), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G358));
  XOR2_X1   g0051(.A(G68), .B(G77), .Z(new_n252));
  XOR2_X1   g0052(.A(G50), .B(G58), .Z(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n254), .B(KEYINPUT69), .ZN(new_n255));
  XOR2_X1   g0055(.A(G87), .B(G97), .Z(new_n256));
  XNOR2_X1  g0056(.A(G107), .B(G116), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n256), .B(new_n257), .ZN(new_n258));
  XNOR2_X1  g0058(.A(new_n255), .B(new_n258), .ZN(G351));
  NAND3_X1  g0059(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G1), .A2(G13), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n210), .A2(G20), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  XOR2_X1   g0065(.A(KEYINPUT8), .B(G58), .Z(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n264), .A2(new_n215), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n267), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT80), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n269), .B(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT16), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n211), .A2(KEYINPUT7), .ZN(new_n273));
  INV_X1    g0073(.A(G33), .ZN(new_n274));
  NOR2_X1   g0074(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n275));
  AOI21_X1  g0075(.A(new_n273), .B1(new_n275), .B2(KEYINPUT78), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n274), .A2(KEYINPUT3), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(G33), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT78), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n277), .A2(new_n279), .A3(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n276), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT7), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n283), .B1(new_n284), .B2(G20), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n203), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G58), .A2(G68), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT77), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(KEYINPUT77), .A2(G58), .A3(G68), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n204), .A2(new_n289), .A3(new_n205), .A4(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G20), .ZN(new_n292));
  NOR2_X1   g0092(.A1(G20), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(G159), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n272), .B1(new_n286), .B2(new_n295), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n291), .A2(G20), .B1(G159), .B2(new_n293), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n277), .A2(new_n279), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(new_n211), .ZN(new_n299));
  INV_X1    g0099(.A(new_n273), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n299), .A2(new_n283), .B1(new_n298), .B2(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(KEYINPUT16), .B(new_n297), .C1(new_n301), .C2(new_n203), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n296), .A2(new_n302), .A3(new_n262), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT79), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n296), .A2(new_n302), .A3(KEYINPUT79), .A4(new_n262), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n271), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n224), .A2(G1698), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n284), .B(new_n308), .C1(G223), .C2(G1698), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G41), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n238), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G41), .ZN(new_n316));
  INV_X1    g0116(.A(G45), .ZN(new_n317));
  AOI21_X1  g0117(.A(G1), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n238), .A2(KEYINPUT70), .A3(new_n312), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(G232), .ZN(new_n323));
  INV_X1    g0123(.A(new_n321), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT70), .B1(new_n238), .B2(new_n312), .ZN(new_n325));
  OAI211_X1 g0125(.A(G274), .B(new_n318), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n315), .A2(new_n323), .A3(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(G190), .ZN(new_n328));
  OR2_X1    g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n327), .A2(G200), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n307), .A2(new_n329), .A3(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT17), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  AOI211_X1 g0134(.A(new_n271), .B(new_n330), .C1(new_n305), .C2(new_n306), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n335), .A2(KEYINPUT17), .A3(new_n329), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT81), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(new_n271), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n299), .A2(new_n283), .B1(new_n276), .B2(new_n281), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n297), .B1(new_n341), .B2(new_n203), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n263), .B1(new_n342), .B2(new_n272), .ZN(new_n343));
  AOI21_X1  g0143(.A(KEYINPUT79), .B1(new_n343), .B2(new_n302), .ZN(new_n344));
  INV_X1    g0144(.A(new_n306), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n340), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n327), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n348), .B1(G169), .B2(new_n327), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT18), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n351), .B(new_n352), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n334), .A2(new_n336), .A3(KEYINPUT81), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n339), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n211), .A2(G33), .ZN(new_n357));
  XOR2_X1   g0157(.A(new_n357), .B(KEYINPUT72), .Z(new_n358));
  AOI22_X1  g0158(.A1(new_n358), .A2(new_n266), .B1(G150), .B2(new_n293), .ZN(new_n359));
  OAI21_X1  g0159(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n262), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n263), .A2(G50), .A3(new_n264), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n268), .A2(new_n223), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(G1698), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n284), .A2(G222), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT71), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n284), .A2(G223), .A3(G1698), .ZN(new_n369));
  INV_X1    g0169(.A(G77), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n368), .B(new_n369), .C1(new_n370), .C2(new_n284), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n314), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n322), .A2(G226), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n326), .A3(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(new_n374), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n365), .B1(new_n375), .B2(G169), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(new_n347), .B2(new_n375), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n374), .A2(G200), .ZN(new_n378));
  NOR2_X1   g0178(.A1(new_n378), .A2(KEYINPUT73), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT73), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n374), .B2(G200), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT10), .ZN(new_n383));
  INV_X1    g0183(.A(new_n365), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(KEYINPUT9), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT9), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n375), .A2(G190), .B1(new_n365), .B2(new_n386), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n382), .A2(new_n383), .A3(new_n385), .A4(new_n387), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n387), .B(new_n385), .C1(new_n379), .C2(new_n381), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT10), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n377), .B1(new_n388), .B2(new_n390), .ZN(new_n391));
  AOI22_X1  g0191(.A1(new_n266), .A2(new_n293), .B1(G20), .B2(G77), .ZN(new_n392));
  XOR2_X1   g0192(.A(KEYINPUT15), .B(G87), .Z(new_n393));
  INV_X1    g0193(.A(new_n393), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n392), .B1(new_n357), .B2(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n395), .A2(new_n262), .B1(new_n370), .B2(new_n268), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n370), .B2(new_n265), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n322), .A2(new_n221), .ZN(new_n398));
  NOR2_X1   g0198(.A1(G232), .A2(G1698), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n366), .A2(G238), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n284), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n314), .C1(G107), .C2(new_n284), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n398), .A2(new_n326), .A3(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n403), .A2(G179), .ZN(new_n404));
  INV_X1    g0204(.A(G169), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n397), .A2(new_n404), .A3(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n356), .A2(new_n391), .A3(new_n407), .ZN(new_n408));
  AOI22_X1  g0208(.A1(new_n358), .A2(G77), .B1(G20), .B2(new_n203), .ZN(new_n409));
  OR2_X1    g0209(.A1(new_n409), .A2(KEYINPUT74), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n293), .A2(G50), .ZN(new_n411));
  XOR2_X1   g0211(.A(new_n411), .B(KEYINPUT75), .Z(new_n412));
  NAND2_X1  g0212(.A1(new_n409), .A2(KEYINPUT74), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n410), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n262), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n415), .A2(KEYINPUT11), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT11), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n414), .A2(new_n417), .A3(new_n262), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n268), .ZN(new_n420));
  NOR3_X1   g0220(.A1(new_n420), .A2(KEYINPUT12), .A3(G68), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT12), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n268), .B2(new_n203), .ZN(new_n423));
  OAI22_X1  g0223(.A1(new_n421), .A2(new_n423), .B1(new_n203), .B2(new_n265), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT76), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n231), .A2(G1698), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(G226), .B2(G1698), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n298), .ZN(new_n431));
  INV_X1    g0231(.A(G97), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n274), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n314), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n318), .ZN(new_n435));
  OAI211_X1 g0235(.A(G238), .B(new_n435), .C1(new_n324), .C2(new_n325), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n326), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(KEYINPUT13), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT13), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n434), .A2(new_n326), .A3(new_n436), .A4(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n428), .B1(new_n441), .B2(G169), .ZN(new_n442));
  AOI211_X1 g0242(.A(KEYINPUT14), .B(new_n405), .C1(new_n438), .C2(new_n440), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(new_n441), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(G179), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n427), .B1(new_n444), .B2(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n441), .A2(G169), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT14), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n441), .A2(new_n428), .A3(G169), .ZN(new_n450));
  AND4_X1   g0250(.A1(new_n427), .A2(new_n449), .A3(new_n446), .A4(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n426), .B1(new_n447), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n445), .A2(G190), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n441), .A2(G200), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n419), .A2(new_n425), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n397), .B1(G200), .B2(new_n403), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n328), .B2(new_n403), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n408), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n210), .A2(G45), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT5), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(G41), .ZN(new_n462));
  OAI21_X1  g0262(.A(KEYINPUT82), .B1(new_n461), .B2(G41), .ZN(new_n463));
  OR3_X1    g0263(.A1(new_n461), .A2(KEYINPUT82), .A3(G41), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n320), .A2(new_n321), .ZN(new_n466));
  AND2_X1   g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n277), .A2(new_n279), .A3(G250), .A4(new_n366), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(KEYINPUT88), .ZN(new_n469));
  XOR2_X1   g0269(.A(KEYINPUT89), .B(G294), .Z(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G33), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT88), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n284), .A2(new_n472), .A3(G250), .A4(new_n366), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n284), .A2(G257), .A3(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n469), .A2(new_n471), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  AOI22_X1  g0275(.A1(new_n467), .A2(G264), .B1(new_n475), .B2(new_n314), .ZN(new_n476));
  AND3_X1   g0276(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n477));
  INV_X1    g0277(.A(G274), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n320), .B2(new_n321), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n476), .A2(new_n328), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n475), .A2(new_n314), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n465), .A2(new_n466), .A3(G264), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n482), .A2(new_n480), .A3(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(G200), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n210), .A2(G33), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n420), .A2(new_n263), .A3(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G107), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT23), .B1(new_n211), .B2(G107), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT23), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n493), .A2(new_n225), .A3(G20), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n211), .A2(G33), .A3(G116), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT86), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n492), .A2(new_n494), .A3(new_n495), .A4(KEYINPUT86), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  AND4_X1   g0301(.A1(new_n211), .A2(new_n277), .A3(new_n279), .A4(G87), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT85), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n284), .A2(new_n503), .A3(new_n211), .A4(G87), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n505), .A2(KEYINPUT22), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT24), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n500), .B(KEYINPUT24), .C1(new_n504), .C2(new_n506), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n509), .A2(new_n262), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n420), .A2(G107), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n512), .B1(KEYINPUT87), .B2(KEYINPUT25), .ZN(new_n513));
  NAND2_X1  g0313(.A1(KEYINPUT87), .A2(KEYINPUT25), .ZN(new_n514));
  MUX2_X1   g0314(.A(new_n512), .B(new_n513), .S(new_n514), .Z(new_n515));
  NAND4_X1  g0315(.A1(new_n487), .A2(new_n491), .A3(new_n511), .A4(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n341), .A2(new_n225), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n293), .A2(G77), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT6), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n432), .A2(new_n225), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G97), .A2(G107), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n225), .A2(KEYINPUT6), .A3(G97), .ZN(new_n523));
  AND2_X1   g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n518), .B1(new_n524), .B2(new_n211), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n262), .B1(new_n517), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n490), .A2(G97), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n268), .A2(new_n432), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n284), .A2(G244), .A3(new_n366), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT4), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(G33), .A2(G283), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n366), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n532), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n314), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n467), .A2(G257), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n538), .A3(new_n480), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n539), .A2(new_n347), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n536), .A2(new_n314), .B1(new_n479), .B2(new_n477), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n405), .B1(new_n541), .B2(new_n538), .ZN(new_n542));
  OAI21_X1  g0342(.A(new_n529), .B1(new_n540), .B2(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n539), .A2(G200), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n541), .A2(G190), .A3(new_n538), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n465), .A2(new_n466), .A3(G270), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n226), .A2(G1698), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(G257), .B2(G1698), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n313), .B1(new_n550), .B2(new_n284), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G303), .B2(new_n284), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n480), .A2(new_n548), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G200), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n420), .A2(G116), .A3(new_n263), .A4(new_n488), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n268), .A2(new_n556), .ZN(new_n557));
  AOI22_X1  g0357(.A1(new_n260), .A2(new_n261), .B1(G20), .B2(new_n556), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n534), .B(new_n211), .C1(G33), .C2(new_n432), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n558), .A2(KEYINPUT20), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT20), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  OAI211_X1 g0361(.A(new_n555), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n554), .B(new_n563), .C1(new_n328), .C2(new_n553), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n516), .A2(new_n543), .A3(new_n547), .A4(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n511), .A2(new_n491), .A3(new_n515), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n484), .A2(new_n405), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n476), .A2(new_n347), .A3(new_n480), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n420), .A2(new_n393), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n284), .A2(new_n211), .A3(G68), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n357), .A2(new_n432), .ZN(new_n572));
  NOR3_X1   g0372(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n573));
  XNOR2_X1  g0373(.A(new_n573), .B(KEYINPUT83), .ZN(new_n574));
  AOI21_X1  g0374(.A(G20), .B1(new_n433), .B2(KEYINPUT19), .ZN(new_n575));
  OAI221_X1 g0375(.A(new_n571), .B1(KEYINPUT19), .B2(new_n572), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n570), .B1(new_n576), .B2(new_n262), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n393), .B(KEYINPUT84), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n490), .ZN(new_n579));
  OR2_X1    g0379(.A1(new_n366), .A2(G244), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n284), .B(new_n580), .C1(G238), .C2(G1698), .ZN(new_n581));
  NAND2_X1  g0381(.A1(G33), .A2(G116), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n314), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n460), .A2(new_n229), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n210), .A2(new_n478), .A3(G45), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n466), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n577), .A2(new_n579), .B1(new_n405), .B2(new_n588), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n584), .A2(new_n587), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n347), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n485), .B1(new_n584), .B2(new_n587), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(G190), .B2(new_n590), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n489), .A2(new_n228), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n570), .B(new_n594), .C1(new_n576), .C2(new_n262), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n589), .A2(new_n591), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n553), .A2(G169), .A3(new_n562), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n553), .A2(new_n347), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n562), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n553), .A2(KEYINPUT21), .A3(new_n562), .A4(G169), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n599), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n569), .A2(new_n596), .A3(new_n603), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n565), .A2(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n459), .A2(new_n605), .ZN(G372));
  AND2_X1   g0406(.A1(new_n589), .A2(new_n591), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT91), .ZN(new_n608));
  XNOR2_X1  g0408(.A(new_n595), .B(new_n608), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n592), .A2(KEYINPUT90), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n590), .A2(G190), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n592), .A2(KEYINPUT90), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n607), .B1(new_n609), .B2(new_n614), .ZN(new_n615));
  AND2_X1   g0415(.A1(new_n547), .A2(new_n543), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n569), .A2(new_n603), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n615), .A2(new_n616), .A3(new_n516), .A4(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT26), .ZN(new_n619));
  INV_X1    g0419(.A(new_n543), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n615), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n589), .A2(new_n591), .ZN(new_n622));
  INV_X1    g0422(.A(new_n596), .ZN(new_n623));
  OAI21_X1  g0423(.A(KEYINPUT26), .B1(new_n623), .B2(new_n543), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n618), .A2(new_n621), .A3(new_n622), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n459), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n339), .A2(new_n354), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n449), .A2(new_n446), .A3(new_n450), .ZN(new_n628));
  XNOR2_X1  g0428(.A(new_n628), .B(KEYINPUT76), .ZN(new_n629));
  INV_X1    g0429(.A(new_n407), .ZN(new_n630));
  AOI22_X1  g0430(.A1(new_n629), .A2(new_n426), .B1(new_n630), .B2(new_n455), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n353), .B1(new_n627), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n388), .A2(new_n390), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n377), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n626), .A2(new_n634), .ZN(G369));
  NOR2_X1   g0435(.A1(new_n215), .A2(G20), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n636), .A2(new_n210), .ZN(new_n637));
  XOR2_X1   g0437(.A(new_n637), .B(KEYINPUT92), .Z(new_n638));
  OR2_X1    g0438(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(KEYINPUT27), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n639), .A2(G213), .A3(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n562), .ZN(new_n644));
  XNOR2_X1  g0444(.A(new_n603), .B(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(new_n564), .ZN(new_n646));
  XNOR2_X1  g0446(.A(new_n646), .B(KEYINPUT93), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(G330), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n566), .B1(new_n481), .B2(new_n486), .ZN(new_n649));
  AND2_X1   g0449(.A1(new_n566), .A2(new_n643), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n569), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  OR2_X1    g0451(.A1(new_n569), .A2(new_n643), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n648), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n603), .A2(new_n643), .ZN(new_n657));
  XNOR2_X1  g0457(.A(new_n657), .B(KEYINPUT94), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g0459(.A1(new_n659), .A2(new_n652), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n217), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n574), .A2(new_n556), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n663), .A2(new_n664), .A3(new_n210), .ZN(new_n665));
  INV_X1    g0465(.A(new_n240), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n665), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  XNOR2_X1  g0467(.A(KEYINPUT95), .B(KEYINPUT28), .ZN(new_n668));
  XNOR2_X1  g0468(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n623), .A2(KEYINPUT26), .A3(new_n543), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n615), .A2(new_n620), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n670), .B1(new_n671), .B2(KEYINPUT26), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n672), .A2(new_n622), .A3(new_n618), .ZN(new_n673));
  INV_X1    g0473(.A(new_n643), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n675), .A2(KEYINPUT29), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n625), .A2(new_n674), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT29), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n541), .A2(new_n590), .A3(new_n538), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n682), .A2(KEYINPUT30), .A3(new_n476), .A4(new_n600), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT30), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n600), .A2(new_n476), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n681), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n539), .A2(new_n347), .A3(new_n484), .A4(new_n553), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n683), .B(new_n686), .C1(new_n590), .C2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n688), .A2(new_n643), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(KEYINPUT31), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT31), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n688), .A2(new_n691), .A3(new_n643), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT96), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n694), .B1(new_n605), .B2(new_n674), .ZN(new_n695));
  NOR4_X1   g0495(.A1(new_n565), .A2(new_n604), .A3(KEYINPUT96), .A4(new_n643), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n693), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G330), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n680), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n669), .B1(new_n700), .B2(G1), .ZN(G364));
  XNOR2_X1  g0501(.A(new_n648), .B(KEYINPUT98), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n210), .B1(new_n636), .B2(G45), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n663), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n647), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT97), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI211_X1 g0508(.A(new_n702), .B(new_n708), .C1(new_n707), .C2(new_n706), .ZN(new_n709));
  INV_X1    g0509(.A(new_n705), .ZN(new_n710));
  NOR2_X1   g0510(.A1(G13), .A2(G33), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n711), .B(KEYINPUT100), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(new_n211), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n710), .B1(new_n646), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n261), .B1(G20), .B2(new_n405), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n211), .A2(new_n328), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n717), .A2(new_n347), .A3(G200), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n211), .A2(G190), .ZN(new_n719));
  NOR2_X1   g0519(.A1(G179), .A2(G200), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI22_X1  g0522(.A1(new_n718), .A2(G322), .B1(G329), .B2(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n347), .A2(new_n485), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n716), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(G326), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n723), .A2(new_n298), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n485), .A2(G179), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(new_n719), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n728), .B1(G283), .B2(new_n731), .ZN(new_n732));
  INV_X1    g0532(.A(new_n719), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n733), .A2(new_n347), .A3(G200), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n724), .A2(new_n719), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  XNOR2_X1  g0536(.A(KEYINPUT33), .B(G317), .ZN(new_n737));
  AOI22_X1  g0537(.A1(new_n734), .A2(G311), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n470), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n211), .B1(new_n720), .B2(G190), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n732), .B(new_n738), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n716), .A2(new_n729), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n741), .B1(G303), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(G87), .ZN(new_n745));
  INV_X1    g0545(.A(new_n734), .ZN(new_n746));
  OR2_X1    g0546(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n746), .A2(KEYINPUT101), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  OAI221_X1 g0549(.A(new_n745), .B1(new_n203), .B2(new_n735), .C1(new_n749), .C2(new_n370), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n730), .A2(new_n225), .ZN(new_n751));
  XOR2_X1   g0551(.A(KEYINPUT102), .B(G159), .Z(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n721), .ZN(new_n754));
  XNOR2_X1  g0554(.A(new_n754), .B(KEYINPUT32), .ZN(new_n755));
  INV_X1    g0555(.A(new_n740), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G97), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n755), .A2(new_n284), .A3(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n718), .ZN(new_n759));
  OAI22_X1  g0559(.A1(new_n759), .A2(new_n202), .B1(new_n725), .B2(new_n223), .ZN(new_n760));
  NOR4_X1   g0560(.A1(new_n750), .A2(new_n751), .A3(new_n758), .A4(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n715), .B1(new_n744), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n254), .A2(G45), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n662), .A2(new_n284), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n763), .B(new_n764), .C1(new_n241), .C2(G45), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n662), .A2(new_n298), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  XOR2_X1   g0567(.A(G355), .B(KEYINPUT99), .Z(new_n768));
  OAI221_X1 g0568(.A(new_n765), .B1(G116), .B2(new_n217), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n713), .A2(new_n715), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n714), .A2(new_n762), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n709), .A2(new_n772), .ZN(G396));
  INV_X1    g0573(.A(G143), .ZN(new_n774));
  INV_X1    g0574(.A(G150), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n759), .A2(new_n774), .B1(new_n775), .B2(new_n735), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G137), .B2(new_n726), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n777), .B1(new_n749), .B2(new_n753), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT34), .ZN(new_n779));
  OAI221_X1 g0579(.A(new_n779), .B1(new_n223), .B2(new_n742), .C1(new_n202), .C2(new_n740), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n730), .A2(new_n203), .ZN(new_n781));
  INV_X1    g0581(.A(G132), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n721), .A2(new_n782), .ZN(new_n783));
  NOR4_X1   g0583(.A1(new_n780), .A2(new_n298), .A3(new_n781), .A4(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(G294), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n757), .B1(new_n785), .B2(new_n759), .C1(new_n749), .C2(new_n556), .ZN(new_n786));
  INV_X1    g0586(.A(G311), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n730), .A2(new_n228), .B1(new_n721), .B2(new_n787), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT104), .ZN(new_n789));
  XOR2_X1   g0589(.A(KEYINPUT103), .B(G283), .Z(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n735), .ZN(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n298), .B1(new_n742), .B2(new_n225), .C1(new_n793), .C2(new_n725), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n786), .A2(new_n789), .A3(new_n792), .A4(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n715), .B1(new_n784), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n643), .A2(new_n397), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n457), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(new_n407), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n407), .A2(new_n643), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(new_n712), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n715), .A2(new_n711), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(new_n370), .ZN(new_n806));
  NAND4_X1  g0606(.A1(new_n796), .A2(new_n705), .A3(new_n804), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n677), .A2(new_n803), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n625), .A2(new_n802), .A3(new_n674), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n710), .B1(new_n810), .B2(new_n698), .ZN(new_n811));
  XOR2_X1   g0611(.A(new_n811), .B(KEYINPUT105), .Z(new_n812));
  AND2_X1   g0612(.A1(new_n810), .A2(new_n698), .ZN(new_n813));
  OAI21_X1  g0613(.A(new_n807), .B1(new_n812), .B2(new_n813), .ZN(G384));
  INV_X1    g0614(.A(KEYINPUT35), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n239), .B1(new_n524), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g0616(.A(new_n816), .B(G116), .C1(new_n815), .C2(new_n524), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT36), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n289), .A2(G77), .A3(new_n290), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n240), .A2(new_n819), .B1(G50), .B2(new_n203), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n820), .A2(G1), .A3(new_n215), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n297), .B1(new_n301), .B2(new_n203), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n272), .A2(KEYINPUT106), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n822), .B(new_n823), .Z(new_n824));
  OAI21_X1  g0624(.A(new_n269), .B1(new_n824), .B2(new_n263), .ZN(new_n825));
  INV_X1    g0625(.A(new_n641), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n355), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g0629(.A1(new_n346), .A2(KEYINPUT107), .A3(new_n826), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT107), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(new_n307), .B2(new_n641), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n335), .A2(new_n329), .B1(new_n346), .B2(new_n350), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT37), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n825), .B1(new_n350), .B2(new_n826), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(new_n332), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n836), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  AND3_X1   g0639(.A1(new_n829), .A2(KEYINPUT38), .A3(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(KEYINPUT38), .B1(new_n829), .B2(new_n839), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n801), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n809), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n426), .A2(new_n643), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n452), .A2(new_n455), .A3(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n629), .A2(new_n426), .A3(new_n643), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  OAI22_X1  g0649(.A1(new_n842), .A2(new_n849), .B1(new_n353), .B2(new_n826), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n452), .A2(new_n643), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT39), .B1(new_n840), .B2(new_n841), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT108), .ZN(new_n853));
  AND3_X1   g0653(.A1(new_n833), .A2(new_n834), .A3(new_n835), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n835), .B1(new_n833), .B2(new_n834), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT107), .B1(new_n346), .B2(new_n826), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n307), .A2(new_n831), .A3(new_n641), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n351), .A2(new_n332), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT37), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n861), .A2(KEYINPUT108), .A3(new_n836), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n351), .B(KEYINPUT18), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n859), .B1(new_n863), .B2(new_n337), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n856), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n829), .A2(KEYINPUT38), .A3(new_n839), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n852), .B1(KEYINPUT39), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n850), .B1(new_n851), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n679), .A2(new_n459), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(new_n634), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n871), .B(new_n873), .Z(new_n874));
  NAND3_X1  g0674(.A1(new_n697), .A2(new_n802), .A3(new_n848), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT40), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n867), .A2(KEYINPUT109), .A3(new_n868), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT109), .B1(new_n867), .B2(new_n868), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n877), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n876), .B1(new_n842), .B2(new_n875), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n880), .A2(G330), .A3(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n698), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n459), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n880), .A2(new_n459), .A3(new_n697), .A4(new_n881), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI22_X1  g0687(.A1(new_n874), .A2(new_n887), .B1(new_n210), .B2(new_n636), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT110), .Z(new_n889));
  AND2_X1   g0689(.A1(new_n874), .A2(new_n887), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n818), .B(new_n821), .C1(new_n889), .C2(new_n890), .ZN(G367));
  NAND2_X1  g0691(.A1(new_n620), .A2(new_n643), .ZN(new_n892));
  XOR2_X1   g0692(.A(new_n892), .B(KEYINPUT112), .Z(new_n893));
  OAI21_X1  g0693(.A(new_n616), .B1(new_n544), .B2(new_n674), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g0695(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n896), .A2(new_n659), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT42), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n543), .B1(new_n896), .B2(new_n569), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(new_n674), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n615), .B1(new_n609), .B2(new_n674), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT111), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n609), .A2(new_n674), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n904), .A2(new_n607), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n901), .A2(new_n902), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n903), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n898), .A2(new_n900), .B1(KEYINPUT43), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n907), .A2(KEYINPUT43), .ZN(new_n909));
  XNOR2_X1  g0709(.A(new_n908), .B(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n655), .A2(new_n895), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n910), .B(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n663), .B(KEYINPUT41), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n660), .A2(new_n895), .ZN(new_n915));
  XOR2_X1   g0715(.A(new_n915), .B(KEYINPUT45), .Z(new_n916));
  NOR2_X1   g0716(.A1(new_n660), .A2(new_n895), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT44), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(new_n656), .ZN(new_n920));
  OAI21_X1  g0720(.A(KEYINPUT113), .B1(new_n653), .B2(new_n658), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(new_n659), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n702), .A2(new_n922), .ZN(new_n923));
  OR2_X1    g0723(.A1(new_n922), .A2(new_n648), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n700), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n920), .A2(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n914), .B1(new_n927), .B2(new_n700), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n703), .B(KEYINPUT114), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n912), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n749), .A2(new_n791), .B1(new_n787), .B2(new_n725), .ZN(new_n931));
  INV_X1    g0731(.A(G317), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n721), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n730), .A2(new_n432), .ZN(new_n934));
  NOR4_X1   g0734(.A1(new_n931), .A2(new_n284), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n736), .A2(new_n470), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n743), .A2(G116), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT46), .ZN(new_n938));
  AOI22_X1  g0738(.A1(new_n718), .A2(G303), .B1(G107), .B2(new_n756), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n935), .A2(new_n936), .A3(new_n938), .A4(new_n939), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n742), .A2(new_n202), .B1(new_n740), .B2(new_n203), .ZN(new_n941));
  INV_X1    g0741(.A(new_n749), .ZN(new_n942));
  AOI22_X1  g0742(.A1(new_n942), .A2(G50), .B1(new_n736), .B2(new_n752), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n943), .A2(KEYINPUT115), .ZN(new_n944));
  AOI211_X1 g0744(.A(new_n941), .B(new_n944), .C1(G150), .C2(new_n718), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n298), .B1(new_n731), .B2(G77), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n722), .A2(G137), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n943), .A2(KEYINPUT115), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n945), .A2(new_n946), .A3(new_n947), .A4(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n725), .A2(new_n774), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n940), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT47), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n715), .ZN(new_n953));
  NAND4_X1  g0753(.A1(new_n903), .A2(new_n713), .A3(new_n905), .A4(new_n906), .ZN(new_n954));
  INV_X1    g0754(.A(new_n764), .ZN(new_n955));
  OAI221_X1 g0755(.A(new_n770), .B1(new_n217), .B2(new_n394), .C1(new_n955), .C2(new_n250), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n953), .A2(new_n705), .A3(new_n954), .A4(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n930), .A2(new_n957), .ZN(G387));
  NAND3_X1  g0758(.A1(new_n923), .A2(new_n924), .A3(new_n929), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n759), .A2(new_n932), .B1(new_n787), .B2(new_n735), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n960), .B1(G322), .B2(new_n726), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n793), .B2(new_n749), .ZN(new_n962));
  XNOR2_X1  g0762(.A(new_n962), .B(KEYINPUT48), .ZN(new_n963));
  OAI221_X1 g0763(.A(new_n963), .B1(new_n739), .B2(new_n742), .C1(new_n740), .C2(new_n791), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n964), .B(KEYINPUT49), .ZN(new_n965));
  AOI22_X1  g0765(.A1(G116), .A2(new_n731), .B1(new_n722), .B2(G326), .ZN(new_n966));
  AND3_X1   g0766(.A1(new_n965), .A2(new_n298), .A3(new_n966), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n742), .A2(new_n370), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n578), .A2(new_n756), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n968), .B(new_n969), .C1(G159), .C2(new_n726), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n736), .A2(new_n266), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n284), .B1(new_n746), .B2(new_n203), .ZN(new_n972));
  AOI211_X1 g0772(.A(new_n934), .B(new_n972), .C1(G150), .C2(new_n722), .ZN(new_n973));
  NAND3_X1  g0773(.A1(new_n970), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(G50), .B2(new_n718), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n715), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n247), .A2(new_n317), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n977), .A2(new_n764), .B1(new_n664), .B2(new_n766), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n266), .A2(new_n223), .ZN(new_n979));
  XNOR2_X1  g0779(.A(KEYINPUT116), .B(KEYINPUT50), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n979), .B(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n203), .A2(new_n370), .ZN(new_n982));
  NOR4_X1   g0782(.A1(new_n981), .A2(G45), .A3(new_n982), .A4(new_n664), .ZN(new_n983));
  OAI22_X1  g0783(.A1(new_n978), .A2(new_n983), .B1(G107), .B2(new_n217), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n770), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n654), .A2(new_n713), .ZN(new_n986));
  NAND4_X1  g0786(.A1(new_n976), .A2(new_n705), .A3(new_n985), .A4(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n700), .B1(new_n923), .B2(new_n924), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(KEYINPUT117), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n663), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n925), .B1(new_n988), .B2(KEYINPUT117), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n959), .B(new_n987), .C1(new_n990), .C2(new_n991), .ZN(G393));
  XOR2_X1   g0792(.A(new_n920), .B(KEYINPUT118), .Z(new_n993));
  NAND2_X1  g0793(.A1(new_n993), .A2(new_n929), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n710), .B1(new_n896), .B2(new_n713), .ZN(new_n995));
  OAI221_X1 g0795(.A(new_n770), .B1(new_n432), .B2(new_n217), .C1(new_n955), .C2(new_n258), .ZN(new_n996));
  AOI22_X1  g0796(.A1(G50), .A2(new_n736), .B1(new_n731), .B2(G87), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n718), .A2(G159), .B1(new_n726), .B2(G150), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n997), .B1(new_n370), .B2(new_n740), .C1(new_n998), .C2(KEYINPUT51), .ZN(new_n999));
  AOI22_X1  g0799(.A1(new_n942), .A2(new_n266), .B1(KEYINPUT51), .B2(new_n998), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n1000), .B(new_n284), .C1(new_n774), .C2(new_n721), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n999), .B(new_n1001), .C1(G68), .C2(new_n743), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n718), .A2(G311), .B1(new_n726), .B2(G317), .ZN(new_n1003));
  XOR2_X1   g0803(.A(new_n1003), .B(KEYINPUT52), .Z(new_n1004));
  NAND2_X1  g0804(.A1(new_n722), .A2(G322), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n743), .A2(new_n790), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n746), .A2(new_n785), .B1(new_n735), .B2(new_n793), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(G116), .B2(new_n756), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1004), .A2(new_n1005), .A3(new_n1006), .A4(new_n1008), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n1009), .A2(new_n284), .A3(new_n751), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n715), .B1(new_n1002), .B2(new_n1010), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n995), .A2(new_n996), .A3(new_n1011), .ZN(new_n1012));
  OR2_X1    g0812(.A1(new_n920), .A2(new_n926), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1013), .A2(new_n663), .A3(new_n927), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n994), .A2(new_n1012), .A3(new_n1014), .ZN(G390));
  XOR2_X1   g0815(.A(KEYINPUT54), .B(G143), .Z(new_n1016));
  AOI22_X1  g0816(.A1(new_n942), .A2(new_n1016), .B1(G137), .B2(new_n736), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n1017), .B(new_n284), .C1(new_n223), .C2(new_n730), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n759), .A2(new_n782), .ZN(new_n1019));
  INV_X1    g0819(.A(G125), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n721), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(G159), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n740), .A2(new_n1022), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1018), .A2(new_n1019), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n742), .A2(new_n775), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT53), .ZN(new_n1026));
  INV_X1    g0826(.A(G128), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1024), .B(new_n1026), .C1(new_n1027), .C2(new_n725), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT120), .ZN(new_n1029));
  NOR2_X1   g0829(.A1(new_n735), .A2(new_n225), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n284), .B1(new_n942), .B2(G97), .ZN(new_n1031));
  OAI221_X1 g0831(.A(new_n1031), .B1(new_n370), .B2(new_n740), .C1(new_n785), .C2(new_n721), .ZN(new_n1032));
  AOI211_X1 g0832(.A(new_n1030), .B(new_n1032), .C1(G116), .C2(new_n718), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n726), .A2(G283), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1033), .A2(new_n745), .A3(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1029), .B1(new_n781), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n710), .B1(new_n1036), .B2(new_n715), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n805), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n712), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1037), .B1(new_n266), .B2(new_n1038), .C1(new_n870), .C2(new_n1039), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n697), .A2(G330), .A3(new_n802), .A4(new_n848), .ZN(new_n1041));
  INV_X1    g0841(.A(new_n851), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n843), .B1(new_n675), .B2(new_n800), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1043), .A2(new_n848), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1042), .B(new_n1044), .C1(new_n878), .C2(new_n879), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n849), .A2(new_n1042), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n852), .B(new_n1046), .C1(KEYINPUT39), .C2(new_n869), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1045), .A2(new_n1047), .A3(new_n1041), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n929), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n1040), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n663), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT119), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1041), .A2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n697), .A2(G330), .A3(new_n802), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n848), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1056), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n1043), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1041), .A2(new_n1057), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1059), .A2(new_n1041), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(new_n844), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  AND3_X1   g0866(.A1(new_n872), .A2(new_n634), .A3(new_n884), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1054), .B1(new_n1051), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1068), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1049), .A2(new_n1070), .A3(new_n1050), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1053), .B1(new_n1069), .B2(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(G378));
  NOR2_X1   g0873(.A1(new_n384), .A2(new_n641), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n391), .B(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1075), .B(new_n1076), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n882), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n880), .A2(new_n1077), .A3(G330), .A4(new_n881), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n1079), .A2(new_n871), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n871), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n1045), .A2(new_n1047), .A3(new_n1041), .ZN(new_n1083));
  NOR3_X1   g0883(.A1(new_n1083), .A2(new_n1048), .A3(new_n1068), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1067), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n1081), .A2(new_n1082), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT57), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1054), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1071), .A2(new_n1067), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1089), .B(KEYINPUT57), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n929), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n710), .B1(new_n1078), .B2(new_n712), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n735), .A2(new_n782), .ZN(new_n1094));
  AOI22_X1  g0894(.A1(new_n718), .A2(G128), .B1(new_n743), .B2(new_n1016), .ZN(new_n1095));
  XNOR2_X1  g0895(.A(new_n1095), .B(KEYINPUT121), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n1096), .B1(new_n1020), .B2(new_n725), .C1(new_n775), .C2(new_n740), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1094), .B(new_n1097), .C1(G137), .C2(new_n734), .ZN(new_n1098));
  INV_X1    g0898(.A(KEYINPUT59), .ZN(new_n1099));
  AOI21_X1  g0899(.A(G33), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g0900(.A(G41), .B1(new_n722), .B2(G124), .ZN(new_n1101));
  OAI211_X1 g0901(.A(new_n1100), .B(new_n1101), .C1(new_n730), .C2(new_n753), .ZN(new_n1102));
  NOR2_X1   g0902(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1103));
  AOI21_X1  g0903(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n1102), .A2(new_n1103), .B1(G50), .B2(new_n1104), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n735), .A2(new_n432), .ZN(new_n1106));
  AOI211_X1 g0906(.A(G41), .B(new_n284), .C1(new_n578), .C2(new_n734), .ZN(new_n1107));
  OAI221_X1 g0907(.A(new_n1107), .B1(new_n202), .B2(new_n730), .C1(new_n556), .C2(new_n725), .ZN(new_n1108));
  AOI211_X1 g0908(.A(new_n1106), .B(new_n1108), .C1(G283), .C2(new_n722), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n968), .B1(G68), .B2(new_n756), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n1109), .B(new_n1110), .C1(new_n225), .C2(new_n759), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT58), .Z(new_n1112));
  OAI21_X1  g0912(.A(new_n715), .B1(new_n1105), .B2(new_n1112), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1093), .B(new_n1113), .C1(G50), .C2(new_n1038), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1092), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1091), .A2(new_n1116), .ZN(G375));
  NAND3_X1  g0917(.A1(new_n1085), .A2(new_n1065), .A3(new_n1063), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n913), .A3(new_n1068), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n711), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n848), .A2(new_n1120), .B1(G68), .B2(new_n1038), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n721), .A2(new_n1027), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1016), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n284), .B1(new_n1022), .B2(new_n742), .C1(new_n1123), .C2(new_n735), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1122), .B(new_n1124), .C1(G150), .C2(new_n734), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n718), .A2(G137), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n756), .A2(G50), .ZN(new_n1127));
  AOI22_X1  g0927(.A1(G132), .A2(new_n726), .B1(new_n731), .B2(G58), .ZN(new_n1128));
  NAND4_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n742), .A2(new_n432), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n1130), .B(new_n969), .C1(G283), .C2(new_n718), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n298), .B1(new_n730), .B2(new_n370), .C1(new_n785), .C2(new_n725), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1132), .B1(G116), .B2(new_n736), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n1131), .B(new_n1133), .C1(new_n225), .C2(new_n749), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n721), .A2(new_n793), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1129), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n710), .B(new_n1121), .C1(new_n715), .C2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(new_n1066), .B2(new_n929), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1119), .A2(new_n1138), .ZN(G381));
  AOI21_X1  g0939(.A(new_n1115), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(new_n1072), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n930), .A2(new_n957), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(G390), .A2(G384), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(G393), .A2(G396), .A3(G381), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n1143), .A3(new_n1144), .A4(new_n1145), .ZN(G407));
  NAND2_X1  g0946(.A1(new_n642), .A2(G213), .ZN(new_n1147));
  OR2_X1    g0947(.A1(new_n1141), .A2(new_n1147), .ZN(new_n1148));
  OR2_X1    g0948(.A1(new_n1148), .A2(KEYINPUT122), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1148), .A2(KEYINPUT122), .ZN(new_n1150));
  NAND4_X1  g0950(.A1(new_n1149), .A2(G213), .A3(G407), .A4(new_n1150), .ZN(G409));
  INV_X1    g0951(.A(KEYINPUT123), .ZN(new_n1152));
  OAI211_X1 g0952(.A(new_n1089), .B(new_n913), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1072), .A2(new_n1153), .A3(new_n1092), .A4(new_n1114), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1147), .B(new_n1154), .C1(new_n1140), .C2(new_n1072), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT60), .ZN(new_n1156));
  OR2_X1    g0956(.A1(new_n1118), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1118), .A2(new_n1156), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1157), .A2(new_n663), .A3(new_n1068), .A4(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n1138), .ZN(new_n1160));
  XNOR2_X1  g0960(.A(new_n1160), .B(G384), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1152), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(G375), .A2(G378), .ZN(new_n1164));
  AND2_X1   g0964(.A1(new_n1154), .A2(new_n1147), .ZN(new_n1165));
  NAND4_X1  g0965(.A1(new_n1164), .A2(KEYINPUT123), .A3(new_n1161), .A4(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT63), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1167), .A2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g0969(.A(G393), .B(G396), .Z(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(G387), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1143), .A2(KEYINPUT125), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1171), .B1(new_n1172), .B2(new_n1170), .ZN(new_n1173));
  INV_X1    g0973(.A(G390), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(G390), .B(new_n1171), .C1(new_n1172), .C2(new_n1170), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1155), .A2(new_n1162), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(KEYINPUT63), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1169), .A2(new_n1177), .A3(new_n1179), .ZN(new_n1180));
  AND3_X1   g0980(.A1(new_n642), .A2(G213), .A3(G2897), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT124), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1181), .B1(new_n1162), .B2(new_n1182), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1161), .B(new_n1182), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n1183), .B(new_n1155), .C1(new_n1184), .C2(new_n1181), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT61), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1180), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT126), .ZN(new_n1189));
  INV_X1    g0989(.A(KEYINPUT62), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1167), .B2(new_n1190), .ZN(new_n1191));
  AOI211_X1 g0991(.A(KEYINPUT126), .B(KEYINPUT62), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1178), .A2(KEYINPUT62), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1187), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  AND3_X1   g0995(.A1(new_n1175), .A2(KEYINPUT127), .A3(new_n1176), .ZN(new_n1196));
  AOI21_X1  g0996(.A(KEYINPUT127), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1188), .B1(new_n1195), .B2(new_n1199), .ZN(G405));
  NAND2_X1  g1000(.A1(new_n1164), .A2(new_n1141), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(new_n1162), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1198), .B(new_n1202), .ZN(G402));
endmodule


