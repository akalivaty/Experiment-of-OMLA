//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 1 1 1 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 0 0 1 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1328, new_n1329;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  XOR2_X1   g0010(.A(new_n210), .B(KEYINPUT64), .Z(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OR2_X1    g0013(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(KEYINPUT65), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n216), .B(G250), .C1(G257), .C2(G264), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT66), .B(KEYINPUT0), .Z(new_n218));
  XNOR2_X1  g0018(.A(new_n217), .B(new_n218), .ZN(new_n219));
  NOR2_X1   g0019(.A1(G58), .A2(G68), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(G50), .ZN(new_n222));
  INV_X1    g0022(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G68), .A2(G238), .B1(G97), .B2(G257), .ZN(new_n228));
  NAND2_X1  g0028(.A1(G116), .A2(G270), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n228), .B(new_n229), .C1(new_n202), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(G50), .B2(G226), .ZN(new_n232));
  NAND2_X1  g0032(.A1(G87), .A2(G250), .ZN(new_n233));
  INV_X1    g0033(.A(G77), .ZN(new_n234));
  INV_X1    g0034(.A(G244), .ZN(new_n235));
  OAI211_X1 g0035(.A(new_n232), .B(new_n233), .C1(new_n234), .C2(new_n235), .ZN(new_n236));
  AND2_X1   g0036(.A1(G107), .A2(G264), .ZN(new_n237));
  OAI21_X1  g0037(.A(new_n212), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n238), .B(KEYINPUT1), .Z(new_n239));
  NAND3_X1  g0039(.A1(new_n219), .A2(new_n227), .A3(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT67), .ZN(G361));
  XNOR2_X1  g0041(.A(G238), .B(G244), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n242), .B(G232), .ZN(new_n243));
  XNOR2_X1  g0043(.A(KEYINPUT2), .B(G226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT68), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G250), .B(G257), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G264), .B(G270), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G358));
  XNOR2_X1  g0050(.A(G50), .B(G58), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n251), .B(KEYINPUT69), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G68), .B(G77), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G87), .B(G97), .ZN(new_n255));
  XNOR2_X1  g0055(.A(G107), .B(G116), .ZN(new_n256));
  XOR2_X1   g0056(.A(new_n255), .B(new_n256), .Z(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  INV_X1    g0058(.A(G1), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n259), .B1(G41), .B2(G45), .ZN(new_n260));
  INV_X1    g0060(.A(G274), .ZN(new_n261));
  NOR2_X1   g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G226), .ZN(new_n263));
  INV_X1    g0063(.A(G1698), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n230), .A2(G1698), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  OAI211_X1 g0068(.A(new_n265), .B(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G97), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n224), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND3_X1   g0076(.A1(new_n276), .A2(G238), .A3(new_n260), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT13), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT13), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n273), .A2(new_n281), .A3(new_n278), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n282), .A3(G190), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT11), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n225), .A2(G33), .A3(G77), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n203), .A2(G20), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n285), .B(new_n286), .C1(new_n288), .C2(new_n201), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT76), .ZN(new_n290));
  NAND3_X1  g0090(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(new_n224), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(new_n289), .B2(new_n292), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n284), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n289), .A2(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT76), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n289), .A2(new_n290), .A3(new_n292), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n297), .A2(KEYINPUT11), .A3(new_n298), .ZN(new_n299));
  NAND4_X1  g0099(.A1(new_n259), .A2(new_n203), .A3(G13), .A4(G20), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT12), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n259), .A2(G20), .ZN(new_n302));
  NAND4_X1  g0102(.A1(new_n302), .A2(new_n291), .A3(G68), .A4(new_n224), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n305));
  AND3_X1   g0105(.A1(new_n301), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AND3_X1   g0106(.A1(new_n295), .A2(new_n299), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n281), .B1(new_n273), .B2(new_n278), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n276), .B1(new_n269), .B2(new_n270), .ZN(new_n309));
  NOR4_X1   g0109(.A1(new_n309), .A2(new_n277), .A3(KEYINPUT13), .A4(new_n262), .ZN(new_n310));
  OAI21_X1  g0110(.A(G200), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n283), .A2(new_n307), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT78), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n283), .A2(new_n307), .A3(new_n311), .A4(KEYINPUT78), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(new_n307), .ZN(new_n317));
  OAI21_X1  g0117(.A(G169), .B1(new_n308), .B2(new_n310), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n318), .A2(KEYINPUT79), .A3(KEYINPUT14), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n280), .A2(new_n282), .ZN(new_n320));
  NAND2_X1  g0120(.A1(KEYINPUT79), .A2(KEYINPUT14), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(G169), .A3(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G179), .ZN(new_n323));
  OAI211_X1 g0123(.A(new_n319), .B(new_n322), .C1(new_n323), .C2(new_n320), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n316), .B1(new_n317), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n259), .A2(G13), .A3(G20), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G50), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  AND2_X1   g0128(.A1(new_n291), .A2(new_n224), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n329), .A2(KEYINPUT72), .A3(new_n326), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT72), .ZN(new_n331));
  INV_X1    g0131(.A(new_n326), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n292), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n330), .A2(new_n333), .A3(G50), .A4(new_n302), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n225), .A2(G33), .ZN(new_n335));
  AND2_X1   g0135(.A1(KEYINPUT8), .A2(G58), .ZN(new_n336));
  NOR2_X1   g0136(.A1(KEYINPUT8), .A2(G58), .ZN(new_n337));
  OAI21_X1  g0137(.A(KEYINPUT70), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT8), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n202), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT70), .ZN(new_n341));
  NAND2_X1  g0141(.A1(KEYINPUT8), .A2(G58), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n335), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(G150), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n288), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT71), .ZN(new_n347));
  AOI211_X1 g0147(.A(new_n347), .B(new_n225), .C1(new_n220), .C2(new_n201), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT71), .B1(new_n204), .B2(G20), .ZN(new_n349));
  NOR4_X1   g0149(.A1(new_n344), .A2(new_n346), .A3(new_n348), .A4(new_n349), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n328), .B(new_n334), .C1(new_n350), .C2(new_n329), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n264), .A2(G223), .ZN(new_n352));
  NOR2_X1   g0152(.A1(G222), .A2(G1698), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n352), .A2(new_n353), .B1(new_n267), .B2(new_n268), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT3), .ZN(new_n355));
  INV_X1    g0155(.A(G33), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n354), .B(new_n272), .C1(G77), .C2(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(new_n262), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n276), .A2(G226), .A3(new_n260), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(G169), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n363), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n323), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n351), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n329), .A2(G77), .A3(new_n302), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n340), .A2(new_n342), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n371), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n372));
  XOR2_X1   g0172(.A(KEYINPUT15), .B(G87), .Z(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n372), .B1(new_n335), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n369), .B1(new_n375), .B2(new_n292), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n326), .A2(G77), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n359), .A2(G232), .A3(new_n264), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n359), .A2(G238), .A3(G1698), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(new_n207), .C2(new_n359), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n272), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n276), .A2(new_n260), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n361), .B1(new_n384), .B2(new_n235), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT73), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  OAI211_X1 g0187(.A(new_n361), .B(KEYINPUT73), .C1(new_n384), .C2(new_n235), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n383), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(new_n364), .ZN(new_n390));
  NAND4_X1  g0190(.A1(new_n383), .A2(new_n323), .A3(new_n387), .A4(new_n388), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n379), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n389), .A2(G200), .ZN(new_n393));
  AOI211_X1 g0193(.A(new_n377), .B(new_n369), .C1(new_n375), .C2(new_n292), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n383), .A2(G190), .A3(new_n387), .A4(new_n388), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n392), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT9), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n351), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n363), .A2(G200), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT74), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n363), .A2(KEYINPUT74), .A3(G200), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n366), .A2(G190), .ZN(new_n406));
  NOR2_X1   g0206(.A1(new_n348), .A2(new_n349), .ZN(new_n407));
  INV_X1    g0207(.A(new_n346), .ZN(new_n408));
  AND2_X1   g0208(.A1(new_n338), .A2(new_n343), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n407), .B(new_n408), .C1(new_n335), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n292), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n411), .A2(KEYINPUT9), .A3(new_n328), .A4(new_n334), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n400), .A2(new_n405), .A3(new_n406), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(KEYINPUT10), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n368), .B(new_n398), .C1(new_n415), .C2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT75), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n325), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(new_n368), .ZN(new_n421));
  INV_X1    g0221(.A(new_n334), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n422), .B1(new_n410), .B2(new_n292), .ZN(new_n423));
  AOI21_X1  g0223(.A(KEYINPUT9), .B1(new_n423), .B2(new_n328), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n344), .A2(new_n346), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n329), .B1(new_n425), .B2(new_n407), .ZN(new_n426));
  NOR4_X1   g0226(.A1(new_n426), .A2(new_n422), .A3(new_n399), .A4(new_n327), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT10), .ZN(new_n429));
  NAND4_X1  g0229(.A1(new_n428), .A2(new_n429), .A3(new_n406), .A4(new_n405), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n421), .B1(new_n430), .B2(new_n414), .ZN(new_n431));
  AOI21_X1  g0231(.A(KEYINPUT75), .B1(new_n431), .B2(new_n398), .ZN(new_n432));
  XNOR2_X1  g0232(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n357), .A2(new_n225), .A3(new_n358), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT7), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n357), .A2(KEYINPUT7), .A3(new_n225), .A4(new_n358), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n203), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n202), .A2(new_n203), .ZN(new_n439));
  OAI21_X1  g0239(.A(G20), .B1(new_n439), .B2(new_n220), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n287), .A2(G159), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n433), .B1(new_n438), .B2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT81), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n436), .A2(new_n437), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n442), .B1(new_n446), .B2(G68), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n329), .B1(new_n447), .B2(KEYINPUT16), .ZN(new_n448));
  OAI211_X1 g0248(.A(KEYINPUT81), .B(new_n433), .C1(new_n438), .C2(new_n442), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n445), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n330), .A2(new_n333), .A3(new_n302), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n451), .A2(new_n409), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n452), .B1(new_n332), .B2(new_n409), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n263), .A2(G1698), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n455), .B1(G223), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n456));
  NAND2_X1  g0256(.A1(G33), .A2(G87), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n458), .A2(new_n272), .ZN(new_n459));
  AND2_X1   g0259(.A1(new_n276), .A2(new_n260), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n262), .B1(new_n460), .B2(G232), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n461), .A3(G179), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n276), .B1(new_n456), .B2(new_n457), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n361), .B1(new_n384), .B2(new_n230), .ZN(new_n464));
  OAI21_X1  g0264(.A(G169), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n454), .A2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT18), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT82), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n454), .A2(KEYINPUT18), .A3(new_n467), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT18), .B1(new_n454), .B2(new_n467), .ZN(new_n474));
  AOI211_X1 g0274(.A(new_n469), .B(new_n466), .C1(new_n450), .C2(new_n453), .ZN(new_n475));
  OAI21_X1  g0275(.A(KEYINPUT82), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n463), .A2(new_n464), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G190), .ZN(new_n478));
  OAI21_X1  g0278(.A(G200), .B1(new_n463), .B2(new_n464), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n450), .A2(new_n478), .A3(new_n453), .A4(new_n479), .ZN(new_n480));
  XNOR2_X1  g0280(.A(new_n480), .B(KEYINPUT17), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n473), .A2(new_n476), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n432), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g0283(.A(KEYINPUT83), .B1(new_n420), .B2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT83), .ZN(new_n485));
  NOR4_X1   g0285(.A1(new_n419), .A2(new_n432), .A3(new_n485), .A4(new_n482), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n267), .A2(new_n268), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(G303), .ZN(new_n489));
  OAI211_X1 g0289(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(new_n264), .C1(new_n267), .C2(new_n268), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n489), .A2(new_n490), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT88), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT88), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n489), .A2(new_n494), .A3(new_n490), .A4(new_n491), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n493), .A2(new_n272), .A3(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G45), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(G1), .ZN(new_n498));
  XNOR2_X1  g0298(.A(KEYINPUT5), .B(G41), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n272), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n259), .A2(G45), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(new_n261), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n500), .A2(G270), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n496), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n332), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n259), .A2(G33), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n326), .A2(new_n507), .A3(new_n224), .A4(new_n291), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(G116), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G283), .ZN(new_n511));
  OAI211_X1 g0311(.A(new_n511), .B(new_n225), .C1(G33), .C2(new_n206), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n292), .C1(new_n225), .C2(G116), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT20), .ZN(new_n514));
  AND2_X1   g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n513), .A2(new_n514), .ZN(new_n516));
  OAI211_X1 g0316(.A(new_n506), .B(new_n510), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND3_X1  g0317(.A1(new_n504), .A2(G169), .A3(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT21), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n496), .A2(G179), .A3(new_n503), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n517), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n504), .A2(KEYINPUT21), .A3(G169), .A4(new_n517), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n520), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(G250), .B(new_n264), .C1(new_n267), .C2(new_n268), .ZN(new_n526));
  OAI211_X1 g0326(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n527));
  NAND2_X1  g0327(.A1(G33), .A2(G294), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(new_n272), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n500), .A2(G264), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n502), .A2(new_n499), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT90), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n272), .A2(new_n529), .B1(new_n500), .B2(G264), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n535), .B1(new_n536), .B2(new_n532), .ZN(new_n537));
  OAI21_X1  g0337(.A(G169), .B1(new_n534), .B2(new_n537), .ZN(new_n538));
  NOR2_X1   g0338(.A1(new_n533), .A2(new_n323), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n225), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n542));
  XNOR2_X1  g0342(.A(KEYINPUT89), .B(KEYINPUT22), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT22), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(KEYINPUT89), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n359), .A2(new_n225), .A3(G87), .A4(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n225), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n544), .A2(new_n547), .A3(new_n551), .A4(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT24), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI22_X1  g0355(.A1(new_n542), .A2(new_n543), .B1(new_n549), .B2(new_n550), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n556), .A2(KEYINPUT24), .A3(new_n547), .A4(new_n552), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n292), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n509), .A2(G107), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n326), .A2(G107), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n560), .B(KEYINPUT25), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n558), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT91), .B1(new_n541), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n536), .A2(new_n535), .A3(new_n532), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n364), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(KEYINPUT91), .B(new_n562), .C1(new_n566), .C2(new_n539), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n525), .B1(new_n563), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n326), .A2(G97), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n446), .A2(G107), .ZN(new_n571));
  NAND2_X1  g0371(.A1(G97), .A2(G107), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n208), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n574), .ZN(new_n576));
  NAND2_X1  g0376(.A1(KEYINPUT6), .A2(G107), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n576), .A2(new_n208), .A3(new_n572), .A4(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(G20), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n288), .A2(new_n234), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n571), .A2(new_n580), .A3(new_n582), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n570), .B1(new_n583), .B2(new_n292), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n508), .A2(new_n206), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  OAI211_X1 g0386(.A(G244), .B(new_n264), .C1(new_n267), .C2(new_n268), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT85), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT4), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n587), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n359), .A2(G250), .A3(G1698), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n588), .A2(new_n589), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n359), .A2(G244), .A3(new_n264), .A4(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(KEYINPUT85), .A2(KEYINPUT4), .B1(G33), .B2(G283), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n590), .A2(new_n591), .A3(new_n593), .A4(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n272), .ZN(new_n596));
  AND2_X1   g0396(.A1(KEYINPUT5), .A2(G41), .ZN(new_n597));
  NOR2_X1   g0397(.A1(KEYINPUT5), .A2(G41), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n498), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n599), .A2(G257), .A3(new_n276), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n600), .A2(new_n532), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n584), .A2(new_n586), .B1(new_n364), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n595), .B2(new_n272), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n323), .ZN(new_n606));
  INV_X1    g0406(.A(G200), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  INV_X1    g0408(.A(G190), .ZN(new_n609));
  AOI211_X1 g0409(.A(new_n609), .B(new_n601), .C1(new_n595), .C2(new_n272), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(new_n570), .ZN(new_n612));
  AOI21_X1  g0412(.A(new_n207), .B1(new_n436), .B2(new_n437), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n225), .B1(new_n575), .B2(new_n578), .ZN(new_n614));
  NOR3_X1   g0414(.A1(new_n613), .A2(new_n614), .A3(new_n581), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n612), .B(new_n586), .C1(new_n615), .C2(new_n329), .ZN(new_n616));
  INV_X1    g0416(.A(new_n616), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n604), .A2(new_n606), .B1(new_n611), .B2(new_n617), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n564), .A2(new_n565), .A3(new_n609), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n533), .A2(new_n607), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n621), .A2(new_n559), .A3(new_n561), .A4(new_n558), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n504), .A2(G200), .ZN(new_n623));
  INV_X1    g0423(.A(new_n517), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n623), .B(new_n624), .C1(new_n609), .C2(new_n504), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n235), .A2(G1698), .ZN(new_n626));
  OAI221_X1 g0426(.A(new_n626), .B1(G238), .B2(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n627));
  NAND2_X1  g0427(.A1(G33), .A2(G116), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n276), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n276), .A2(G250), .A3(new_n501), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NOR3_X1   g0431(.A1(new_n629), .A2(new_n502), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n323), .ZN(new_n633));
  NOR2_X1   g0433(.A1(new_n373), .A2(new_n326), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n359), .A2(new_n225), .A3(G68), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT19), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n636), .B1(new_n335), .B2(new_n206), .ZN(new_n637));
  NOR3_X1   g0437(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT86), .ZN(new_n639));
  XNOR2_X1  g0439(.A(new_n638), .B(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n270), .A2(new_n636), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(G20), .ZN(new_n642));
  OAI211_X1 g0442(.A(new_n635), .B(new_n637), .C1(new_n640), .C2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n634), .B1(new_n643), .B2(new_n292), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n509), .A2(new_n373), .ZN(new_n645));
  INV_X1    g0445(.A(new_n502), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n627), .A2(new_n628), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n646), .B(new_n630), .C1(new_n647), .C2(new_n276), .ZN(new_n648));
  AOI22_X1  g0448(.A1(new_n644), .A2(new_n645), .B1(new_n364), .B2(new_n648), .ZN(new_n649));
  NOR4_X1   g0449(.A1(new_n629), .A2(new_n631), .A3(new_n609), .A4(new_n502), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n650), .B1(G200), .B2(new_n648), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n643), .A2(new_n292), .ZN(new_n652));
  INV_X1    g0452(.A(new_n634), .ZN(new_n653));
  INV_X1    g0453(.A(G87), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n508), .A2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(KEYINPUT87), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n655), .B(new_n656), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n652), .A2(new_n653), .A3(new_n657), .ZN(new_n658));
  AOI22_X1  g0458(.A1(new_n633), .A2(new_n649), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n618), .A2(new_n622), .A3(new_n625), .A4(new_n659), .ZN(new_n660));
  NOR3_X1   g0460(.A1(new_n487), .A2(new_n569), .A3(new_n660), .ZN(G372));
  NOR2_X1   g0461(.A1(new_n474), .A2(new_n475), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n392), .A2(KEYINPUT92), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT92), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n379), .A2(new_n390), .A3(new_n665), .A4(new_n391), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n667), .A2(new_n312), .B1(new_n324), .B2(new_n317), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT17), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n480), .B(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n663), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n430), .A2(new_n414), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n421), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n603), .A2(G200), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n605), .A2(G190), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n674), .A2(new_n584), .A3(new_n586), .A4(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n603), .A2(new_n364), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n677), .A2(new_n616), .A3(new_n606), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n562), .B1(new_n619), .B2(new_n620), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n652), .A2(new_n645), .A3(new_n653), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n648), .A2(new_n364), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(new_n633), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n648), .A2(G200), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n632), .A2(G190), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(new_n644), .A4(new_n657), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n679), .A2(new_n680), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n562), .B1(new_n566), .B2(new_n539), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n689), .A2(new_n522), .A3(new_n523), .A4(new_n520), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n683), .ZN(new_n692));
  INV_X1    g0492(.A(new_n678), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n659), .A2(new_n693), .A3(KEYINPUT26), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT26), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n687), .B2(new_n678), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n692), .B1(new_n694), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g0497(.A1(new_n691), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n673), .B1(new_n487), .B2(new_n698), .ZN(G369));
  INV_X1    g0499(.A(G13), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n700), .A2(G20), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  OR3_X1    g0502(.A1(new_n702), .A2(KEYINPUT27), .A3(G1), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT27), .B1(new_n702), .B2(G1), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n703), .A2(G213), .A3(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(G343), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n707), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n624), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g0509(.A(new_n524), .B(new_n709), .ZN(new_n710));
  AND2_X1   g0510(.A1(new_n710), .A2(new_n625), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n711), .A2(G330), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT91), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n689), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(new_n567), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n680), .B1(new_n562), .B2(new_n707), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n541), .A2(new_n562), .A3(new_n707), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n712), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n524), .A2(new_n708), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT93), .ZN(new_n722));
  AND2_X1   g0522(.A1(new_n541), .A2(new_n562), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n722), .A2(new_n719), .B1(new_n723), .B2(new_n708), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n720), .A2(new_n724), .ZN(G399));
  INV_X1    g0525(.A(new_n216), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G41), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n640), .A2(new_n505), .ZN(new_n728));
  NOR3_X1   g0528(.A1(new_n727), .A2(new_n259), .A3(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n223), .B2(new_n727), .ZN(new_n730));
  XOR2_X1   g0530(.A(new_n730), .B(KEYINPUT28), .Z(new_n731));
  AOI21_X1  g0531(.A(new_n707), .B1(new_n691), .B2(new_n697), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT29), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n569), .A2(new_n688), .ZN(new_n735));
  AOI21_X1  g0535(.A(new_n707), .B1(new_n735), .B2(new_n697), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n734), .B1(new_n736), .B2(new_n733), .ZN(new_n737));
  INV_X1    g0537(.A(G330), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n524), .B1(new_n714), .B2(new_n567), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n739), .A2(new_n688), .A3(new_n625), .A4(new_n708), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n632), .A2(new_n536), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND4_X1  g0542(.A1(new_n521), .A2(new_n742), .A3(KEYINPUT30), .A4(new_n605), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT30), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n605), .A2(new_n496), .A3(G179), .A4(new_n503), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n744), .B1(new_n745), .B2(new_n741), .ZN(new_n746));
  AOI21_X1  g0546(.A(G179), .B1(new_n496), .B2(new_n503), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n747), .A2(new_n533), .A3(new_n603), .A4(new_n648), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n743), .A2(new_n746), .A3(new_n748), .ZN(new_n749));
  AND3_X1   g0549(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n750));
  AOI21_X1  g0550(.A(KEYINPUT31), .B1(new_n749), .B2(new_n707), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n738), .B1(new_n740), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n737), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n731), .B1(new_n754), .B2(G1), .ZN(G364));
  NAND2_X1  g0555(.A1(G355), .A2(new_n359), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n223), .A2(G45), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n757), .B1(new_n254), .B2(G45), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n216), .B(new_n756), .C1(new_n758), .C2(new_n359), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n274), .B1(new_n225), .B2(G169), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n760), .A2(KEYINPUT94), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n760), .A2(KEYINPUT94), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(G13), .A2(G33), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n765), .A2(G20), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n759), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n768), .B1(G116), .B2(new_n726), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n609), .A2(G20), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT97), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n771), .A2(new_n323), .A3(new_n607), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT98), .ZN(new_n773));
  OR2_X1    g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n772), .A2(new_n773), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g0576(.A(G159), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NAND2_X1  g0579(.A1(G20), .A2(G179), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT95), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n609), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT96), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n609), .A2(new_n607), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n784), .A2(new_n202), .B1(new_n201), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n771), .A2(new_n323), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G107), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n781), .A2(new_n609), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n790), .B(new_n359), .C1(new_n234), .C2(new_n793), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n791), .A2(new_n607), .ZN(new_n795));
  AOI211_X1 g0595(.A(new_n787), .B(new_n794), .C1(G68), .C2(new_n795), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n785), .A2(G20), .A3(new_n323), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT99), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT99), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G87), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n225), .B1(new_n782), .B2(new_n323), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n803), .A2(new_n206), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n779), .A2(new_n796), .A3(new_n802), .A4(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n776), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G329), .ZN(new_n808));
  INV_X1    g0608(.A(G294), .ZN(new_n809));
  INV_X1    g0609(.A(new_n795), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT33), .B(G317), .Z(new_n811));
  OAI221_X1 g0611(.A(new_n808), .B1(new_n809), .B2(new_n803), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G283), .B2(new_n789), .ZN(new_n813));
  INV_X1    g0613(.A(G303), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n488), .B1(new_n800), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n786), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n815), .B1(G326), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(G311), .ZN(new_n818));
  OAI211_X1 g0618(.A(new_n813), .B(new_n817), .C1(new_n818), .C2(new_n793), .ZN(new_n819));
  INV_X1    g0619(.A(G322), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n783), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n806), .B1(new_n819), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n769), .B1(new_n822), .B2(new_n763), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n259), .B1(new_n701), .B2(G45), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n727), .A2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n766), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n823), .B(new_n826), .C1(new_n711), .C2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n711), .A2(G330), .ZN(new_n830));
  NOR3_X1   g0630(.A1(new_n712), .A2(new_n830), .A3(new_n826), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n832), .ZN(G396));
  NOR2_X1   g0633(.A1(new_n763), .A2(new_n764), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n826), .B1(G77), .B2(new_n835), .ZN(new_n836));
  XOR2_X1   g0636(.A(new_n836), .B(KEYINPUT100), .Z(new_n837));
  NAND2_X1  g0637(.A1(new_n379), .A2(new_n707), .ZN(new_n838));
  AND3_X1   g0638(.A1(new_n392), .A2(new_n396), .A3(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n838), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(new_n667), .B2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n789), .A2(G87), .ZN(new_n843));
  INV_X1    g0643(.A(G283), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n843), .B1(new_n793), .B2(new_n505), .C1(new_n844), .C2(new_n810), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n804), .B(new_n845), .C1(G303), .C2(new_n816), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n807), .A2(G311), .ZN(new_n847));
  INV_X1    g0647(.A(new_n783), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n801), .A2(G107), .B1(G294), .B2(new_n848), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n488), .A3(new_n847), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n795), .A2(G150), .B1(new_n816), .B2(G137), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n851), .B1(new_n777), .B2(new_n793), .ZN(new_n852));
  INV_X1    g0652(.A(new_n784), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n852), .B1(G143), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g0654(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n854), .A2(new_n855), .B1(G50), .B2(new_n801), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n856), .B1(new_n855), .B2(new_n854), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n788), .A2(new_n203), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n359), .B1(new_n803), .B2(new_n202), .ZN(new_n859));
  OR3_X1    g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g0660(.A(G132), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n776), .A2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n850), .B1(new_n860), .B2(new_n862), .ZN(new_n863));
  XOR2_X1   g0663(.A(new_n863), .B(KEYINPUT102), .Z(new_n864));
  INV_X1    g0664(.A(new_n763), .ZN(new_n865));
  OAI221_X1 g0665(.A(new_n837), .B1(new_n765), .B2(new_n842), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  XNOR2_X1  g0666(.A(new_n732), .B(new_n842), .ZN(new_n867));
  XNOR2_X1  g0667(.A(new_n867), .B(new_n753), .ZN(new_n868));
  INV_X1    g0668(.A(new_n826), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n866), .A2(new_n870), .ZN(G384));
  INV_X1    g0671(.A(new_n487), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n317), .B(new_n707), .C1(new_n316), .C2(new_n324), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n324), .A2(new_n317), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n317), .A2(new_n707), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n875), .A2(new_n312), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n841), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NOR3_X1   g0678(.A1(new_n569), .A2(new_n660), .A3(new_n707), .ZN(new_n879));
  INV_X1    g0679(.A(new_n751), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n749), .A2(KEYINPUT31), .A3(new_n707), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n878), .B1(new_n879), .B2(new_n882), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT105), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(KEYINPUT40), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n740), .A2(new_n752), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(KEYINPUT105), .A3(new_n878), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT38), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT37), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n466), .A2(new_n705), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n447), .A2(KEYINPUT16), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n292), .A3(new_n443), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n453), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n480), .B2(new_n895), .ZN(new_n896));
  AND4_X1   g0696(.A1(new_n478), .A2(new_n450), .A3(new_n453), .A4(new_n479), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n450), .A2(new_n453), .B1(new_n466), .B2(new_n705), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n899), .B2(new_n890), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n705), .B1(new_n893), .B2(new_n453), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n889), .B(new_n900), .C1(new_n482), .C2(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(KEYINPUT37), .B1(new_n897), .B2(new_n898), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(KEYINPUT104), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n899), .A2(new_n890), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT104), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(KEYINPUT37), .C1(new_n897), .C2(new_n898), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n705), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n454), .B(new_n909), .C1(new_n670), .C2(new_n662), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT38), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n888), .B1(new_n902), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(KEYINPUT106), .B1(new_n886), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT40), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n883), .B2(new_n884), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n908), .A2(new_n910), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n889), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n482), .A2(new_n901), .ZN(new_n918));
  INV_X1    g0718(.A(new_n900), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(KEYINPUT38), .A3(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n917), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT106), .ZN(new_n922));
  NAND4_X1  g0722(.A1(new_n915), .A2(new_n921), .A3(new_n922), .A4(new_n888), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n913), .A2(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n883), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n918), .B2(new_n919), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n925), .B1(new_n926), .B2(new_n902), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n914), .ZN(new_n928));
  AND4_X1   g0728(.A1(new_n872), .A2(new_n924), .A3(new_n887), .A4(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n738), .B1(new_n927), .B2(new_n914), .ZN(new_n930));
  AOI22_X1  g0730(.A1(new_n925), .A2(KEYINPUT105), .B1(new_n917), .B2(new_n920), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n922), .B1(new_n931), .B2(new_n915), .ZN(new_n932));
  AND4_X1   g0732(.A1(new_n922), .A2(new_n915), .A3(new_n888), .A4(new_n921), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n930), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(G330), .B(new_n887), .C1(new_n484), .C2(new_n486), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n929), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT107), .Z(new_n937));
  OAI21_X1  g0737(.A(KEYINPUT39), .B1(new_n926), .B2(new_n902), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT39), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n917), .A2(new_n920), .A3(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n324), .A2(new_n317), .A3(new_n708), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OR2_X1    g0743(.A1(new_n392), .A2(new_n707), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT103), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n732), .B2(new_n842), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n873), .A2(new_n877), .ZN(new_n948));
  OAI211_X1 g0748(.A(new_n947), .B(new_n948), .C1(new_n902), .C2(new_n926), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n663), .B2(new_n909), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n943), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n737), .B1(new_n484), .B2(new_n486), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n952), .A2(new_n673), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n951), .B(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n937), .A2(new_n954), .B1(G1), .B2(new_n702), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n955), .B(KEYINPUT108), .Z(new_n956));
  OAI21_X1  g0756(.A(new_n956), .B1(new_n937), .B2(new_n954), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n505), .B1(new_n579), .B2(KEYINPUT35), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n958), .B(new_n226), .C1(KEYINPUT35), .C2(new_n579), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n959), .B(KEYINPUT36), .ZN(new_n960));
  OAI21_X1  g0760(.A(G77), .B1(new_n202), .B2(new_n203), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n222), .A2(new_n961), .B1(G50), .B2(new_n203), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(G1), .A3(new_n700), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n957), .A2(new_n960), .A3(new_n963), .ZN(G367));
  OAI21_X1  g0764(.A(new_n618), .B1(new_n617), .B2(new_n708), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n678), .B2(new_n708), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n722), .A2(new_n719), .A3(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT42), .Z(new_n968));
  OAI21_X1  g0768(.A(new_n678), .B1(new_n965), .B2(new_n715), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n708), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n658), .A2(new_n708), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n687), .A2(new_n971), .ZN(new_n972));
  OR2_X1    g0772(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n692), .A2(new_n971), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(KEYINPUT109), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n968), .A2(new_n970), .B1(KEYINPUT43), .B2(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n977), .B(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n720), .ZN(new_n980));
  AND2_X1   g0780(.A1(new_n980), .A2(new_n966), .ZN(new_n981));
  OR2_X1    g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n979), .A2(new_n981), .ZN(new_n983));
  XNOR2_X1  g0783(.A(KEYINPUT110), .B(KEYINPUT41), .ZN(new_n984));
  XOR2_X1   g0784(.A(new_n727), .B(new_n984), .Z(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n712), .B(new_n719), .ZN(new_n987));
  INV_X1    g0787(.A(new_n722), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n754), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT111), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n724), .A2(new_n992), .A3(new_n966), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT45), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n724), .B2(new_n966), .ZN(new_n996));
  OR3_X1    g0796(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n724), .A2(new_n966), .ZN(new_n998));
  XNOR2_X1  g0798(.A(new_n998), .B(KEYINPUT44), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n995), .B1(new_n994), .B2(new_n996), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n997), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n980), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n997), .A2(new_n720), .A3(new_n999), .A4(new_n1000), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n991), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n986), .B1(new_n1004), .B2(new_n754), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n982), .B(new_n983), .C1(new_n1005), .C2(new_n825), .ZN(new_n1006));
  INV_X1    g0806(.A(new_n976), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n869), .B1(new_n1007), .B2(new_n766), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n216), .A2(new_n488), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n767), .B1(new_n216), .B2(new_n374), .C1(new_n1009), .C2(new_n249), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n807), .A2(G137), .B1(G58), .B2(new_n801), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT112), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(new_n789), .A2(G77), .B1(new_n792), .B2(G50), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1013), .A2(new_n359), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n795), .A2(G159), .B1(new_n848), .B2(G150), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n203), .B2(new_n803), .C1(new_n1011), .C2(new_n1012), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n1015), .B(new_n1017), .C1(G143), .C2(new_n816), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n792), .A2(G283), .B1(new_n816), .B2(G311), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n1019), .B1(new_n809), .B2(new_n810), .C1(new_n784), .C2(new_n814), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n800), .A2(new_n505), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n1021), .A2(KEYINPUT46), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n359), .B1(new_n1021), .B2(KEYINPUT46), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n803), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(G107), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n789), .A2(G97), .ZN(new_n1026));
  NAND4_X1  g0826(.A1(new_n1022), .A2(new_n1023), .A3(new_n1025), .A4(new_n1026), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n1020), .B(new_n1027), .C1(G317), .C2(new_n807), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n1018), .A2(new_n1028), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT47), .ZN(new_n1030));
  OAI211_X1 g0830(.A(new_n1008), .B(new_n1010), .C1(new_n1030), .C2(new_n865), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1006), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(KEYINPUT113), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT113), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1006), .A2(new_n1034), .A3(new_n1031), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(G387));
  INV_X1    g0836(.A(new_n991), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n727), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n989), .B2(new_n990), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n719), .A2(new_n827), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n371), .A2(new_n201), .ZN(new_n1042));
  AOI21_X1  g0842(.A(G45), .B1(new_n1042), .B2(KEYINPUT50), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(KEYINPUT50), .B2(new_n1042), .C1(new_n203), .C2(new_n234), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n728), .B1(new_n1044), .B2(new_n488), .ZN(new_n1045));
  NOR3_X1   g0845(.A1(new_n245), .A2(new_n497), .A3(new_n359), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n216), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1047), .B(new_n767), .C1(new_n207), .C2(new_n216), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n800), .A2(new_n234), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n359), .B1(new_n803), .B2(new_n374), .C1(new_n793), .C2(new_n203), .ZN(new_n1050));
  AOI211_X1 g0850(.A(new_n1049), .B(new_n1050), .C1(G159), .C2(new_n816), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n807), .A2(G150), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n409), .ZN(new_n1053));
  AOI22_X1  g0853(.A1(new_n795), .A2(new_n1053), .B1(new_n848), .B2(G50), .ZN(new_n1054));
  AND4_X1   g0854(.A1(new_n1026), .A2(new_n1051), .A3(new_n1052), .A4(new_n1054), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n792), .A2(G303), .B1(new_n816), .B2(G322), .ZN(new_n1056));
  INV_X1    g0856(.A(G317), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n1056), .B1(new_n818), .B2(new_n810), .C1(new_n784), .C2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT48), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n844), .B2(new_n803), .C1(new_n809), .C2(new_n800), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT49), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n488), .B1(new_n788), .B2(new_n505), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(new_n807), .B2(G326), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1055), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n826), .B(new_n1048), .C1(new_n1064), .C2(new_n865), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1041), .B1(new_n1065), .B2(KEYINPUT114), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n1066), .B1(KEYINPUT114), .B2(new_n1065), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n1040), .B(new_n1067), .C1(new_n824), .C2(new_n989), .ZN(G393));
  NAND2_X1  g0868(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1037), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1070), .A2(new_n727), .A3(new_n1004), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1002), .A2(new_n825), .A3(new_n1003), .ZN(new_n1072));
  OR2_X1    g0872(.A1(new_n966), .A2(new_n827), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n810), .A2(new_n814), .B1(new_n505), .B2(new_n803), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n359), .B1(new_n1074), .B2(KEYINPUT115), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1075), .B1(KEYINPUT115), .B2(new_n1074), .C1(new_n844), .C2(new_n800), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n790), .B1(new_n809), .B2(new_n793), .C1(new_n776), .C2(new_n820), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n818), .A2(new_n783), .B1(new_n786), .B2(new_n1057), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n1078), .B(KEYINPUT52), .Z(new_n1079));
  NOR3_X1   g0879(.A1(new_n1076), .A2(new_n1077), .A3(new_n1079), .ZN(new_n1080));
  OAI22_X1  g0880(.A1(new_n345), .A2(new_n786), .B1(new_n783), .B2(new_n777), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT51), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n488), .B1(new_n795), .B2(G50), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n803), .A2(new_n234), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n792), .B2(new_n371), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .A4(new_n843), .ZN(new_n1087));
  INV_X1    g0887(.A(G143), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n776), .A2(new_n1088), .B1(new_n1082), .B2(new_n1081), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n1087), .B(new_n1089), .C1(G68), .C2(new_n801), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n763), .B1(new_n1080), .B2(new_n1090), .ZN(new_n1091));
  OAI221_X1 g0891(.A(new_n767), .B1(new_n206), .B2(new_n216), .C1(new_n1009), .C2(new_n257), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1073), .A2(new_n826), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n1071), .A2(new_n1072), .A3(new_n1093), .ZN(G390));
  INV_X1    g0894(.A(new_n948), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n942), .B1(new_n946), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n938), .A2(new_n940), .A3(new_n1096), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n945), .B1(new_n736), .B2(new_n842), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n921), .B(new_n942), .C1(new_n1095), .C2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1097), .A2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n887), .A2(G330), .A3(new_n842), .A4(new_n948), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n1101), .A2(KEYINPUT116), .ZN(new_n1102));
  INV_X1    g0902(.A(KEYINPUT116), .ZN(new_n1103));
  NAND4_X1  g0903(.A1(new_n753), .A2(new_n1103), .A3(new_n842), .A4(new_n948), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1100), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(KEYINPUT117), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1097), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1108));
  INV_X1    g0908(.A(KEYINPUT117), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1100), .A2(new_n1109), .A3(new_n1105), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n887), .A2(G330), .A3(new_n842), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n1095), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1102), .A2(new_n1104), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1101), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n948), .B1(new_n753), .B2(new_n842), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  AOI22_X1  g0917(.A1(new_n1114), .A2(new_n947), .B1(new_n1117), .B2(new_n1098), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n935), .A2(new_n673), .A3(new_n952), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1111), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g0922(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .A4(new_n1120), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n727), .A3(new_n1123), .ZN(new_n1124));
  AND3_X1   g0924(.A1(new_n1107), .A2(new_n1108), .A3(new_n1110), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n941), .A2(new_n764), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n826), .B1(new_n1053), .B2(new_n835), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n802), .A2(new_n488), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n1129), .A2(KEYINPUT118), .B1(G283), .B2(new_n816), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n848), .A2(G116), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT118), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1128), .A2(new_n1132), .B1(G97), .B2(new_n792), .ZN(new_n1133));
  AOI211_X1 g0933(.A(new_n1085), .B(new_n858), .C1(G107), .C2(new_n795), .ZN(new_n1134));
  NAND4_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .A4(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G294), .B2(new_n807), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT119), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n788), .A2(new_n201), .ZN(new_n1138));
  XOR2_X1   g0938(.A(KEYINPUT54), .B(G143), .Z(new_n1139));
  AOI22_X1  g0939(.A1(new_n792), .A2(new_n1139), .B1(G159), .B2(new_n1024), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1140), .B(new_n359), .C1(new_n1141), .C2(new_n786), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1142), .B1(G132), .B2(new_n848), .ZN(new_n1143));
  NOR2_X1   g0943(.A1(new_n800), .A2(new_n345), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1145), .A2(KEYINPUT53), .B1(G137), .B2(new_n795), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT53), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n807), .A2(G125), .B1(new_n1147), .B2(new_n1144), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1143), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1137), .B1(new_n1138), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1127), .B1(new_n1150), .B2(new_n763), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(new_n1125), .A2(new_n825), .B1(new_n1126), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1124), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(KEYINPUT120), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT120), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1124), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1154), .A2(new_n1156), .ZN(G378));
  XNOR2_X1  g0957(.A(new_n431), .B(KEYINPUT121), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n351), .A2(new_n909), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1158), .A2(new_n351), .A3(new_n909), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n1161), .A2(new_n1164), .A3(new_n1162), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n1168), .A2(new_n765), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n201), .B1(new_n267), .B2(G41), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n810), .A2(new_n861), .B1(new_n345), .B2(new_n803), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G125), .A2(new_n816), .B1(new_n848), .B2(G128), .ZN(new_n1172));
  INV_X1    g0972(.A(G137), .ZN(new_n1173));
  OAI21_X1  g0973(.A(new_n1172), .B1(new_n1173), .B2(new_n793), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n1171), .B(new_n1174), .C1(new_n801), .C2(new_n1139), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT59), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G33), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(G41), .B1(new_n807), .B2(G124), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n1177), .B(new_n1178), .C1(new_n777), .C2(new_n788), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1170), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n783), .A2(new_n207), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n792), .A2(new_n373), .ZN(new_n1183));
  AOI21_X1  g0983(.A(G41), .B1(new_n1024), .B2(G68), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n816), .A2(G116), .ZN(new_n1185));
  NAND4_X1  g0985(.A1(new_n1183), .A2(new_n488), .A3(new_n1184), .A4(new_n1185), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n1182), .B(new_n1186), .C1(G97), .C2(new_n795), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1049), .B1(G58), .B2(new_n789), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1187), .B(new_n1188), .C1(new_n844), .C2(new_n776), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT58), .Z(new_n1190));
  OAI21_X1  g0990(.A(new_n763), .B1(new_n1181), .B2(new_n1190), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1191), .B(new_n826), .C1(G50), .C2(new_n835), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n1169), .A2(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n949), .B1(new_n663), .B2(new_n909), .C1(new_n941), .C2(new_n942), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n924), .A2(new_n930), .A3(new_n1168), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1168), .B1(new_n924), .B2(new_n930), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n1194), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1168), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n934), .A2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n924), .A2(new_n1168), .A3(new_n930), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1199), .A2(new_n951), .A3(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1197), .A2(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1193), .B1(new_n1202), .B2(new_n825), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1119), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1201), .A2(new_n1197), .B1(new_n1123), .B2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n727), .B1(new_n1205), .B2(KEYINPUT57), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1123), .A2(new_n1204), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1202), .A2(new_n1207), .A3(KEYINPUT57), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1206), .B2(new_n1209), .ZN(G375));
  AOI21_X1  g1010(.A(new_n869), .B1(new_n1095), .B2(new_n764), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n792), .A2(G150), .B1(G50), .B2(new_n1024), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(KEYINPUT122), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n488), .B1(new_n795), .B2(new_n1139), .ZN(new_n1214));
  OAI211_X1 g1014(.A(new_n1213), .B(new_n1214), .C1(new_n776), .C2(new_n1141), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n853), .A2(G137), .B1(G132), .B2(new_n816), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(KEYINPUT122), .B2(new_n1212), .C1(new_n202), .C2(new_n788), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1215), .B(new_n1217), .C1(G159), .C2(new_n801), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(G107), .A2(new_n792), .B1(new_n795), .B2(G116), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1219), .B(new_n488), .C1(new_n206), .C2(new_n800), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n816), .A2(G294), .B1(new_n373), .B2(new_n1024), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1221), .B1(new_n234), .B2(new_n788), .C1(new_n776), .C2(new_n814), .ZN(new_n1222));
  AOI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(G283), .C2(new_n848), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n763), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1211), .B(new_n1224), .C1(G68), .C2(new_n835), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1118), .B2(new_n824), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1121), .A2(new_n985), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1114), .A2(new_n947), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1117), .A2(new_n1098), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NOR2_X1   g1031(.A1(new_n1204), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1227), .B1(new_n1228), .B2(new_n1232), .ZN(G381));
  INV_X1    g1033(.A(G390), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1033), .A2(new_n1035), .A3(new_n1234), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1235), .A2(G384), .A3(G381), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G375), .A2(new_n1153), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G393), .A2(G396), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1236), .A2(new_n1237), .A3(new_n1238), .ZN(G407));
  NAND2_X1  g1039(.A1(new_n1237), .A2(new_n706), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(G407), .A2(G213), .A3(new_n1240), .ZN(G409));
  XNOR2_X1  g1041(.A(G393), .B(new_n832), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1032), .A2(G390), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1242), .B1(new_n1235), .B2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1234), .A2(new_n1031), .A3(new_n1006), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1243), .A2(new_n1245), .A3(new_n1242), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT61), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT60), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1250), .B1(new_n1204), .B2(new_n1231), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1251), .A2(new_n1121), .A3(new_n727), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1118), .A2(new_n1119), .A3(KEYINPUT60), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1253), .B(KEYINPUT124), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1252), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G384), .B1(new_n1255), .B2(new_n1227), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G384), .ZN(new_n1258));
  AOI211_X1 g1058(.A(new_n1258), .B(new_n1226), .C1(new_n1252), .C2(new_n1254), .ZN(new_n1259));
  INV_X1    g1059(.A(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(G213), .ZN(new_n1261));
  NOR2_X1   g1061(.A1(new_n1261), .A2(G343), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(G2897), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1257), .A2(new_n1260), .A3(new_n1263), .ZN(new_n1264));
  OAI211_X1 g1064(.A(G2897), .B(new_n1262), .C1(new_n1256), .C2(new_n1259), .ZN(new_n1265));
  AND2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1203), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1202), .A2(new_n1207), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT57), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1038), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1267), .B1(new_n1270), .B2(new_n1208), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1202), .A2(new_n1207), .A3(new_n985), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT123), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1205), .A2(KEYINPUT123), .A3(new_n985), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1274), .A2(new_n1275), .A3(new_n1203), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1153), .ZN(new_n1277));
  AOI22_X1  g1077(.A1(new_n1271), .A2(G378), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1266), .B1(new_n1278), .B2(new_n1262), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1257), .A2(new_n1260), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1281), .A2(new_n727), .A3(new_n1208), .ZN(new_n1282));
  AOI21_X1  g1082(.A(new_n1155), .B1(new_n1124), .B2(new_n1152), .ZN(new_n1283));
  AND3_X1   g1083(.A1(new_n1124), .A2(new_n1152), .A3(new_n1155), .ZN(new_n1284));
  OAI211_X1 g1084(.A(new_n1282), .B(new_n1203), .C1(new_n1283), .C2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1286));
  AOI211_X1 g1086(.A(new_n1262), .B(new_n1280), .C1(new_n1285), .C2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT62), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1249), .B(new_n1279), .C1(new_n1287), .C2(new_n1288), .ZN(new_n1289));
  INV_X1    g1089(.A(new_n1262), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1280), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1284), .A2(new_n1283), .ZN(new_n1292));
  NOR2_X1   g1092(.A1(new_n1292), .A2(G375), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1276), .A2(new_n1277), .ZN(new_n1294));
  OAI211_X1 g1094(.A(new_n1290), .B(new_n1291), .C1(new_n1293), .C2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1295), .A2(KEYINPUT62), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1248), .B1(new_n1289), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT125), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT63), .B1(new_n1287), .B2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n1242), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1035), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1034), .B1(new_n1006), .B2(new_n1031), .ZN(new_n1302));
  NOR3_X1   g1102(.A1(new_n1301), .A2(new_n1302), .A3(G390), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1243), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1300), .B1(new_n1303), .B2(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1246), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1290), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1307));
  AOI21_X1  g1107(.A(KEYINPUT61), .B1(new_n1307), .B2(new_n1266), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT63), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1295), .A2(KEYINPUT125), .A3(new_n1309), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1299), .A2(new_n1306), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1297), .A2(new_n1311), .ZN(G405));
  NAND2_X1  g1112(.A1(G375), .A2(new_n1277), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1285), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT126), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1291), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  AOI211_X1 g1116(.A(KEYINPUT126), .B(new_n1280), .C1(new_n1285), .C2(new_n1313), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(new_n1316), .A2(new_n1317), .ZN(new_n1318));
  INV_X1    g1118(.A(KEYINPUT127), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1285), .A2(new_n1313), .A3(KEYINPUT126), .ZN(new_n1320));
  NAND4_X1  g1120(.A1(new_n1318), .A2(new_n1306), .A3(new_n1319), .A4(new_n1320), .ZN(new_n1321));
  AOI21_X1  g1121(.A(new_n1153), .B1(new_n1282), .B2(new_n1203), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1315), .B1(new_n1293), .B2(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1323), .A2(new_n1280), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1314), .A2(new_n1315), .A3(new_n1291), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1324), .A2(new_n1320), .A3(new_n1325), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1305), .A2(KEYINPUT127), .A3(new_n1246), .ZN(new_n1327));
  OAI21_X1  g1127(.A(new_n1319), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1326), .A2(new_n1327), .A3(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1321), .A2(new_n1329), .ZN(G402));
endmodule


