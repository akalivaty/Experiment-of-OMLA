//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 0 0 0 0 1 0 0 1 1 1 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 1 0 0 1 0 0 0 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n437, new_n447, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n460, new_n461, new_n462, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n570, new_n571, new_n573, new_n574, new_n575,
    new_n576, new_n577, new_n578, new_n579, new_n580, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n615, new_n616,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1203;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n437));
  XNOR2_X1  g012(.A(new_n436), .B(new_n437), .ZN(G220));
  INV_X1    g013(.A(G96), .ZN(G221));
  INV_X1    g014(.A(G69), .ZN(G235));
  INV_X1    g015(.A(G120), .ZN(G236));
  INV_X1    g016(.A(G57), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XOR2_X1   g028(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  INV_X1    g033(.A(G325), .ZN(G261));
  NAND2_X1  g034(.A1(new_n455), .A2(G2106), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n457), .A2(G567), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(G319));
  INV_X1    g038(.A(G101), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT67), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n465), .B1(G2104), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR3_X1   g043(.A1(new_n468), .A2(KEYINPUT67), .A3(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  INV_X1    g047(.A(G137), .ZN(new_n473));
  OAI22_X1  g048(.A1(new_n464), .A2(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n466), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n474), .A2(new_n477), .ZN(G160));
  INV_X1    g053(.A(new_n472), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n471), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G124), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n466), .A2(G112), .ZN(new_n484));
  OAI21_X1  g059(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n480), .B(new_n483), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT68), .ZN(G162));
  OAI21_X1  g062(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  AOI21_X1  g064(.A(new_n488), .B1(new_n489), .B2(G2105), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n471), .A2(G138), .A3(new_n466), .ZN(new_n491));
  NAND2_X1  g066(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n471), .A2(G138), .A3(new_n466), .A4(new_n492), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT69), .ZN(new_n497));
  INV_X1    g072(.A(G126), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n481), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g074(.A1(new_n471), .A2(KEYINPUT69), .A3(G126), .A4(G2105), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT5), .B(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  AND3_X1   g082(.A1(new_n507), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n508));
  AOI21_X1  g083(.A(KEYINPUT71), .B1(new_n507), .B2(KEYINPUT6), .ZN(new_n509));
  OAI211_X1 g084(.A(new_n504), .B(new_n506), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT72), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT71), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n505), .B2(G651), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n507), .A2(KEYINPUT71), .A3(KEYINPUT6), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g091(.A1(new_n516), .A2(KEYINPUT72), .A3(new_n504), .A4(new_n506), .ZN(new_n517));
  AND2_X1   g092(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n516), .A2(G543), .A3(new_n506), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(G75), .A2(G543), .ZN(new_n522));
  OR2_X1    g097(.A1(KEYINPUT5), .A2(G543), .ZN(new_n523));
  NAND2_X1  g098(.A1(KEYINPUT5), .A2(G543), .ZN(new_n524));
  AND2_X1   g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n522), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g102(.A1(new_n521), .A2(G50), .B1(new_n527), .B2(G651), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n519), .A2(new_n528), .ZN(G303));
  INV_X1    g104(.A(G303), .ZN(G166));
  NAND2_X1  g105(.A1(new_n521), .A2(G51), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n504), .A2(KEYINPUT73), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT73), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n523), .A2(new_n533), .A3(new_n524), .ZN(new_n534));
  NAND4_X1  g109(.A1(new_n532), .A2(G63), .A3(G651), .A4(new_n534), .ZN(new_n535));
  XOR2_X1   g110(.A(KEYINPUT74), .B(KEYINPUT7), .Z(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n531), .A2(new_n535), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n518), .A2(G89), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n539), .A2(new_n540), .ZN(G286));
  INV_X1    g116(.A(G286), .ZN(G168));
  NAND2_X1  g117(.A1(new_n518), .A2(G90), .ZN(new_n543));
  NAND2_X1  g118(.A1(G77), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n532), .A2(new_n534), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g122(.A1(new_n547), .A2(G651), .B1(G52), .B2(new_n521), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n543), .A2(new_n548), .ZN(G301));
  INV_X1    g124(.A(G301), .ZN(G171));
  NAND3_X1  g125(.A1(new_n532), .A2(G56), .A3(new_n534), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(KEYINPUT75), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT75), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n551), .A2(new_n555), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n554), .A2(G651), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n512), .A2(G81), .A3(new_n517), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n521), .A2(G43), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n558), .A2(KEYINPUT76), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT76), .B1(new_n558), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g136(.A(new_n557), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  OAI211_X1 g139(.A(KEYINPUT77), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n567), .A2(G860), .ZN(G153));
  NAND4_X1  g143(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  NAND2_X1  g147(.A1(new_n518), .A2(G91), .ZN(new_n573));
  INV_X1    g148(.A(G53), .ZN(new_n574));
  OR3_X1    g149(.A1(new_n520), .A2(KEYINPUT9), .A3(new_n574), .ZN(new_n575));
  OAI21_X1  g150(.A(KEYINPUT9), .B1(new_n520), .B2(new_n574), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g152(.A1(new_n504), .A2(G65), .ZN(new_n578));
  AND2_X1   g153(.A1(G78), .A2(G543), .ZN(new_n579));
  OAI21_X1  g154(.A(G651), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n573), .A2(new_n577), .A3(new_n580), .ZN(G299));
  AND2_X1   g156(.A1(G49), .A2(G543), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n516), .A2(new_n506), .A3(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n583), .B(new_n584), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n512), .A2(G87), .A3(new_n517), .ZN(new_n586));
  AND2_X1   g161(.A1(new_n532), .A2(new_n534), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n587), .B2(G74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n585), .A2(new_n586), .A3(new_n588), .ZN(G288));
  NAND2_X1  g164(.A1(G73), .A2(G543), .ZN(new_n590));
  INV_X1    g165(.A(G61), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n525), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n521), .A2(G48), .B1(new_n592), .B2(G651), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n512), .A2(G86), .A3(new_n517), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(G305));
  NAND2_X1  g170(.A1(G72), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G60), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n545), .B2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT79), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n507), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(new_n599), .B2(new_n598), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n518), .A2(G85), .B1(G47), .B2(new_n521), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n601), .A2(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n521), .A2(G54), .ZN(new_n605));
  AOI22_X1  g180(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n507), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n518), .A2(G92), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n518), .A2(KEYINPUT10), .A3(G92), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n604), .B1(new_n612), .B2(G868), .ZN(G284));
  OAI21_X1  g188(.A(new_n604), .B1(new_n612), .B2(G868), .ZN(G321));
  NAND2_X1  g189(.A1(G286), .A2(G868), .ZN(new_n615));
  INV_X1    g190(.A(G299), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G297));
  OAI21_X1  g192(.A(new_n615), .B1(new_n616), .B2(G868), .ZN(G280));
  INV_X1    g193(.A(G559), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(G860), .ZN(G148));
  INV_X1    g195(.A(G868), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n566), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n612), .A2(new_n619), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT80), .Z(new_n624));
  OAI21_X1  g199(.A(new_n622), .B1(new_n624), .B2(new_n621), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n470), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(new_n471), .ZN(new_n628));
  XNOR2_X1  g203(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(KEYINPUT13), .Z(new_n631));
  OR2_X1    g206(.A1(new_n631), .A2(G2100), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n631), .A2(G2100), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n479), .A2(G135), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT82), .Z(new_n635));
  OAI21_X1  g210(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n636));
  INV_X1    g211(.A(G111), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n636), .B1(new_n637), .B2(G2105), .ZN(new_n638));
  AOI21_X1  g213(.A(new_n638), .B1(new_n482), .B2(G123), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n635), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2096), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n632), .A2(new_n633), .A3(new_n641), .ZN(G156));
  XOR2_X1   g217(.A(KEYINPUT15), .B(G2435), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g221(.A(KEYINPUT84), .B(KEYINPUT14), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n645), .ZN(new_n648));
  NAND3_X1  g223(.A1(new_n646), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2451), .B(G2454), .Z(new_n654));
  XNOR2_X1  g229(.A(G2443), .B(G2446), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  OR2_X1    g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n653), .A2(new_n656), .ZN(new_n658));
  AND3_X1   g233(.A1(new_n657), .A2(G14), .A3(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT85), .Z(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT17), .ZN(new_n662));
  XNOR2_X1  g237(.A(G2084), .B(G2090), .ZN(new_n663));
  XNOR2_X1  g238(.A(G2067), .B(G2678), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT87), .ZN(new_n666));
  INV_X1    g241(.A(new_n664), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n667), .A2(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n662), .A2(new_n664), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n672), .B(new_n663), .C1(new_n661), .C2(new_n664), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n666), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2096), .B(G2100), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(G1971), .B(G1976), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(KEYINPUT19), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n679), .A2(new_n680), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n683), .A2(new_n681), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n683), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT88), .B(KEYINPUT20), .Z(new_n686));
  OAI221_X1 g261(.A(new_n682), .B1(new_n684), .B2(new_n678), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n687), .B1(new_n685), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(new_n690));
  XNOR2_X1  g265(.A(G1991), .B(G1996), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XOR2_X1   g267(.A(G1981), .B(G1986), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G229));
  INV_X1    g269(.A(G29), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(G26), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT28), .Z(new_n697));
  NAND2_X1  g272(.A1(new_n479), .A2(G140), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n482), .A2(G128), .ZN(new_n699));
  NOR2_X1   g274(.A1(new_n466), .A2(G116), .ZN(new_n700));
  OAI21_X1  g275(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n698), .B(new_n699), .C1(new_n700), .C2(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n697), .B1(new_n702), .B2(G29), .ZN(new_n703));
  INV_X1    g278(.A(G2067), .ZN(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  XNOR2_X1  g280(.A(KEYINPUT31), .B(G11), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT30), .B(G28), .Z(new_n707));
  OAI21_X1  g282(.A(new_n706), .B1(new_n707), .B2(G29), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n640), .B2(G29), .ZN(new_n709));
  AOI22_X1  g284(.A1(G105), .A2(new_n627), .B1(new_n479), .B2(G141), .ZN(new_n710));
  NAND3_X1  g285(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT26), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(new_n482), .B2(G129), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G32), .B(new_n714), .S(G29), .Z(new_n715));
  XOR2_X1   g290(.A(KEYINPUT27), .B(G1996), .Z(new_n716));
  OAI21_X1  g291(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n705), .B(new_n717), .C1(new_n715), .C2(new_n716), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT24), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n695), .B1(new_n719), .B2(G34), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(new_n719), .B2(G34), .ZN(new_n721));
  AOI21_X1  g296(.A(new_n721), .B1(G160), .B2(G29), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(G2084), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT98), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(G2084), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT94), .Z(new_n726));
  NOR2_X1   g301(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n695), .A2(G33), .ZN(new_n728));
  NAND3_X1  g303(.A1(new_n466), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT92), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT25), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n479), .A2(G139), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n731), .B(new_n732), .C1(new_n466), .C2(new_n733), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n728), .B1(new_n734), .B2(G29), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT93), .ZN(new_n738));
  INV_X1    g313(.A(G16), .ZN(new_n739));
  NOR2_X1   g314(.A1(G171), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G5), .B2(new_n739), .ZN(new_n741));
  INV_X1    g316(.A(G1961), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND4_X1  g318(.A1(new_n718), .A2(new_n727), .A3(new_n738), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n739), .A2(G20), .ZN(new_n745));
  XOR2_X1   g320(.A(new_n745), .B(KEYINPUT23), .Z(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G299), .B2(G16), .ZN(new_n747));
  INV_X1    g322(.A(G1956), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n735), .A2(new_n736), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n695), .A2(G27), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G164), .B2(new_n695), .ZN(new_n753));
  INV_X1    g328(.A(G2078), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  OAI211_X1 g330(.A(new_n751), .B(new_n755), .C1(new_n742), .C2(new_n741), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n744), .A2(new_n749), .A3(new_n756), .ZN(new_n757));
  NOR2_X1   g332(.A1(G286), .A2(new_n739), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(KEYINPUT96), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT96), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G16), .B2(G21), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(new_n758), .B2(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(G1966), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT97), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n739), .A2(G4), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n765), .B1(new_n612), .B2(new_n739), .ZN(new_n766));
  INV_X1    g341(.A(G1348), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n762), .A2(G1966), .ZN(new_n769));
  NOR2_X1   g344(.A1(G29), .A2(G35), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G162), .B2(G29), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(KEYINPUT29), .Z(new_n772));
  INV_X1    g347(.A(G2090), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n769), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n774), .B1(new_n773), .B2(new_n772), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n757), .A2(new_n764), .A3(new_n768), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n739), .A2(G19), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n567), .B2(new_n739), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1341), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  AND2_X1   g356(.A1(new_n739), .A2(G22), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G303), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT90), .ZN(new_n784));
  OR2_X1    g359(.A1(new_n784), .A2(G1971), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(G1971), .ZN(new_n786));
  NOR2_X1   g361(.A1(G6), .A2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G305), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(G16), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT32), .B(G1981), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n785), .A2(new_n786), .A3(new_n791), .ZN(new_n792));
  AND2_X1   g367(.A1(new_n739), .A2(G23), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G288), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT33), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n794), .A2(new_n795), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G1976), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  NOR3_X1   g375(.A1(new_n792), .A2(KEYINPUT34), .A3(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(KEYINPUT91), .ZN(new_n803));
  INV_X1    g378(.A(G290), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(G16), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G16), .B2(G24), .ZN(new_n806));
  INV_X1    g381(.A(G1986), .ZN(new_n807));
  AND2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NOR2_X1   g384(.A1(G25), .A2(G29), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n479), .A2(G131), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n482), .A2(G119), .ZN(new_n812));
  OR2_X1    g387(.A1(G95), .A2(G2105), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n813), .B(G2104), .C1(G107), .C2(new_n466), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n811), .A2(new_n812), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n810), .B1(new_n816), .B2(G29), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT35), .B(G1991), .Z(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT89), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n817), .B(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n808), .A2(new_n809), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n802), .A2(new_n803), .A3(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(new_n821), .ZN(new_n823));
  OAI21_X1  g398(.A(KEYINPUT91), .B1(new_n801), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(KEYINPUT34), .B1(new_n792), .B2(new_n800), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n827), .A2(KEYINPUT36), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT36), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n825), .A2(new_n829), .A3(new_n826), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n781), .B1(new_n828), .B2(new_n830), .ZN(G311));
  NAND2_X1  g406(.A1(new_n828), .A2(new_n830), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(new_n780), .ZN(G150));
  NAND2_X1  g408(.A1(G80), .A2(G543), .ZN(new_n834));
  INV_X1    g409(.A(G67), .ZN(new_n835));
  OAI21_X1  g410(.A(new_n834), .B1(new_n545), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n836), .A2(G651), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n512), .A2(G93), .A3(new_n517), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n521), .A2(G55), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT37), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n612), .A2(G559), .ZN(new_n844));
  XOR2_X1   g419(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n840), .B(new_n557), .C1(new_n560), .C2(new_n561), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(new_n840), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n848), .B1(new_n566), .B2(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n846), .B(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(KEYINPUT39), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n841), .B1(new_n852), .B2(KEYINPUT39), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n843), .B1(new_n853), .B2(new_n854), .ZN(G145));
  XOR2_X1   g430(.A(G162), .B(G160), .Z(new_n856));
  XOR2_X1   g431(.A(new_n856), .B(new_n640), .Z(new_n857));
  INV_X1    g432(.A(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n859));
  AND3_X1   g434(.A1(new_n496), .A2(new_n859), .A3(new_n501), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n859), .B1(new_n496), .B2(new_n501), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n862), .B(new_n702), .Z(new_n863));
  XNOR2_X1  g438(.A(new_n863), .B(new_n714), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n734), .B2(KEYINPUT102), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n482), .A2(G130), .ZN(new_n869));
  NOR2_X1   g444(.A1(new_n466), .A2(G118), .ZN(new_n870));
  OAI21_X1  g445(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n872), .B1(G142), .B2(new_n479), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(new_n816), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(new_n630), .Z(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n867), .B1(new_n866), .B2(new_n734), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n864), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n868), .A2(new_n876), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g455(.A(new_n876), .B1(new_n868), .B2(new_n878), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n858), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(new_n857), .A3(new_n879), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n882), .A2(new_n884), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n886), .B(new_n887), .ZN(G395));
  XNOR2_X1  g463(.A(new_n624), .B(new_n850), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n610), .A2(new_n611), .ZN(new_n890));
  INV_X1    g465(.A(new_n607), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n892), .A2(G299), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n612), .A2(new_n616), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n895), .A2(KEYINPUT41), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n893), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n889), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(new_n895), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n889), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(G290), .A2(G166), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n601), .A2(G303), .A3(new_n602), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n788), .A2(G288), .ZN(new_n906));
  INV_X1    g481(.A(G288), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n907), .A2(G305), .ZN(new_n908));
  AND4_X1   g483(.A1(new_n904), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n904), .A2(new_n905), .B1(new_n906), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n911), .B(KEYINPUT42), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n901), .A2(new_n903), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n913), .B1(new_n901), .B2(new_n903), .ZN(new_n915));
  OAI21_X1  g490(.A(G868), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n916), .B1(G868), .B2(new_n840), .ZN(G295));
  OAI21_X1  g492(.A(new_n916), .B1(G868), .B2(new_n840), .ZN(G331));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n558), .A2(new_n559), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT76), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n558), .A2(KEYINPUT76), .A3(new_n559), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(KEYINPUT77), .B1(new_n924), .B2(new_n557), .ZN(new_n925));
  INV_X1    g500(.A(new_n565), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n849), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G286), .A2(G301), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n540), .A2(new_n539), .A3(new_n543), .A4(new_n548), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n847), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n840), .B1(new_n564), .B2(new_n565), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n930), .B1(new_n933), .B2(new_n848), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n911), .B1(new_n935), .B2(new_n899), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  OAI211_X1 g513(.A(KEYINPUT104), .B(new_n930), .C1(new_n933), .C2(new_n848), .ZN(new_n939));
  AOI21_X1  g514(.A(KEYINPUT105), .B1(new_n850), .B2(new_n931), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT105), .ZN(new_n941));
  NOR4_X1   g516(.A1(new_n933), .A2(new_n941), .A3(new_n930), .A4(new_n848), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n938), .B(new_n939), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n919), .B(new_n936), .C1(new_n943), .C2(new_n895), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n932), .A2(new_n941), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n850), .A2(KEYINPUT105), .A3(new_n931), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n948), .A2(new_n902), .A3(new_n938), .A4(new_n939), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n919), .B1(new_n949), .B2(new_n936), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n945), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT43), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n902), .A2(KEYINPUT107), .A3(new_n897), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n898), .A2(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n953), .A2(new_n896), .A3(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n935), .ZN(new_n957));
  AOI22_X1  g532(.A1(new_n943), .A2(new_n956), .B1(new_n957), .B2(new_n902), .ZN(new_n958));
  INV_X1    g533(.A(new_n911), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n885), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n951), .A2(new_n952), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n936), .B1(new_n943), .B2(new_n895), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(new_n944), .ZN(new_n964));
  OAI22_X1  g539(.A1(new_n943), .A2(new_n895), .B1(new_n900), .B2(new_n957), .ZN(new_n965));
  AOI21_X1  g540(.A(G37), .B1(new_n965), .B2(new_n911), .ZN(new_n966));
  AOI21_X1  g541(.A(KEYINPUT43), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  NOR3_X1   g544(.A1(new_n951), .A2(KEYINPUT43), .A3(new_n960), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n952), .B1(new_n964), .B2(new_n966), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n968), .A2(new_n972), .ZN(G397));
  NAND2_X1  g548(.A1(new_n804), .A2(new_n807), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n974), .B(KEYINPUT108), .ZN(new_n975));
  INV_X1    g550(.A(G1996), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n714), .B(new_n976), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n702), .B(new_n704), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n816), .A2(new_n818), .ZN(new_n979));
  OR2_X1    g554(.A1(new_n816), .A2(new_n818), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n977), .A2(new_n978), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n981), .B1(G1986), .B2(G290), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n975), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(G1384), .ZN(new_n984));
  AOI21_X1  g559(.A(KEYINPUT45), .B1(new_n862), .B2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G40), .ZN(new_n986));
  NOR3_X1   g561(.A1(new_n474), .A2(new_n477), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n983), .A2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT54), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n496), .B2(new_n501), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n987), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  AOI211_X1 g569(.A(KEYINPUT50), .B(G1384), .C1(new_n496), .C2(new_n501), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  XOR2_X1   g571(.A(KEYINPUT123), .B(G1961), .Z(new_n997));
  NOR2_X1   g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n987), .A2(KEYINPUT53), .A3(new_n754), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n985), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n502), .A2(KEYINPUT100), .ZN(new_n1001));
  NAND3_X1  g576(.A1(new_n496), .A2(new_n859), .A3(new_n501), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(G1384), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1001), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1005), .A2(KEYINPUT109), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT109), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n1001), .A2(new_n1007), .A3(new_n1002), .A4(new_n1004), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n998), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT124), .B(KEYINPUT53), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n987), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n1012), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1013));
  AOI211_X1 g588(.A(KEYINPUT125), .B(new_n1011), .C1(new_n1013), .C2(new_n754), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT125), .ZN(new_n1015));
  INV_X1    g590(.A(new_n987), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n502), .A2(new_n984), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1016), .B1(new_n1017), .B2(new_n1003), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1007), .B1(new_n862), .B2(new_n1004), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1008), .ZN(new_n1020));
  OAI211_X1 g595(.A(new_n754), .B(new_n1018), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(new_n1011), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1015), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  OAI211_X1 g598(.A(G301), .B(new_n1010), .C1(new_n1014), .C2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT126), .ZN(new_n1025));
  INV_X1    g600(.A(new_n998), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n502), .A2(new_n1004), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1018), .A2(KEYINPUT53), .A3(new_n754), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  AOI211_X1 g604(.A(G2078), .B(new_n1012), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT125), .B1(new_n1030), .B2(new_n1011), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1021), .A2(new_n1015), .A3(new_n1022), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI22_X1  g608(.A1(new_n1024), .A2(new_n1025), .B1(new_n1033), .B2(G301), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1010), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1035), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT126), .B1(new_n1036), .B2(G301), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n991), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G1966), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1027), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1039), .B1(new_n1012), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1017), .A2(KEYINPUT50), .ZN(new_n1042));
  INV_X1    g617(.A(G2084), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n502), .A2(new_n993), .A3(new_n984), .ZN(new_n1044));
  NAND4_X1  g619(.A1(new_n1042), .A2(new_n1043), .A3(new_n987), .A4(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1041), .A2(new_n1045), .A3(G168), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1046), .A2(G8), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT51), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1966), .B1(new_n1018), .B2(new_n1027), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n994), .A2(G2084), .A3(new_n995), .ZN(new_n1051));
  OAI21_X1  g626(.A(G286), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(G8), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n1052), .A2(new_n1046), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(G303), .A2(G8), .ZN(new_n1058));
  XNOR2_X1  g633(.A(new_n1058), .B(KEYINPUT55), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1016), .B1(new_n1017), .B2(KEYINPUT50), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1044), .A2(KEYINPUT114), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n992), .B2(new_n993), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n773), .B(new_n1060), .C1(new_n1061), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(G1971), .ZN(new_n1066));
  OAI21_X1  g641(.A(new_n1018), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1059), .B1(new_n1068), .B2(new_n1053), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1059), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1013), .A2(G1971), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n996), .A2(new_n773), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1072), .ZN(new_n1073));
  OAI211_X1 g648(.A(G8), .B(new_n1070), .C1(new_n1071), .C2(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n502), .A2(new_n987), .A3(new_n984), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1075), .A2(G8), .ZN(new_n1076));
  XNOR2_X1  g651(.A(KEYINPUT111), .B(G1981), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n788), .A2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT112), .ZN(new_n1079));
  AND3_X1   g654(.A1(G305), .A2(new_n1079), .A3(G1981), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1079), .B1(G305), .B2(G1981), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1078), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT49), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1076), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  OAI211_X1 g659(.A(KEYINPUT49), .B(new_n1078), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n585), .A2(new_n588), .A3(G1976), .A4(new_n586), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1075), .A2(G8), .A3(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(KEYINPUT52), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT110), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(KEYINPUT110), .A3(KEYINPUT52), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1088), .ZN(new_n1093));
  AOI21_X1  g668(.A(KEYINPUT52), .B1(G288), .B2(new_n799), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1091), .A2(new_n1092), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1086), .A2(new_n1095), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1057), .A2(new_n1069), .A3(new_n1074), .A4(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1010), .B1(new_n1014), .B2(new_n1023), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n991), .B1(new_n1098), .B2(G171), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1033), .A2(G301), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1097), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1038), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(new_n736), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1018), .B(new_n1104), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1060), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(new_n748), .ZN(new_n1107));
  XOR2_X1   g682(.A(G299), .B(KEYINPUT57), .Z(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(KEYINPUT121), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1105), .A2(new_n1112), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1111), .A2(new_n1113), .A3(KEYINPUT61), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n767), .B1(new_n994), .B2(new_n995), .ZN(new_n1115));
  INV_X1    g690(.A(new_n1075), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n704), .ZN(new_n1117));
  AOI21_X1  g692(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(KEYINPUT60), .A3(new_n1117), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n612), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1115), .A2(new_n892), .A3(KEYINPUT60), .A4(new_n1117), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT59), .ZN(new_n1123));
  AOI211_X1 g698(.A(G1996), .B(new_n1012), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1124));
  XOR2_X1   g699(.A(KEYINPUT119), .B(KEYINPUT58), .Z(new_n1125));
  XNOR2_X1  g700(.A(new_n1125), .B(G1341), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1116), .A2(new_n1126), .ZN(new_n1127));
  OAI221_X1 g702(.A(new_n567), .B1(KEYINPUT120), .B2(new_n1123), .C1(new_n1124), .C2(new_n1127), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1123), .A2(KEYINPUT120), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1127), .B1(new_n1013), .B2(new_n976), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1129), .B1(new_n1130), .B2(new_n566), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1122), .B1(new_n1128), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1109), .A2(KEYINPUT118), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT61), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT118), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1105), .A2(new_n1108), .A3(new_n1107), .A4(new_n1135), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1133), .A2(new_n1134), .A3(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1114), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT122), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n892), .B1(new_n1117), .B2(new_n1115), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1140), .B1(new_n1110), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1138), .A2(new_n1139), .A3(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1139), .B1(new_n1138), .B2(new_n1142), .ZN(new_n1144));
  NOR3_X1   g719(.A1(new_n1102), .A2(new_n1143), .A3(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1086), .A2(new_n1095), .A3(KEYINPUT113), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT113), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1067), .A2(new_n1066), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1053), .B1(new_n1148), .B2(new_n1072), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1146), .A2(new_n1147), .B1(new_n1070), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT116), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI221_X1 g727(.A(KEYINPUT116), .B1(new_n1149), .B2(new_n1070), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1153));
  AOI211_X1 g728(.A(new_n1053), .B(G286), .C1(new_n1041), .C2(new_n1045), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n1074), .A2(KEYINPUT63), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1152), .A2(new_n1153), .A3(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1069), .A2(new_n1074), .A3(new_n1096), .A4(new_n1154), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT115), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1157), .A2(KEYINPUT115), .A3(new_n1158), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1156), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1164));
  OAI211_X1 g739(.A(new_n1026), .B(new_n1028), .C1(new_n1014), .C2(new_n1023), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT62), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1049), .A2(new_n1055), .A3(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1166), .B1(new_n1049), .B2(new_n1055), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(G171), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1069), .A2(new_n1074), .A3(new_n1096), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1164), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1170), .ZN(new_n1172));
  INV_X1    g747(.A(new_n1168), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1049), .A2(new_n1055), .A3(new_n1166), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1033), .A2(G301), .ZN(new_n1176));
  NAND4_X1  g751(.A1(new_n1172), .A2(new_n1175), .A3(new_n1176), .A4(KEYINPUT127), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1086), .A2(new_n799), .A3(new_n907), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1076), .B1(new_n1179), .B2(new_n1078), .ZN(new_n1180));
  OR2_X1    g755(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1181));
  INV_X1    g756(.A(new_n1074), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1180), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1163), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n990), .B1(new_n1145), .B2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n975), .A2(new_n988), .ZN(new_n1186));
  OR2_X1    g761(.A1(new_n1186), .A2(KEYINPUT48), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(KEYINPUT48), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n989), .A2(new_n981), .ZN(new_n1189));
  NAND3_X1  g764(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n977), .A2(new_n978), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1191), .A2(new_n979), .B1(G2067), .B2(new_n702), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n989), .A2(new_n1192), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n988), .A2(G1996), .ZN(new_n1194));
  NOR2_X1   g769(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1195));
  AND2_X1   g770(.A1(new_n1194), .A2(KEYINPUT46), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n978), .A2(new_n710), .A3(new_n713), .ZN(new_n1197));
  AOI211_X1 g772(.A(new_n1195), .B(new_n1196), .C1(new_n989), .C2(new_n1197), .ZN(new_n1198));
  OAI211_X1 g773(.A(new_n1190), .B(new_n1193), .C1(KEYINPUT47), .C2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g774(.A(new_n1199), .B1(KEYINPUT47), .B2(new_n1198), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1185), .A2(new_n1200), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g776(.A1(G229), .A2(new_n462), .A3(G401), .A4(G227), .ZN(new_n1203));
  OAI211_X1 g777(.A(new_n886), .B(new_n1203), .C1(new_n970), .C2(new_n971), .ZN(G225));
  INV_X1    g778(.A(G225), .ZN(G308));
endmodule


