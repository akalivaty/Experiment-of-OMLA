//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 0 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034;
  INV_X1    g000(.A(KEYINPUT30), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT0), .A4(G128), .ZN(new_n192));
  XNOR2_X1  g006(.A(G143), .B(G146), .ZN(new_n193));
  OR2_X1    g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND2_X1  g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT64), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  INV_X1    g014(.A(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G137), .ZN(new_n202));
  INV_X1    g016(.A(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT11), .A3(G134), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(G137), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G131), .ZN(new_n207));
  INV_X1    g021(.A(G131), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n202), .A2(new_n204), .A3(new_n208), .A4(new_n205), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n207), .A2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT65), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n192), .B(KEYINPUT64), .C1(new_n193), .C2(new_n196), .ZN(new_n212));
  NAND4_X1  g026(.A1(new_n199), .A2(new_n210), .A3(new_n211), .A4(new_n212), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n201), .A2(G137), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n203), .A2(G134), .ZN(new_n215));
  OAI21_X1  g029(.A(G131), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n189), .A2(new_n191), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n218), .A2(KEYINPUT1), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  AOI21_X1  g035(.A(G128), .B1(new_n189), .B2(new_n191), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT1), .ZN(new_n223));
  NOR3_X1   g037(.A1(new_n223), .A2(new_n188), .A3(G143), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n221), .B1(new_n222), .B2(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n188), .A2(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n227), .B(KEYINPUT66), .C1(new_n193), .C2(G128), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n220), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n213), .B1(new_n217), .B2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n212), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n218), .A2(new_n195), .A3(new_n194), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT64), .B1(new_n232), .B2(new_n192), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n211), .B1(new_n234), .B2(new_n210), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n187), .B1(new_n230), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G119), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT67), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT67), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G119), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(new_n240), .A3(G116), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n245), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(new_n241), .A3(new_n243), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n209), .A2(new_n216), .A3(KEYINPUT68), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(KEYINPUT68), .B1(new_n209), .B2(new_n216), .ZN(new_n252));
  NOR3_X1   g066(.A1(new_n229), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n210), .A2(new_n192), .A3(new_n232), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT30), .ZN(new_n255));
  OAI21_X1  g069(.A(KEYINPUT69), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n193), .A2(new_n223), .A3(G128), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n190), .A2(G146), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n219), .B1(new_n258), .B2(new_n226), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT66), .B1(new_n259), .B2(new_n227), .ZN(new_n260));
  NOR3_X1   g074(.A1(new_n222), .A2(new_n221), .A3(new_n224), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n257), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n252), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n262), .A2(new_n250), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n265));
  NAND4_X1  g079(.A1(new_n264), .A2(new_n265), .A3(KEYINPUT30), .A4(new_n254), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n236), .A2(new_n249), .A3(new_n256), .A4(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(new_n249), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n264), .A2(new_n268), .A3(new_n254), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(G237), .ZN(new_n271));
  INV_X1    g085(.A(G953), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(new_n272), .A3(G210), .ZN(new_n273));
  XOR2_X1   g087(.A(new_n273), .B(KEYINPUT27), .Z(new_n274));
  XNOR2_X1  g088(.A(KEYINPUT26), .B(G101), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n267), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT31), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n277), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n269), .A2(KEYINPUT28), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n197), .B1(new_n209), .B2(new_n207), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n225), .A2(new_n228), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n252), .B1(new_n284), .B2(new_n257), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n285), .B2(new_n250), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT28), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(new_n268), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n199), .A2(new_n210), .A3(new_n212), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(KEYINPUT65), .ZN(new_n290));
  OAI211_X1 g104(.A(new_n290), .B(new_n213), .C1(new_n217), .C2(new_n229), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n282), .A2(new_n288), .B1(new_n249), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n276), .ZN(new_n293));
  OAI21_X1  g107(.A(KEYINPUT70), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n249), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n287), .B1(new_n286), .B2(new_n268), .ZN(new_n296));
  NOR4_X1   g110(.A1(new_n253), .A2(KEYINPUT28), .A3(new_n283), .A4(new_n249), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT70), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n298), .A2(new_n299), .A3(new_n276), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n280), .A2(new_n281), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(G472), .A2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT71), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n299), .B1(new_n298), .B2(new_n276), .ZN(new_n306));
  NOR3_X1   g120(.A1(new_n292), .A2(KEYINPUT70), .A3(new_n293), .ZN(new_n307));
  AND3_X1   g121(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n277), .ZN(new_n308));
  AOI21_X1  g122(.A(KEYINPUT31), .B1(new_n267), .B2(new_n277), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n306), .A2(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT71), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n311), .A3(new_n302), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(new_n305), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n280), .A2(new_n281), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n294), .A2(new_n300), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n303), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(G902), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n264), .A2(new_n254), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(new_n249), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n296), .B2(new_n297), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n293), .A2(KEYINPUT29), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT29), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n322), .B1(new_n298), .B2(new_n276), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n293), .B1(new_n267), .B2(new_n269), .ZN(new_n324));
  OAI221_X1 g138(.A(new_n317), .B1(new_n320), .B2(new_n321), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  AOI22_X1  g139(.A1(new_n316), .A2(KEYINPUT32), .B1(new_n325), .B2(G472), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n313), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G125), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n328), .A2(G140), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT16), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G140), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G125), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n328), .A2(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n331), .B1(new_n335), .B2(new_n330), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n188), .ZN(new_n337));
  OAI211_X1 g151(.A(new_n331), .B(G146), .C1(new_n335), .C2(new_n330), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n237), .A2(G128), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT73), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n238), .A2(new_n240), .A3(G128), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT67), .B(G119), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n344), .A2(KEYINPUT73), .A3(G128), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XNOR2_X1  g160(.A(KEYINPUT24), .B(G110), .ZN(new_n347));
  INV_X1    g161(.A(G110), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT23), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n344), .B2(G128), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n340), .A2(KEYINPUT23), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n350), .A2(new_n351), .A3(new_n342), .ZN(new_n352));
  OAI221_X1 g166(.A(new_n339), .B1(new_n346), .B2(new_n347), .C1(new_n348), .C2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n350), .A2(new_n348), .A3(new_n351), .A4(new_n342), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n343), .A2(new_n347), .A3(new_n345), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT74), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n333), .A2(new_n334), .A3(new_n188), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n338), .A2(new_n358), .ZN(new_n359));
  AND3_X1   g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n357), .B1(new_n356), .B2(new_n359), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n272), .A2(G221), .A3(G234), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(KEYINPUT75), .ZN(new_n364));
  XNOR2_X1  g178(.A(KEYINPUT22), .B(G137), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n364), .B(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n362), .A2(new_n367), .ZN(new_n368));
  OAI211_X1 g182(.A(new_n353), .B(new_n366), .C1(new_n360), .C2(new_n361), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT76), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT25), .ZN(new_n371));
  AOI21_X1  g185(.A(G902), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n370), .A2(new_n371), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g189(.A(KEYINPUT72), .B(G217), .Z(new_n376));
  AOI21_X1  g190(.A(new_n376), .B1(G234), .B2(new_n317), .ZN(new_n377));
  INV_X1    g191(.A(new_n374), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n368), .A2(new_n369), .A3(new_n378), .A4(new_n372), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n375), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n368), .A2(new_n369), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n377), .A2(G902), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(KEYINPUT77), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT9), .B(G234), .ZN(new_n387));
  OAI21_X1  g201(.A(G221), .B1(new_n387), .B2(G902), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n388), .B(KEYINPUT78), .ZN(new_n389));
  INV_X1    g203(.A(G104), .ZN(new_n390));
  OAI21_X1  g204(.A(KEYINPUT3), .B1(new_n390), .B2(G107), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT3), .ZN(new_n392));
  INV_X1    g206(.A(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n393), .A3(G104), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n390), .A2(G107), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT4), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n396), .A2(new_n397), .A3(G101), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(new_n197), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n396), .A2(G101), .ZN(new_n400));
  AOI21_X1  g214(.A(G101), .B1(new_n390), .B2(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n391), .A2(new_n401), .A3(new_n394), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n402), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT79), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n402), .A2(KEYINPUT4), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n400), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n399), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n210), .ZN(new_n409));
  NOR2_X1   g223(.A1(new_n390), .A2(G107), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n393), .A2(G104), .ZN(new_n411));
  OAI21_X1  g225(.A(G101), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n402), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(KEYINPUT80), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n402), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n262), .A2(new_n417), .A3(KEYINPUT10), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n222), .A2(new_n224), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(new_n257), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n420), .A2(new_n402), .A3(new_n412), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT10), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n408), .A2(new_n409), .A3(new_n418), .A4(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  INV_X1    g239(.A(G227), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n425), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n424), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT84), .ZN(new_n431));
  AOI21_X1  g245(.A(KEYINPUT12), .B1(new_n210), .B2(KEYINPUT81), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n413), .B1(new_n257), .B2(new_n419), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n412), .A2(new_n402), .A3(new_n415), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n415), .B1(new_n412), .B2(new_n402), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n433), .B1(new_n436), .B2(new_n229), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n432), .B1(new_n437), .B2(new_n409), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n421), .B1(new_n262), .B2(new_n417), .ZN(new_n439));
  INV_X1    g253(.A(new_n432), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n210), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT84), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n424), .A2(new_n443), .A3(new_n429), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n431), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n408), .A2(new_n418), .A3(new_n423), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n210), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n429), .B1(new_n447), .B2(new_n424), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  AOI211_X1 g263(.A(G469), .B(G902), .C1(new_n445), .C2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n429), .B1(new_n442), .B2(new_n424), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n424), .A2(KEYINPUT82), .A3(new_n429), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n452), .A2(new_n447), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT82), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n430), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n451), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G469), .B1(new_n456), .B2(G902), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n450), .B1(new_n457), .B2(KEYINPUT83), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n455), .A2(new_n447), .A3(new_n452), .ZN(new_n459));
  INV_X1    g273(.A(new_n451), .ZN(new_n460));
  AOI21_X1  g274(.A(G902), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G469), .ZN(new_n462));
  NOR3_X1   g276(.A1(new_n461), .A2(KEYINPUT83), .A3(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n389), .B1(new_n458), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g279(.A(G214), .B1(G237), .B2(G902), .ZN(new_n466));
  XNOR2_X1  g280(.A(G110), .B(G122), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n467), .B(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n398), .B1(new_n246), .B2(new_n248), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT85), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n470), .B(new_n471), .C1(new_n404), .C2(new_n407), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n241), .A2(KEYINPUT5), .A3(new_n243), .ZN(new_n473));
  OAI211_X1 g287(.A(new_n473), .B(G113), .C1(KEYINPUT5), .C2(new_n241), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n474), .B(new_n248), .C1(new_n434), .C2(new_n435), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n403), .A2(KEYINPUT79), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n406), .A2(new_n405), .A3(new_n400), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n471), .B1(new_n479), .B2(new_n470), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n469), .B1(new_n476), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n470), .B1(new_n404), .B2(new_n407), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(KEYINPUT85), .ZN(new_n483));
  XNOR2_X1  g297(.A(new_n467), .B(KEYINPUT86), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n475), .A4(new_n472), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(KEYINPUT6), .A3(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT87), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n197), .A2(new_n487), .A3(G125), .ZN(new_n488));
  INV_X1    g302(.A(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n487), .B1(new_n197), .B2(G125), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n229), .A2(new_n328), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n272), .A2(G224), .ZN(new_n494));
  XOR2_X1   g308(.A(new_n493), .B(new_n494), .Z(new_n495));
  INV_X1    g309(.A(KEYINPUT6), .ZN(new_n496));
  OAI211_X1 g310(.A(new_n496), .B(new_n469), .C1(new_n476), .C2(new_n480), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n486), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n494), .A2(KEYINPUT7), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n197), .A2(G125), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n499), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT8), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n484), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n469), .A2(KEYINPUT8), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n473), .ZN(new_n506));
  OAI21_X1  g320(.A(G113), .B1(new_n241), .B2(KEYINPUT5), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n248), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n413), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n505), .B1(new_n475), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n490), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n492), .A2(new_n511), .A3(new_n488), .A4(new_n499), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT88), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n491), .A2(new_n514), .A3(new_n492), .A4(new_n499), .ZN(new_n515));
  AOI211_X1 g329(.A(new_n501), .B(new_n510), .C1(new_n513), .C2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n516), .B2(new_n485), .ZN(new_n517));
  OAI21_X1  g331(.A(G210), .B1(G237), .B2(G902), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(KEYINPUT89), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n498), .A2(new_n517), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n520), .B1(new_n498), .B2(new_n517), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n466), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n271), .A2(new_n272), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n190), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n271), .A2(new_n272), .A3(G143), .A4(G214), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n208), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(G131), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n339), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n527), .A2(KEYINPUT17), .A3(G131), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n534), .A2(KEYINPUT96), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(KEYINPUT96), .ZN(new_n536));
  OAI211_X1 g350(.A(new_n532), .B(new_n533), .C1(new_n535), .C2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(G113), .B(G122), .ZN(new_n538));
  XNOR2_X1  g352(.A(KEYINPUT94), .B(G104), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n540), .B(KEYINPUT95), .Z(new_n541));
  INV_X1    g355(.A(KEYINPUT90), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n332), .A2(G125), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n542), .B1(new_n329), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n333), .A2(new_n334), .A3(KEYINPUT90), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(G146), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n358), .ZN(new_n547));
  AND4_X1   g361(.A1(KEYINPUT91), .A2(new_n528), .A3(KEYINPUT18), .A4(G131), .ZN(new_n548));
  AOI22_X1  g362(.A1(new_n528), .A2(KEYINPUT91), .B1(KEYINPUT18), .B2(G131), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n537), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n544), .A2(KEYINPUT19), .A3(new_n545), .ZN(new_n552));
  OR2_X1    g366(.A1(new_n335), .A2(KEYINPUT19), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n188), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT92), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n552), .A2(KEYINPUT92), .A3(new_n188), .A4(new_n553), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n556), .A2(KEYINPUT93), .A3(new_n338), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n529), .A2(new_n531), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND2_X1   g374(.A1(new_n557), .A2(new_n338), .ZN(new_n561));
  AOI21_X1  g375(.A(KEYINPUT93), .B1(new_n561), .B2(new_n556), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n550), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n551), .B1(new_n563), .B2(new_n540), .ZN(new_n564));
  NOR2_X1   g378(.A1(G475), .A2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(KEYINPUT20), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT20), .ZN(new_n568));
  INV_X1    g382(.A(new_n540), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT93), .ZN(new_n570));
  INV_X1    g384(.A(new_n556), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n557), .A2(new_n338), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n573), .A2(new_n559), .A3(new_n558), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n574), .B2(new_n550), .ZN(new_n575));
  OAI211_X1 g389(.A(new_n568), .B(new_n565), .C1(new_n575), .C2(new_n551), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n537), .A2(new_n550), .ZN(new_n577));
  NOR2_X1   g391(.A1(new_n577), .A2(new_n569), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n317), .B1(new_n578), .B2(new_n551), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n567), .A2(new_n576), .B1(G475), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(G478), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n581), .A2(KEYINPUT15), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n376), .A2(G953), .A3(new_n387), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n190), .A2(G128), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT13), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n219), .A2(G143), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n586), .A2(new_n587), .ZN(new_n591));
  OAI21_X1  g405(.A(G134), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n586), .A2(new_n589), .A3(new_n201), .ZN(new_n593));
  XNOR2_X1  g407(.A(G116), .B(G122), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(new_n393), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n393), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n592), .B(new_n593), .C1(new_n595), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n593), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n201), .B1(new_n586), .B2(new_n589), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT14), .ZN(new_n601));
  AND2_X1   g415(.A1(new_n594), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n242), .A2(KEYINPUT14), .A3(G122), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G107), .ZN(new_n604));
  OAI221_X1 g418(.A(new_n596), .B1(new_n599), .B2(new_n600), .C1(new_n602), .C2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT97), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n606), .B1(new_n598), .B2(new_n605), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n585), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n598), .A2(new_n605), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT97), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n584), .A3(new_n607), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n583), .B1(new_n614), .B2(new_n317), .ZN(new_n615));
  AOI211_X1 g429(.A(G902), .B(new_n582), .C1(new_n610), .C2(new_n613), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n272), .A2(G952), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(G234), .B2(G237), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(KEYINPUT21), .B(G898), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT98), .ZN(new_n622));
  NAND2_X1  g436(.A1(G234), .A2(G237), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(G902), .A3(G953), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n580), .A2(new_n617), .A3(new_n625), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n523), .A2(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n327), .A2(new_n386), .A3(new_n465), .A4(new_n627), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G101), .ZN(G3));
  INV_X1    g443(.A(new_n389), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n424), .A2(new_n443), .A3(new_n429), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n443), .B1(new_n424), .B2(new_n429), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n438), .A2(new_n441), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n462), .B(new_n317), .C1(new_n634), .C2(new_n448), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n452), .A2(new_n447), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT82), .B1(new_n424), .B2(new_n429), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n408), .A2(new_n418), .A3(new_n423), .ZN(new_n638));
  AOI22_X1  g452(.A1(new_n638), .A2(new_n409), .B1(new_n438), .B2(new_n441), .ZN(new_n639));
  OAI22_X1  g453(.A1(new_n636), .A2(new_n637), .B1(new_n639), .B2(new_n429), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n462), .B1(new_n640), .B2(new_n317), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT83), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n635), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n630), .B1(new_n643), .B2(new_n463), .ZN(new_n644));
  OAI21_X1  g458(.A(G472), .B1(new_n301), .B2(G902), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n304), .A2(new_n645), .A3(new_n312), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n644), .A2(new_n646), .A3(new_n385), .ZN(new_n647));
  OAI211_X1 g461(.A(new_n625), .B(new_n466), .C1(new_n521), .C2(new_n522), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n614), .B(KEYINPUT33), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n581), .A2(G902), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n608), .A2(new_n609), .A3(new_n585), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n584), .B1(new_n612), .B2(new_n607), .ZN(new_n652));
  OAI21_X1  g466(.A(new_n317), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n649), .A2(new_n650), .B1(new_n581), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n567), .A2(new_n576), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n579), .A2(G475), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n655), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n648), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n647), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT34), .B(G104), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G6));
  NAND2_X1  g477(.A1(new_n653), .A2(new_n582), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n614), .A2(new_n317), .A3(new_n583), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n580), .A2(new_n666), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n648), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n647), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  INV_X1    g485(.A(new_n646), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n362), .A2(KEYINPUT99), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT99), .ZN(new_n674));
  OAI211_X1 g488(.A(new_n353), .B(new_n674), .C1(new_n360), .C2(new_n361), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n367), .A2(KEYINPUT36), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n673), .A2(new_n677), .A3(new_n675), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n383), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n380), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n672), .A2(new_n465), .A3(new_n627), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  OAI211_X1 g499(.A(new_n466), .B(new_n682), .C1(new_n521), .C2(new_n522), .ZN(new_n686));
  INV_X1    g500(.A(G900), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(G953), .ZN(new_n688));
  AOI211_X1 g502(.A(new_n317), .B(new_n688), .C1(G234), .C2(G237), .ZN(new_n689));
  OR2_X1    g503(.A1(new_n689), .A2(KEYINPUT100), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(KEYINPUT100), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n620), .A3(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n580), .A2(new_n666), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n686), .A2(new_n693), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n327), .A2(new_n465), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT101), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT101), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n327), .A2(new_n697), .A3(new_n465), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G128), .ZN(G30));
  XNOR2_X1  g514(.A(new_n692), .B(KEYINPUT39), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n465), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT40), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n702), .B(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n617), .B1(new_n656), .B2(new_n657), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n709), .A2(new_n380), .A3(new_n466), .A4(new_n681), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT102), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n267), .A2(new_n269), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(new_n293), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n270), .A2(new_n293), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n319), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n316), .A2(KEYINPUT32), .B1(G472), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n313), .A2(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n498), .A2(new_n517), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n519), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n498), .A2(new_n517), .A3(new_n520), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XOR2_X1   g537(.A(new_n723), .B(KEYINPUT38), .Z(new_n724));
  NOR3_X1   g538(.A1(new_n711), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n705), .A2(new_n708), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G143), .ZN(G45));
  NAND3_X1  g541(.A1(new_n655), .A2(new_n658), .A3(new_n692), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n686), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n327), .A2(new_n465), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G146), .ZN(G48));
  NOR2_X1   g545(.A1(new_n462), .A2(KEYINPUT104), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n634), .A2(new_n448), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n732), .B1(new_n733), .B2(G902), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n445), .A2(new_n449), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n735), .B(new_n317), .C1(KEYINPUT104), .C2(new_n462), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n734), .A2(new_n736), .A3(new_n630), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n327), .A2(new_n386), .A3(new_n660), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND4_X1  g555(.A1(new_n327), .A2(new_n386), .A3(new_n668), .A4(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  NOR3_X1   g557(.A1(new_n737), .A2(new_n686), .A3(new_n626), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n327), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G119), .ZN(G21));
  INV_X1    g560(.A(new_n709), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n737), .A3(new_n648), .ZN(new_n748));
  AOI21_X1  g562(.A(new_n293), .B1(new_n320), .B2(KEYINPUT105), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n749), .B1(KEYINPUT105), .B2(new_n320), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n314), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n302), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n645), .A2(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(new_n385), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n748), .A2(new_n754), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G122), .ZN(G24));
  AND3_X1   g570(.A1(new_n645), .A2(new_n752), .A3(new_n682), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n737), .A2(new_n523), .ZN(new_n758));
  INV_X1    g572(.A(new_n728), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n757), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G125), .ZN(G27));
  OAI21_X1  g575(.A(new_n630), .B1(new_n450), .B2(new_n641), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n721), .A2(new_n466), .A3(new_n722), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n385), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n327), .A2(new_n764), .A3(new_n759), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT42), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n305), .B1(new_n301), .B2(new_n303), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n326), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n728), .A2(new_n766), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AOI22_X1  g584(.A1(new_n765), .A2(new_n766), .B1(new_n770), .B2(new_n764), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n208), .ZN(G33));
  INV_X1    g586(.A(new_n693), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n327), .A2(new_n764), .A3(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(new_n774), .B(G134), .ZN(G36));
  OR2_X1    g589(.A1(new_n456), .A2(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n456), .A2(KEYINPUT45), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(G469), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(KEYINPUT106), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n462), .A2(new_n317), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(KEYINPUT107), .A3(KEYINPUT46), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT106), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n778), .B(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(new_n780), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n784), .A2(KEYINPUT46), .A3(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT107), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n782), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n635), .B1(new_n781), .B2(KEYINPUT46), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n389), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n655), .A2(new_n580), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(KEYINPUT43), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n646), .A2(new_n682), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(KEYINPUT44), .ZN(new_n797));
  XOR2_X1   g611(.A(new_n763), .B(KEYINPUT108), .Z(new_n798));
  NAND4_X1  g612(.A1(new_n792), .A2(new_n701), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G137), .ZN(G39));
  NOR4_X1   g614(.A1(new_n327), .A2(new_n386), .A3(new_n728), .A4(new_n763), .ZN(new_n801));
  INV_X1    g615(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n792), .A2(KEYINPUT47), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT47), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n790), .B1(new_n788), .B2(new_n782), .ZN(new_n805));
  OAI21_X1  g619(.A(new_n804), .B1(new_n805), .B2(new_n389), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n802), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(new_n332), .ZN(G42));
  INV_X1    g622(.A(KEYINPUT53), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n723), .A2(new_n709), .A3(new_n466), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n635), .B1(new_n462), .B2(new_n461), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n380), .A2(new_n681), .A3(new_n692), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n630), .A3(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n810), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n814), .A2(new_n718), .ZN(new_n815));
  AND3_X1   g629(.A1(new_n730), .A2(new_n815), .A3(new_n760), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n699), .A2(KEYINPUT52), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT52), .B1(new_n699), .B2(new_n816), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n820), .B1(new_n615), .B2(new_n616), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n664), .A2(KEYINPUT110), .A3(new_n665), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n821), .A2(new_n822), .A3(new_n692), .ZN(new_n823));
  AOI21_X1  g637(.A(KEYINPUT112), .B1(new_n823), .B2(new_n580), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n721), .A2(new_n682), .A3(new_n466), .A4(new_n722), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n823), .A2(new_n580), .A3(KEYINPUT112), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n327), .A2(new_n826), .A3(new_n465), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n762), .A2(new_n763), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n757), .A2(new_n759), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n774), .A3(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n771), .A2(new_n831), .ZN(new_n832));
  AND4_X1   g646(.A1(new_n304), .A2(new_n645), .A3(new_n312), .A4(new_n386), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT109), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n648), .B2(new_n659), .ZN(new_n835));
  INV_X1    g649(.A(new_n466), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n836), .B1(new_n721), .B2(new_n722), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n580), .A2(new_n654), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n838), .A3(KEYINPUT109), .A4(new_n625), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n833), .A2(new_n835), .A3(new_n465), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(new_n628), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT111), .ZN(new_n842));
  INV_X1    g656(.A(new_n821), .ZN(new_n843));
  INV_X1    g657(.A(new_n822), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n580), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n648), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n833), .A2(new_n846), .A3(new_n465), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n683), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n841), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n683), .A2(new_n847), .A3(KEYINPUT111), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n739), .A2(new_n742), .A3(new_n755), .A4(new_n745), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n832), .A2(new_n849), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n809), .B1(new_n819), .B2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n831), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n765), .A2(new_n766), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n770), .A2(new_n764), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n848), .A2(new_n842), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n859), .A2(new_n628), .A3(new_n850), .A4(new_n840), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n644), .B1(new_n313), .B2(new_n326), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n697), .B1(new_n863), .B2(new_n694), .ZN(new_n864));
  AND4_X1   g678(.A1(new_n697), .A2(new_n327), .A3(new_n465), .A4(new_n694), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n730), .A2(new_n815), .A3(new_n760), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n862), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n699), .A2(new_n816), .A3(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n861), .A2(new_n870), .A3(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n853), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g686(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n873));
  NOR2_X1   g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n874), .B1(KEYINPUT54), .B2(new_n872), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT116), .ZN(new_n876));
  OR3_X1    g690(.A1(new_n737), .A2(new_n763), .A3(new_n876), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n876), .B1(new_n737), .B2(new_n763), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n877), .A2(new_n619), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(new_n794), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n768), .A2(new_n386), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g696(.A(KEYINPUT118), .B(KEYINPUT48), .ZN(new_n883));
  XNOR2_X1  g697(.A(new_n882), .B(new_n883), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n794), .A2(new_n385), .A3(new_n620), .A4(new_n753), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n618), .B1(new_n885), .B2(new_n758), .ZN(new_n886));
  OR3_X1    g700(.A1(new_n879), .A2(new_n385), .A3(new_n718), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n884), .B(new_n886), .C1(new_n659), .C2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n734), .A2(new_n736), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(new_n389), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n803), .A2(new_n806), .A3(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n885), .A2(new_n798), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR3_X1   g707(.A1(new_n887), .A2(new_n658), .A3(new_n655), .ZN(new_n894));
  INV_X1    g708(.A(new_n757), .ZN(new_n895));
  OR3_X1    g709(.A1(new_n880), .A2(KEYINPUT117), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(KEYINPUT117), .B1(new_n880), .B2(new_n895), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n894), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n738), .A2(new_n836), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(KEYINPUT114), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n900), .A2(new_n724), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(KEYINPUT115), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT115), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n900), .A2(new_n904), .A3(new_n724), .A4(new_n901), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n885), .A3(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT50), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(KEYINPUT50), .A3(new_n885), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n893), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT51), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n888), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n893), .A2(new_n911), .A3(KEYINPUT51), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n875), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n916), .B1(G952), .B2(G953), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n889), .B(KEYINPUT49), .ZN(new_n918));
  NOR4_X1   g732(.A1(new_n793), .A2(new_n385), .A3(new_n389), .A4(new_n836), .ZN(new_n919));
  NAND4_X1  g733(.A1(new_n918), .A2(new_n719), .A3(new_n724), .A4(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n917), .A2(new_n920), .ZN(G75));
  NAND2_X1  g735(.A1(new_n486), .A2(new_n497), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n495), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT55), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(KEYINPUT56), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n928), .B1(new_n872), .B2(G902), .ZN(new_n929));
  AOI211_X1 g743(.A(KEYINPUT119), .B(new_n317), .C1(new_n853), .C2(new_n871), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  AOI21_X1  g745(.A(new_n927), .B1(new_n931), .B2(new_n519), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n272), .A2(G952), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n317), .B1(new_n853), .B2(new_n871), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT56), .B1(new_n935), .B2(new_n519), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n936), .B2(new_n925), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT120), .B1(new_n932), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n935), .A2(new_n519), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n926), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n933), .B1(new_n940), .B2(new_n924), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n929), .A2(new_n930), .A3(new_n520), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n941), .B(new_n942), .C1(new_n943), .C2(new_n927), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n938), .A2(new_n944), .ZN(G51));
  XNOR2_X1  g759(.A(new_n780), .B(KEYINPUT57), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n872), .A2(new_n873), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(new_n874), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n735), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n931), .A2(new_n779), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n933), .B1(new_n950), .B2(new_n951), .ZN(G54));
  AND2_X1   g766(.A1(KEYINPUT58), .A2(G475), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n931), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n954), .A2(new_n564), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n931), .B(new_n953), .C1(new_n551), .C2(new_n575), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n955), .A2(new_n934), .A3(new_n956), .ZN(G60));
  INV_X1    g771(.A(KEYINPUT121), .ZN(new_n958));
  INV_X1    g772(.A(new_n649), .ZN(new_n959));
  NAND2_X1  g773(.A1(G478), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT59), .Z(new_n961));
  NOR2_X1   g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n962), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n872), .A2(new_n873), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n947), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n958), .B1(new_n965), .B2(new_n933), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n962), .B1(new_n948), .B2(new_n874), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n967), .A2(KEYINPUT121), .A3(new_n934), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n959), .B1(new_n875), .B2(new_n961), .ZN(new_n969));
  AND3_X1   g783(.A1(new_n966), .A2(new_n968), .A3(new_n969), .ZN(G63));
  INV_X1    g784(.A(new_n872), .ZN(new_n971));
  XNOR2_X1  g785(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n972));
  NAND2_X1  g786(.A1(G217), .A2(G902), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n975), .A2(new_n680), .A3(new_n679), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n381), .B(KEYINPUT123), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n977), .B1(new_n971), .B2(new_n974), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n976), .A2(new_n934), .A3(new_n978), .ZN(new_n979));
  INV_X1    g793(.A(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n976), .A2(KEYINPUT61), .A3(new_n934), .A4(new_n978), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(G66));
  AOI21_X1  g797(.A(new_n272), .B1(new_n622), .B2(G224), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT124), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n986));
  INV_X1    g800(.A(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n985), .B1(new_n987), .B2(G953), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT125), .Z(new_n989));
  OAI21_X1  g803(.A(new_n922), .B1(G898), .B2(new_n272), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G69));
  OAI21_X1  g805(.A(G953), .B1(new_n426), .B2(new_n687), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n236), .A2(new_n256), .A3(new_n266), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n552), .A2(new_n553), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  XNOR2_X1  g810(.A(new_n996), .B(KEYINPUT126), .ZN(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  AND3_X1   g812(.A1(new_n699), .A2(new_n730), .A3(new_n760), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n726), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  XNOR2_X1  g815(.A(new_n1000), .B(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n803), .A2(new_n806), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(new_n801), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n763), .B1(new_n659), .B2(new_n845), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n703), .A2(new_n327), .A3(new_n386), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n799), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1002), .A2(new_n1004), .A3(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n998), .B1(new_n1008), .B2(new_n272), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n881), .A2(new_n810), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n792), .A2(new_n701), .A3(new_n1011), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n857), .A2(new_n774), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n799), .A2(new_n1012), .A3(new_n999), .A4(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n272), .B1(new_n1014), .B2(new_n807), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n996), .B1(new_n1015), .B2(new_n688), .ZN(new_n1016));
  INV_X1    g830(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n993), .B1(new_n1010), .B2(new_n1017), .ZN(new_n1018));
  NOR3_X1   g832(.A1(new_n1009), .A2(new_n1016), .A3(new_n992), .ZN(new_n1019));
  NOR2_X1   g833(.A1(new_n1018), .A2(new_n1019), .ZN(G72));
  NAND4_X1  g834(.A1(new_n1002), .A2(new_n1007), .A3(new_n1004), .A4(new_n987), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  AOI21_X1  g837(.A(new_n713), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n1024), .A2(KEYINPUT127), .ZN(new_n1025));
  NOR3_X1   g839(.A1(new_n1014), .A2(new_n807), .A3(new_n986), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1023), .ZN(new_n1027));
  OAI211_X1 g841(.A(new_n267), .B(new_n714), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n324), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1027), .B1(new_n1029), .B2(new_n278), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n933), .B1(new_n872), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1028), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT127), .ZN(new_n1033));
  AOI211_X1 g847(.A(new_n1033), .B(new_n713), .C1(new_n1021), .C2(new_n1023), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1025), .A2(new_n1032), .A3(new_n1034), .ZN(G57));
endmodule


