

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734;

  OR2_X1 U364 ( .A1(n375), .A2(n598), .ZN(n374) );
  OR2_X1 U365 ( .A1(n610), .A2(n649), .ZN(n596) );
  XNOR2_X1 U366 ( .A(n419), .B(KEYINPUT87), .ZN(n415) );
  XNOR2_X1 U367 ( .A(n522), .B(n521), .ZN(n647) );
  XNOR2_X2 U368 ( .A(KEYINPUT64), .B(KEYINPUT79), .ZN(n440) );
  INV_X1 U369 ( .A(n629), .ZN(n342) );
  BUF_X1 U370 ( .A(n690), .Z(n702) );
  AND2_X1 U371 ( .A1(n693), .A2(G475), .ZN(n695) );
  AND2_X1 U372 ( .A1(n382), .A2(n379), .ZN(n378) );
  NAND2_X1 U373 ( .A1(n377), .A2(n349), .ZN(n376) );
  XNOR2_X1 U374 ( .A(n427), .B(KEYINPUT41), .ZN(n677) );
  XNOR2_X1 U375 ( .A(n590), .B(n577), .ZN(n598) );
  XNOR2_X1 U376 ( .A(n415), .B(KEYINPUT19), .ZN(n574) );
  XNOR2_X1 U377 ( .A(n389), .B(G469), .ZN(n538) );
  OR2_X1 U378 ( .A1(n687), .A2(G902), .ZN(n389) );
  XNOR2_X1 U379 ( .A(n464), .B(n463), .ZN(n706) );
  XNOR2_X1 U380 ( .A(n495), .B(n442), .ZN(n454) );
  XNOR2_X1 U381 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U382 ( .A(n461), .B(n460), .ZN(n471) );
  BUF_X1 U383 ( .A(n732), .Z(n343) );
  INV_X1 U384 ( .A(n601), .ZN(n344) );
  NOR2_X2 U385 ( .A1(n714), .A2(n726), .ZN(n615) );
  XNOR2_X2 U386 ( .A(n368), .B(n435), .ZN(n714) );
  XNOR2_X1 U387 ( .A(n538), .B(n388), .ZN(n610) );
  BUF_X1 U388 ( .A(n714), .Z(n345) );
  XNOR2_X1 U389 ( .A(n390), .B(n351), .ZN(n346) );
  BUF_X1 U390 ( .A(n590), .Z(n347) );
  XNOR2_X1 U391 ( .A(n390), .B(n351), .ZN(n391) );
  INV_X1 U392 ( .A(n505), .ZN(n424) );
  NAND2_X1 U393 ( .A1(n561), .A2(n562), .ZN(n667) );
  XNOR2_X1 U394 ( .A(G101), .B(G110), .ZN(n460) );
  XOR2_X1 U395 ( .A(G104), .B(G107), .Z(n461) );
  XNOR2_X1 U396 ( .A(KEYINPUT10), .B(n477), .ZN(n721) );
  INV_X1 U397 ( .A(KEYINPUT4), .ZN(n442) );
  NOR2_X1 U398 ( .A1(n413), .A2(n411), .ZN(n423) );
  XNOR2_X1 U399 ( .A(n414), .B(n358), .ZN(n413) );
  NOR2_X1 U400 ( .A1(G953), .A2(G237), .ZN(n484) );
  NAND2_X1 U401 ( .A1(n409), .A2(n406), .ZN(n655) );
  OR2_X1 U402 ( .A1(n503), .A2(n407), .ZN(n406) );
  AND2_X1 U403 ( .A1(n405), .A2(n410), .ZN(n409) );
  NAND2_X1 U404 ( .A1(n504), .A2(n408), .ZN(n407) );
  XNOR2_X1 U405 ( .A(G116), .B(G113), .ZN(n444) );
  XNOR2_X1 U406 ( .A(n493), .B(n492), .ZN(n432) );
  XNOR2_X1 U407 ( .A(n494), .B(n431), .ZN(n430) );
  XNOR2_X1 U408 ( .A(G134), .B(G116), .ZN(n494) );
  XNOR2_X1 U409 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n431) );
  XOR2_X1 U410 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n499) );
  XNOR2_X1 U411 ( .A(G131), .B(G143), .ZN(n481) );
  XOR2_X1 U412 ( .A(G122), .B(G140), .Z(n475) );
  XNOR2_X1 U413 ( .A(n720), .B(n472), .ZN(n687) );
  NAND2_X1 U414 ( .A1(n429), .A2(n428), .ZN(n427) );
  INV_X1 U415 ( .A(n667), .ZN(n428) );
  INV_X1 U416 ( .A(n661), .ZN(n429) );
  XNOR2_X1 U417 ( .A(n426), .B(n551), .ZN(n566) );
  NOR2_X1 U418 ( .A1(n564), .A2(n550), .ZN(n426) );
  XNOR2_X1 U419 ( .A(n402), .B(n401), .ZN(n552) );
  INV_X1 U420 ( .A(KEYINPUT108), .ZN(n401) );
  NAND2_X1 U421 ( .A1(n403), .A2(n342), .ZN(n402) );
  XNOR2_X1 U422 ( .A(n502), .B(n350), .ZN(n562) );
  NOR2_X1 U423 ( .A1(n548), .A2(n649), .ZN(n579) );
  INV_X1 U424 ( .A(KEYINPUT1), .ZN(n388) );
  XNOR2_X1 U425 ( .A(n517), .B(n516), .ZN(n704) );
  XNOR2_X1 U426 ( .A(n721), .B(n506), .ZN(n517) );
  XNOR2_X1 U427 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U428 ( .A(n505), .B(KEYINPUT23), .ZN(n506) );
  XNOR2_X1 U429 ( .A(n685), .B(n684), .ZN(n686) );
  INV_X1 U430 ( .A(G953), .ZN(n728) );
  XNOR2_X1 U431 ( .A(n644), .B(n643), .ZN(n645) );
  INV_X1 U432 ( .A(G902), .ZN(n408) );
  NAND2_X1 U433 ( .A1(G472), .A2(G902), .ZN(n410) );
  XOR2_X1 U434 ( .A(G146), .B(G125), .Z(n476) );
  XNOR2_X1 U435 ( .A(KEYINPUT100), .B(KEYINPUT12), .ZN(n478) );
  XOR2_X1 U436 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n479) );
  XOR2_X1 U437 ( .A(G902), .B(KEYINPUT15), .Z(n611) );
  INV_X1 U438 ( .A(KEYINPUT18), .ZN(n455) );
  XNOR2_X1 U439 ( .A(n533), .B(n404), .ZN(n403) );
  INV_X1 U440 ( .A(KEYINPUT107), .ZN(n404) );
  AND2_X1 U441 ( .A1(n386), .A2(n600), .ZN(n385) );
  OR2_X1 U442 ( .A1(n679), .A2(n355), .ZN(n375) );
  XNOR2_X1 U443 ( .A(G131), .B(G134), .ZN(n443) );
  XNOR2_X1 U444 ( .A(G101), .B(KEYINPUT75), .ZN(n449) );
  XOR2_X1 U445 ( .A(KEYINPUT5), .B(G137), .Z(n447) );
  INV_X1 U446 ( .A(KEYINPUT45), .ZN(n435) );
  XOR2_X1 U447 ( .A(G137), .B(G140), .Z(n505) );
  NOR2_X1 U448 ( .A1(n383), .A2(n381), .ZN(n380) );
  XNOR2_X1 U449 ( .A(n655), .B(KEYINPUT6), .ZN(n603) );
  NAND2_X1 U450 ( .A1(n655), .A2(n664), .ZN(n545) );
  XNOR2_X1 U451 ( .A(KEYINPUT66), .B(KEYINPUT22), .ZN(n591) );
  XNOR2_X1 U452 ( .A(n471), .B(n462), .ZN(n463) );
  XOR2_X1 U453 ( .A(G122), .B(KEYINPUT16), .Z(n462) );
  XNOR2_X1 U454 ( .A(n432), .B(n430), .ZN(n497) );
  XNOR2_X1 U455 ( .A(G113), .B(G104), .ZN(n474) );
  XNOR2_X1 U456 ( .A(n544), .B(KEYINPUT42), .ZN(n733) );
  XNOR2_X1 U457 ( .A(n425), .B(KEYINPUT40), .ZN(n734) );
  NAND2_X1 U458 ( .A1(n566), .A2(n342), .ZN(n425) );
  NAND2_X1 U459 ( .A1(n555), .A2(n601), .ZN(n637) );
  AND2_X1 U460 ( .A1(n579), .A2(n606), .ZN(n366) );
  XNOR2_X1 U461 ( .A(n703), .B(n704), .ZN(n395) );
  XNOR2_X1 U462 ( .A(n691), .B(n692), .ZN(n394) );
  INV_X1 U463 ( .A(KEYINPUT56), .ZN(n420) );
  INV_X1 U464 ( .A(KEYINPUT53), .ZN(n397) );
  NAND2_X1 U465 ( .A1(n400), .A2(n399), .ZN(n398) );
  AND2_X1 U466 ( .A1(n682), .A2(n728), .ZN(n399) );
  AND2_X1 U467 ( .A1(n578), .A2(n366), .ZN(n348) );
  AND2_X1 U468 ( .A1(n383), .A2(n381), .ZN(n349) );
  XOR2_X1 U469 ( .A(n491), .B(KEYINPUT105), .Z(n350) );
  AND2_X1 U470 ( .A1(n473), .A2(G210), .ZN(n351) );
  XOR2_X1 U471 ( .A(KEYINPUT3), .B(G119), .Z(n352) );
  XOR2_X1 U472 ( .A(KEYINPUT81), .B(n627), .Z(n353) );
  NOR2_X1 U473 ( .A1(n537), .A2(n346), .ZN(n354) );
  XNOR2_X1 U474 ( .A(KEYINPUT78), .B(n599), .ZN(n355) );
  XNOR2_X1 U475 ( .A(n387), .B(n424), .ZN(n720) );
  XOR2_X1 U476 ( .A(n697), .B(n696), .Z(n356) );
  XOR2_X1 U477 ( .A(n503), .B(KEYINPUT62), .Z(n357) );
  XOR2_X1 U478 ( .A(KEYINPUT46), .B(KEYINPUT85), .Z(n358) );
  NOR2_X1 U479 ( .A1(G952), .A2(n728), .ZN(n705) );
  INV_X1 U480 ( .A(n705), .ZN(n392) );
  NOR2_X1 U481 ( .A1(n714), .A2(n726), .ZN(n359) );
  AND2_X1 U482 ( .A1(n393), .A2(n392), .ZN(n699) );
  XNOR2_X1 U483 ( .A(n698), .B(n356), .ZN(n393) );
  NAND2_X1 U484 ( .A1(n614), .A2(n613), .ZN(n360) );
  NAND2_X1 U485 ( .A1(n614), .A2(n613), .ZN(n694) );
  XNOR2_X1 U486 ( .A(n398), .B(n397), .ZN(G75) );
  XNOR2_X1 U487 ( .A(n423), .B(n438), .ZN(n565) );
  NAND2_X1 U488 ( .A1(n645), .A2(n693), .ZN(n400) );
  NOR2_X1 U489 ( .A1(n353), .A2(n560), .ZN(n412) );
  NAND2_X1 U490 ( .A1(n454), .A2(n437), .ZN(n363) );
  NAND2_X1 U491 ( .A1(n361), .A2(n362), .ZN(n364) );
  NAND2_X1 U492 ( .A1(n363), .A2(n364), .ZN(n436) );
  INV_X1 U493 ( .A(n454), .ZN(n361) );
  INV_X1 U494 ( .A(n437), .ZN(n362) );
  XNOR2_X1 U495 ( .A(n458), .B(KEYINPUT77), .ZN(n437) );
  XNOR2_X1 U496 ( .A(n436), .B(n457), .ZN(n466) );
  XNOR2_X1 U497 ( .A(n466), .B(n465), .ZN(n683) );
  AND2_X1 U498 ( .A1(n373), .A2(n616), .ZN(n369) );
  XNOR2_X1 U499 ( .A(n700), .B(n701), .ZN(n396) );
  XNOR2_X1 U500 ( .A(n418), .B(n357), .ZN(n417) );
  XNOR2_X1 U501 ( .A(n422), .B(n686), .ZN(n365) );
  NAND2_X1 U502 ( .A1(n365), .A2(n392), .ZN(n421) );
  NAND2_X1 U503 ( .A1(n417), .A2(n392), .ZN(n416) );
  NAND2_X1 U504 ( .A1(n623), .A2(n367), .ZN(n372) );
  XNOR2_X1 U505 ( .A(n367), .B(G119), .ZN(G21) );
  XNOR2_X2 U506 ( .A(n433), .B(n605), .ZN(n367) );
  NAND2_X1 U507 ( .A1(n370), .A2(n369), .ZN(n368) );
  XNOR2_X1 U508 ( .A(n371), .B(KEYINPUT44), .ZN(n370) );
  NOR2_X2 U509 ( .A1(n732), .A2(n372), .ZN(n371) );
  NAND2_X1 U510 ( .A1(n378), .A2(n376), .ZN(n732) );
  NAND2_X1 U511 ( .A1(n587), .A2(n586), .ZN(n373) );
  NAND2_X1 U512 ( .A1(n385), .A2(n374), .ZN(n384) );
  XNOR2_X2 U513 ( .A(n576), .B(n575), .ZN(n590) );
  XNOR2_X1 U514 ( .A(n597), .B(KEYINPUT33), .ZN(n679) );
  INV_X1 U515 ( .A(n384), .ZN(n377) );
  INV_X1 U516 ( .A(n380), .ZN(n379) );
  INV_X1 U517 ( .A(KEYINPUT35), .ZN(n381) );
  NAND2_X1 U518 ( .A1(n384), .A2(KEYINPUT35), .ZN(n382) );
  NAND2_X1 U519 ( .A1(n598), .A2(n355), .ZN(n383) );
  NAND2_X1 U520 ( .A1(n679), .A2(n355), .ZN(n386) );
  XNOR2_X1 U521 ( .A(n387), .B(n453), .ZN(n503) );
  XNOR2_X1 U522 ( .A(n454), .B(n443), .ZN(n387) );
  NAND2_X1 U523 ( .A1(n391), .A2(n664), .ZN(n419) );
  NAND2_X1 U524 ( .A1(n683), .A2(n518), .ZN(n390) );
  XNOR2_X1 U525 ( .A(n346), .B(KEYINPUT38), .ZN(n550) );
  NAND2_X1 U526 ( .A1(n600), .A2(n346), .ZN(n563) );
  NOR2_X1 U527 ( .A1(n394), .A2(n705), .ZN(G54) );
  NOR2_X1 U528 ( .A1(n395), .A2(n705), .ZN(G66) );
  NAND2_X1 U529 ( .A1(n615), .A2(n611), .ZN(n614) );
  NOR2_X1 U530 ( .A1(n396), .A2(n705), .ZN(G63) );
  NAND2_X1 U531 ( .A1(n552), .A2(n415), .ZN(n553) );
  NAND2_X1 U532 ( .A1(n503), .A2(G472), .ZN(n405) );
  NAND2_X1 U533 ( .A1(n733), .A2(n734), .ZN(n414) );
  NAND2_X1 U534 ( .A1(n412), .A2(n637), .ZN(n411) );
  XNOR2_X1 U535 ( .A(n416), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U536 ( .A1(n690), .A2(G472), .ZN(n418) );
  XNOR2_X1 U537 ( .A(n421), .B(n420), .ZN(G51) );
  NAND2_X1 U538 ( .A1(n690), .A2(G210), .ZN(n422) );
  NOR2_X2 U539 ( .A1(n574), .A2(n573), .ZN(n576) );
  NAND2_X1 U540 ( .A1(n607), .A2(n604), .ZN(n433) );
  XNOR2_X2 U541 ( .A(n434), .B(n591), .ZN(n607) );
  NOR2_X2 U542 ( .A1(n590), .A2(n589), .ZN(n434) );
  XOR2_X1 U543 ( .A(KEYINPUT48), .B(KEYINPUT84), .Z(n438) );
  INV_X1 U544 ( .A(G146), .ZN(n448) );
  XNOR2_X1 U545 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U546 ( .A(G128), .B(G143), .ZN(n439) );
  XNOR2_X1 U547 ( .A(n451), .B(n450), .ZN(n452) );
  INV_X1 U548 ( .A(KEYINPUT91), .ZN(n577) );
  XNOR2_X1 U549 ( .A(n459), .B(n452), .ZN(n453) );
  XNOR2_X1 U550 ( .A(n471), .B(n470), .ZN(n472) );
  INV_X1 U551 ( .A(KEYINPUT80), .ZN(n643) );
  XNOR2_X1 U552 ( .A(n520), .B(KEYINPUT25), .ZN(n521) );
  INV_X1 U553 ( .A(G472), .ZN(n504) );
  INV_X1 U554 ( .A(KEYINPUT39), .ZN(n551) );
  INV_X1 U555 ( .A(n439), .ZN(n441) );
  XNOR2_X2 U556 ( .A(n441), .B(n440), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n352), .B(n444), .ZN(n445) );
  XNOR2_X1 U558 ( .A(KEYINPUT71), .B(n445), .ZN(n459) );
  NAND2_X1 U559 ( .A1(n484), .A2(G210), .ZN(n446) );
  XNOR2_X1 U560 ( .A(n447), .B(n446), .ZN(n451) );
  XOR2_X1 U561 ( .A(n476), .B(KEYINPUT17), .Z(n456) );
  NAND2_X1 U562 ( .A1(G224), .A2(n728), .ZN(n458) );
  INV_X1 U563 ( .A(n459), .ZN(n464) );
  INV_X1 U564 ( .A(n706), .ZN(n465) );
  INV_X1 U565 ( .A(n611), .ZN(n518) );
  NOR2_X1 U566 ( .A1(G237), .A2(G902), .ZN(n467) );
  XOR2_X1 U567 ( .A(KEYINPUT74), .B(n467), .Z(n473) );
  XOR2_X1 U568 ( .A(G146), .B(KEYINPUT76), .Z(n469) );
  NAND2_X1 U569 ( .A1(G227), .A2(n728), .ZN(n468) );
  XNOR2_X1 U570 ( .A(n469), .B(n468), .ZN(n470) );
  INV_X1 U571 ( .A(n610), .ZN(n601) );
  NAND2_X1 U572 ( .A1(G214), .A2(n473), .ZN(n664) );
  XNOR2_X1 U573 ( .A(n475), .B(n474), .ZN(n488) );
  INV_X1 U574 ( .A(n476), .ZN(n477) );
  XNOR2_X1 U575 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U576 ( .A(n480), .B(KEYINPUT11), .Z(n482) );
  XNOR2_X1 U577 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U578 ( .A(n721), .B(n483), .Z(n486) );
  NAND2_X1 U579 ( .A1(G214), .A2(n484), .ZN(n485) );
  XNOR2_X1 U580 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U581 ( .A(n488), .B(n487), .ZN(n697) );
  NOR2_X1 U582 ( .A1(G902), .A2(n697), .ZN(n490) );
  XNOR2_X1 U583 ( .A(KEYINPUT13), .B(G475), .ZN(n489) );
  XNOR2_X1 U584 ( .A(n490), .B(n489), .ZN(n558) );
  XNOR2_X1 U585 ( .A(G478), .B(KEYINPUT104), .ZN(n491) );
  XOR2_X1 U586 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n493) );
  XNOR2_X1 U587 ( .A(G107), .B(G122), .ZN(n492) );
  XNOR2_X1 U588 ( .A(n495), .B(KEYINPUT103), .ZN(n496) );
  XNOR2_X1 U589 ( .A(n497), .B(n496), .ZN(n501) );
  NAND2_X1 U590 ( .A1(G234), .A2(n728), .ZN(n498) );
  XNOR2_X1 U591 ( .A(n499), .B(n498), .ZN(n513) );
  NAND2_X1 U592 ( .A1(G217), .A2(n513), .ZN(n500) );
  XOR2_X1 U593 ( .A(n501), .B(n500), .Z(n701) );
  NOR2_X1 U594 ( .A1(G902), .A2(n701), .ZN(n502) );
  NAND2_X1 U595 ( .A1(n558), .A2(n562), .ZN(n629) );
  XOR2_X1 U596 ( .A(KEYINPUT93), .B(G110), .Z(n508) );
  XNOR2_X1 U597 ( .A(G128), .B(G119), .ZN(n507) );
  XNOR2_X1 U598 ( .A(n508), .B(n507), .ZN(n512) );
  XOR2_X1 U599 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n510) );
  XNOR2_X1 U600 ( .A(KEYINPUT82), .B(KEYINPUT72), .ZN(n509) );
  XNOR2_X1 U601 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U602 ( .A(n512), .B(n511), .ZN(n515) );
  NAND2_X1 U603 ( .A1(G221), .A2(n513), .ZN(n514) );
  NOR2_X1 U604 ( .A1(G902), .A2(n704), .ZN(n522) );
  NAND2_X1 U605 ( .A1(n518), .A2(G234), .ZN(n519) );
  XNOR2_X1 U606 ( .A(n519), .B(KEYINPUT20), .ZN(n528) );
  NAND2_X1 U607 ( .A1(n528), .A2(G217), .ZN(n520) );
  NAND2_X1 U608 ( .A1(G234), .A2(G237), .ZN(n523) );
  XNOR2_X1 U609 ( .A(n523), .B(KEYINPUT14), .ZN(n524) );
  NAND2_X1 U610 ( .A1(G952), .A2(n524), .ZN(n676) );
  NOR2_X1 U611 ( .A1(G953), .A2(n676), .ZN(n572) );
  AND2_X1 U612 ( .A1(G953), .A2(n524), .ZN(n525) );
  NAND2_X1 U613 ( .A1(G902), .A2(n525), .ZN(n568) );
  NOR2_X1 U614 ( .A1(G900), .A2(n568), .ZN(n526) );
  XNOR2_X1 U615 ( .A(n526), .B(KEYINPUT106), .ZN(n527) );
  NOR2_X1 U616 ( .A1(n572), .A2(n527), .ZN(n547) );
  NAND2_X1 U617 ( .A1(G221), .A2(n528), .ZN(n529) );
  XNOR2_X1 U618 ( .A(KEYINPUT21), .B(n529), .ZN(n588) );
  NOR2_X1 U619 ( .A1(n547), .A2(n588), .ZN(n530) );
  XOR2_X1 U620 ( .A(KEYINPUT70), .B(n530), .Z(n531) );
  NOR2_X1 U621 ( .A1(n647), .A2(n531), .ZN(n532) );
  XNOR2_X1 U622 ( .A(n532), .B(KEYINPUT69), .ZN(n539) );
  NOR2_X1 U623 ( .A1(n603), .A2(n539), .ZN(n533) );
  NAND2_X1 U624 ( .A1(n664), .A2(n552), .ZN(n534) );
  XOR2_X1 U625 ( .A(KEYINPUT109), .B(n534), .Z(n535) );
  NOR2_X1 U626 ( .A1(n601), .A2(n535), .ZN(n536) );
  XNOR2_X1 U627 ( .A(n536), .B(KEYINPUT43), .ZN(n537) );
  INV_X1 U628 ( .A(n538), .ZN(n548) );
  XNOR2_X1 U629 ( .A(n548), .B(KEYINPUT110), .ZN(n543) );
  XNOR2_X1 U630 ( .A(KEYINPUT111), .B(KEYINPUT28), .ZN(n541) );
  INV_X1 U631 ( .A(n655), .ZN(n606) );
  NOR2_X1 U632 ( .A1(n606), .A2(n539), .ZN(n540) );
  XNOR2_X1 U633 ( .A(n541), .B(n540), .ZN(n542) );
  NOR2_X1 U634 ( .A1(n543), .A2(n542), .ZN(n557) );
  INV_X1 U635 ( .A(n550), .ZN(n665) );
  NAND2_X1 U636 ( .A1(n665), .A2(n664), .ZN(n661) );
  INV_X1 U637 ( .A(n558), .ZN(n561) );
  NAND2_X1 U638 ( .A1(n557), .A2(n677), .ZN(n544) );
  XNOR2_X1 U639 ( .A(KEYINPUT30), .B(n545), .ZN(n546) );
  NOR2_X1 U640 ( .A1(n547), .A2(n546), .ZN(n549) );
  INV_X1 U641 ( .A(n588), .ZN(n646) );
  NAND2_X1 U642 ( .A1(n647), .A2(n646), .ZN(n649) );
  NAND2_X1 U643 ( .A1(n549), .A2(n579), .ZN(n564) );
  XOR2_X1 U644 ( .A(KEYINPUT112), .B(KEYINPUT36), .Z(n554) );
  XNOR2_X1 U645 ( .A(n554), .B(n553), .ZN(n555) );
  INV_X1 U646 ( .A(n574), .ZN(n556) );
  NAND2_X1 U647 ( .A1(n557), .A2(n556), .ZN(n628) );
  NOR2_X1 U648 ( .A1(n558), .A2(n562), .ZN(n633) );
  NOR2_X1 U649 ( .A1(n342), .A2(n633), .ZN(n662) );
  NOR2_X1 U650 ( .A1(n628), .A2(n662), .ZN(n559) );
  XOR2_X1 U651 ( .A(KEYINPUT47), .B(n559), .Z(n560) );
  NOR2_X1 U652 ( .A1(n562), .A2(n561), .ZN(n600) );
  NOR2_X1 U653 ( .A1(n564), .A2(n563), .ZN(n627) );
  NOR2_X1 U654 ( .A1(n354), .A2(n565), .ZN(n567) );
  NAND2_X1 U655 ( .A1(n633), .A2(n566), .ZN(n638) );
  NAND2_X1 U656 ( .A1(n567), .A2(n638), .ZN(n726) );
  INV_X1 U657 ( .A(n568), .ZN(n569) );
  XNOR2_X1 U658 ( .A(KEYINPUT89), .B(G898), .ZN(n712) );
  NAND2_X1 U659 ( .A1(n569), .A2(n712), .ZN(n570) );
  XOR2_X1 U660 ( .A(KEYINPUT90), .B(n570), .Z(n571) );
  NOR2_X1 U661 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U662 ( .A(KEYINPUT0), .ZN(n575) );
  INV_X1 U663 ( .A(n598), .ZN(n578) );
  NOR2_X1 U664 ( .A1(n596), .A2(n606), .ZN(n580) );
  XNOR2_X1 U665 ( .A(n580), .B(KEYINPUT94), .ZN(n657) );
  INV_X1 U666 ( .A(n347), .ZN(n581) );
  NAND2_X1 U667 ( .A1(n657), .A2(n581), .ZN(n584) );
  XOR2_X1 U668 ( .A(KEYINPUT96), .B(KEYINPUT31), .Z(n582) );
  XNOR2_X1 U669 ( .A(KEYINPUT95), .B(n582), .ZN(n583) );
  XNOR2_X1 U670 ( .A(n584), .B(n583), .ZN(n632) );
  NOR2_X1 U671 ( .A1(n348), .A2(n632), .ZN(n585) );
  XNOR2_X1 U672 ( .A(n585), .B(KEYINPUT97), .ZN(n587) );
  INV_X1 U673 ( .A(n662), .ZN(n586) );
  INV_X1 U674 ( .A(n647), .ZN(n594) );
  OR2_X1 U675 ( .A1(n667), .A2(n588), .ZN(n589) );
  NAND2_X1 U676 ( .A1(n607), .A2(n603), .ZN(n592) );
  XNOR2_X1 U677 ( .A(KEYINPUT86), .B(n592), .ZN(n593) );
  NOR2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n344), .A2(n595), .ZN(n616) );
  NOR2_X1 U680 ( .A1(n596), .A2(n603), .ZN(n597) );
  XOR2_X1 U681 ( .A(KEYINPUT73), .B(KEYINPUT34), .Z(n599) );
  XOR2_X1 U682 ( .A(KEYINPUT65), .B(KEYINPUT32), .Z(n605) );
  NOR2_X1 U683 ( .A1(n344), .A2(n647), .ZN(n602) );
  AND2_X1 U684 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  NOR2_X1 U686 ( .A1(n647), .A2(n608), .ZN(n609) );
  NAND2_X1 U687 ( .A1(n344), .A2(n609), .ZN(n623) );
  NAND2_X1 U688 ( .A1(n611), .A2(KEYINPUT2), .ZN(n612) );
  XOR2_X1 U689 ( .A(KEYINPUT67), .B(n612), .Z(n613) );
  NAND2_X1 U690 ( .A1(n359), .A2(KEYINPUT2), .ZN(n693) );
  AND2_X2 U691 ( .A1(n694), .A2(n693), .ZN(n690) );
  XNOR2_X1 U692 ( .A(G101), .B(n616), .ZN(G3) );
  NAND2_X1 U693 ( .A1(n348), .A2(n342), .ZN(n617) );
  XNOR2_X1 U694 ( .A(n617), .B(G104), .ZN(G6) );
  XOR2_X1 U695 ( .A(KEYINPUT114), .B(KEYINPUT27), .Z(n619) );
  XNOR2_X1 U696 ( .A(G107), .B(KEYINPUT26), .ZN(n618) );
  XNOR2_X1 U697 ( .A(n619), .B(n618), .ZN(n620) );
  XOR2_X1 U698 ( .A(KEYINPUT113), .B(n620), .Z(n622) );
  NAND2_X1 U699 ( .A1(n348), .A2(n633), .ZN(n621) );
  XNOR2_X1 U700 ( .A(n622), .B(n621), .ZN(G9) );
  XNOR2_X1 U701 ( .A(G110), .B(n623), .ZN(G12) );
  INV_X1 U702 ( .A(n633), .ZN(n624) );
  NOR2_X1 U703 ( .A1(n624), .A2(n628), .ZN(n626) );
  XNOR2_X1 U704 ( .A(G128), .B(KEYINPUT29), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n626), .B(n625), .ZN(G30) );
  XOR2_X1 U706 ( .A(G143), .B(n627), .Z(G45) );
  NOR2_X1 U707 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U708 ( .A(G146), .B(n630), .Z(G48) );
  NAND2_X1 U709 ( .A1(n632), .A2(n342), .ZN(n631) );
  XNOR2_X1 U710 ( .A(n631), .B(G113), .ZN(G15) );
  XOR2_X1 U711 ( .A(G116), .B(KEYINPUT115), .Z(n635) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U713 ( .A(n635), .B(n634), .ZN(G18) );
  XOR2_X1 U714 ( .A(G125), .B(KEYINPUT37), .Z(n636) );
  XNOR2_X1 U715 ( .A(n637), .B(n636), .ZN(G27) );
  XNOR2_X1 U716 ( .A(G134), .B(n638), .ZN(G36) );
  XOR2_X1 U717 ( .A(G140), .B(n354), .Z(G42) );
  INV_X1 U718 ( .A(KEYINPUT2), .ZN(n640) );
  AND2_X1 U719 ( .A1(n640), .A2(n726), .ZN(n639) );
  XNOR2_X1 U720 ( .A(n639), .B(KEYINPUT83), .ZN(n642) );
  NAND2_X1 U721 ( .A1(n640), .A2(n345), .ZN(n641) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n644) );
  NOR2_X1 U723 ( .A1(n647), .A2(n646), .ZN(n648) );
  XNOR2_X1 U724 ( .A(KEYINPUT49), .B(n648), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n649), .A2(n344), .ZN(n650) );
  XNOR2_X1 U726 ( .A(n650), .B(KEYINPUT50), .ZN(n651) );
  XNOR2_X1 U727 ( .A(KEYINPUT116), .B(n651), .ZN(n652) );
  NAND2_X1 U728 ( .A1(n653), .A2(n652), .ZN(n654) );
  NOR2_X1 U729 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U730 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U731 ( .A(KEYINPUT51), .B(n658), .ZN(n659) );
  NAND2_X1 U732 ( .A1(n659), .A2(n677), .ZN(n660) );
  XNOR2_X1 U733 ( .A(n660), .B(KEYINPUT117), .ZN(n673) );
  NOR2_X1 U734 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U735 ( .A(KEYINPUT119), .B(n663), .Z(n670) );
  NOR2_X1 U736 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U738 ( .A(KEYINPUT118), .B(n668), .ZN(n669) );
  NOR2_X1 U739 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U740 ( .A1(n679), .A2(n671), .ZN(n672) );
  NOR2_X1 U741 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U742 ( .A(n674), .B(KEYINPUT52), .ZN(n675) );
  NOR2_X1 U743 ( .A1(n676), .A2(n675), .ZN(n681) );
  INV_X1 U744 ( .A(n677), .ZN(n678) );
  NOR2_X1 U745 ( .A1(n679), .A2(n678), .ZN(n680) );
  NOR2_X1 U746 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U747 ( .A(KEYINPUT88), .B(KEYINPUT55), .Z(n685) );
  XNOR2_X1 U748 ( .A(n683), .B(KEYINPUT54), .ZN(n684) );
  XOR2_X1 U749 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n689) );
  XNOR2_X1 U750 ( .A(n687), .B(KEYINPUT120), .ZN(n688) );
  XNOR2_X1 U751 ( .A(n689), .B(n688), .ZN(n692) );
  NAND2_X1 U752 ( .A1(n702), .A2(G469), .ZN(n691) );
  NAND2_X1 U753 ( .A1(n695), .A2(n360), .ZN(n698) );
  INV_X1 U754 ( .A(KEYINPUT59), .ZN(n696) );
  XNOR2_X1 U755 ( .A(KEYINPUT60), .B(n699), .ZN(G60) );
  NAND2_X1 U756 ( .A1(G478), .A2(n702), .ZN(n700) );
  NAND2_X1 U757 ( .A1(G217), .A2(n702), .ZN(n703) );
  NAND2_X1 U758 ( .A1(n712), .A2(G953), .ZN(n707) );
  NAND2_X1 U759 ( .A1(n707), .A2(n706), .ZN(n708) );
  XNOR2_X1 U760 ( .A(n708), .B(KEYINPUT124), .ZN(n719) );
  NAND2_X1 U761 ( .A1(G224), .A2(G953), .ZN(n709) );
  XNOR2_X1 U762 ( .A(n709), .B(KEYINPUT61), .ZN(n710) );
  XNOR2_X1 U763 ( .A(n710), .B(KEYINPUT121), .ZN(n711) );
  NOR2_X1 U764 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U765 ( .A(n713), .B(KEYINPUT122), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n345), .A2(G953), .ZN(n715) );
  NOR2_X1 U767 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U768 ( .A(n717), .B(KEYINPUT123), .Z(n718) );
  XNOR2_X1 U769 ( .A(n719), .B(n718), .ZN(G69) );
  XOR2_X1 U770 ( .A(n720), .B(n721), .Z(n722) );
  XOR2_X1 U771 ( .A(KEYINPUT125), .B(n722), .Z(n727) );
  XOR2_X1 U772 ( .A(KEYINPUT126), .B(n727), .Z(n723) );
  XNOR2_X1 U773 ( .A(G227), .B(n723), .ZN(n724) );
  NAND2_X1 U774 ( .A1(n724), .A2(G900), .ZN(n725) );
  NAND2_X1 U775 ( .A1(n725), .A2(G953), .ZN(n731) );
  XOR2_X1 U776 ( .A(n727), .B(n726), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U778 ( .A1(n731), .A2(n730), .ZN(G72) );
  XOR2_X1 U779 ( .A(G122), .B(n343), .Z(G24) );
  XNOR2_X1 U780 ( .A(G137), .B(n733), .ZN(G39) );
  XNOR2_X1 U781 ( .A(G131), .B(n734), .ZN(G33) );
endmodule

