//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n733, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n835,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n894, new_n895, new_n896, new_n897, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941;
  INV_X1    g000(.A(G29gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(KEYINPUT14), .ZN(new_n203));
  INV_X1    g002(.A(G36gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n204), .B1(new_n202), .B2(KEYINPUT14), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n203), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(G43gat), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(G50gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT89), .B(G50gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(new_n209), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n210), .B1(new_n212), .B2(KEYINPUT90), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(KEYINPUT90), .B2(new_n212), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT15), .ZN(new_n215));
  AOI21_X1  g014(.A(new_n208), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G43gat), .B(G50gat), .Z(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(KEYINPUT88), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(KEYINPUT88), .ZN(new_n219));
  NOR3_X1   g018(.A1(new_n218), .A2(new_n219), .A3(new_n215), .ZN(new_n220));
  OR2_X1    g019(.A1(new_n216), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(new_n208), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  OR2_X1    g023(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(KEYINPUT17), .ZN(new_n226));
  NAND2_X1  g025(.A1(G85gat), .A2(G92gat), .ZN(new_n227));
  XNOR2_X1  g026(.A(new_n227), .B(KEYINPUT7), .ZN(new_n228));
  NAND2_X1  g027(.A1(G99gat), .A2(G106gat), .ZN(new_n229));
  INV_X1    g028(.A(G85gat), .ZN(new_n230));
  INV_X1    g029(.A(G92gat), .ZN(new_n231));
  AOI22_X1  g030(.A1(KEYINPUT8), .A2(new_n229), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G99gat), .B(G106gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n225), .A2(new_n226), .A3(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT41), .ZN(new_n238));
  NAND2_X1  g037(.A1(G232gat), .A2(G233gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT96), .Z(new_n240));
  OAI221_X1 g039(.A(new_n237), .B1(new_n238), .B2(new_n240), .C1(new_n224), .C2(new_n236), .ZN(new_n241));
  XNOR2_X1  g040(.A(G190gat), .B(G218gat), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n240), .A2(new_n238), .ZN(new_n244));
  XOR2_X1   g043(.A(G134gat), .B(G162gat), .Z(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n246), .A2(KEYINPUT97), .ZN(new_n247));
  OR2_X1    g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g047(.A1(new_n246), .A2(KEYINPUT97), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n243), .B1(new_n249), .B2(new_n247), .ZN(new_n250));
  AND2_X1   g049(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  XNOR2_X1  g050(.A(G15gat), .B(G22gat), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT16), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(G1gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n254), .B1(G1gat), .B2(new_n252), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n255), .B(G8gat), .Z(new_n256));
  INV_X1    g055(.A(KEYINPUT21), .ZN(new_n257));
  AOI21_X1  g056(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n258));
  AND2_X1   g057(.A1(G57gat), .A2(G64gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(G57gat), .A2(G64gat), .ZN(new_n260));
  OR3_X1    g059(.A1(new_n258), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(G71gat), .A2(G78gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT9), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n262), .B1(new_n263), .B2(KEYINPUT93), .ZN(new_n264));
  NOR2_X1   g063(.A1(G71gat), .A2(G78gat), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  OR2_X1    g065(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n261), .A2(new_n266), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n256), .B1(new_n257), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT95), .ZN(new_n271));
  NAND2_X1  g070(.A1(G231gat), .A2(G233gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(KEYINPUT94), .ZN(new_n273));
  XOR2_X1   g072(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n271), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n257), .ZN(new_n277));
  XOR2_X1   g076(.A(G127gat), .B(G155gat), .Z(new_n278));
  XNOR2_X1  g077(.A(new_n277), .B(new_n278), .ZN(new_n279));
  XOR2_X1   g078(.A(G183gat), .B(G211gat), .Z(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n276), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n251), .A2(KEYINPUT98), .A3(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT98), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n248), .A2(new_n250), .ZN(new_n285));
  INV_X1    g084(.A(new_n282), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n283), .A2(new_n287), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n235), .B(new_n269), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT10), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n235), .A2(KEYINPUT10), .A3(new_n267), .A4(new_n268), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g092(.A1(G230gat), .A2(G233gat), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n289), .A2(new_n294), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(G120gat), .B(G148gat), .Z(new_n298));
  XNOR2_X1  g097(.A(G176gat), .B(G204gat), .ZN(new_n299));
  XNOR2_X1  g098(.A(new_n298), .B(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g100(.A(new_n301), .B(KEYINPUT99), .Z(new_n302));
  NOR2_X1   g101(.A1(new_n297), .A2(new_n300), .ZN(new_n303));
  XNOR2_X1  g102(.A(new_n303), .B(KEYINPUT100), .ZN(new_n304));
  AND2_X1   g103(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT101), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g106(.A1(new_n302), .A2(new_n306), .A3(new_n304), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n288), .A2(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(G113gat), .B(G141gat), .ZN(new_n312));
  XNOR2_X1  g111(.A(new_n312), .B(G197gat), .ZN(new_n313));
  XOR2_X1   g112(.A(KEYINPUT11), .B(G169gat), .Z(new_n314));
  XNOR2_X1  g113(.A(new_n313), .B(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n315), .B(KEYINPUT12), .Z(new_n316));
  INV_X1    g115(.A(new_n224), .ZN(new_n317));
  INV_X1    g116(.A(new_n256), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n319), .B(KEYINPUT91), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n225), .A2(new_n256), .A3(new_n226), .ZN(new_n321));
  AND2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G229gat), .A2(G233gat), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n322), .A2(KEYINPUT18), .A3(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  XOR2_X1   g124(.A(new_n323), .B(KEYINPUT13), .Z(new_n326));
  NAND2_X1  g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT18), .B1(new_n322), .B2(new_n323), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n316), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n322), .A2(new_n323), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT18), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n316), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n333), .A2(new_n334), .A3(new_n324), .A4(new_n327), .ZN(new_n335));
  AND3_X1   g134(.A1(new_n330), .A2(KEYINPUT92), .A3(new_n335), .ZN(new_n336));
  AOI21_X1  g135(.A(KEYINPUT92), .B1(new_n330), .B2(new_n335), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(G183gat), .A2(G190gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(G169gat), .A2(G176gat), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n340), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n340), .A2(KEYINPUT67), .ZN(new_n342));
  INV_X1    g141(.A(KEYINPUT26), .ZN(new_n343));
  INV_X1    g142(.A(G169gat), .ZN(new_n344));
  INV_X1    g143(.A(G176gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n343), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n339), .B(new_n341), .C1(new_n342), .C2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT28), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT66), .B(G190gat), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT27), .B(G183gat), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n350), .A2(new_n351), .A3(new_n349), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n348), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  AND2_X1   g154(.A1(G169gat), .A2(G176gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(KEYINPUT23), .B2(new_n340), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n360));
  INV_X1    g159(.A(G183gat), .ZN(new_n361));
  INV_X1    g160(.A(G190gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n359), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT64), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n365), .B(new_n366), .C1(G169gat), .C2(G176gat), .ZN(new_n367));
  OAI21_X1  g166(.A(KEYINPUT64), .B1(new_n340), .B2(KEYINPUT23), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n357), .A2(new_n364), .A3(new_n367), .A4(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT25), .ZN(new_n370));
  AND2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  OR2_X1    g170(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n372));
  NAND2_X1  g171(.A1(KEYINPUT65), .A2(KEYINPUT24), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n372), .A2(new_n339), .A3(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n362), .A2(KEYINPUT66), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT66), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(G190gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n377), .A3(new_n361), .ZN(new_n378));
  AND3_X1   g177(.A1(new_n374), .A2(new_n378), .A3(new_n360), .ZN(new_n379));
  NAND4_X1  g178(.A1(new_n357), .A2(KEYINPUT25), .A3(new_n367), .A4(new_n368), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n355), .B1(new_n371), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(G113gat), .ZN(new_n383));
  INV_X1    g182(.A(G120gat), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT1), .ZN(new_n386));
  NAND2_X1  g185(.A1(G113gat), .A2(G120gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n385), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  AND2_X1   g187(.A1(G127gat), .A2(G134gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(G127gat), .A2(G134gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT69), .ZN(new_n393));
  AND2_X1   g192(.A1(G113gat), .A2(G120gat), .ZN(new_n394));
  NOR2_X1   g193(.A1(G113gat), .A2(G120gat), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n385), .A2(KEYINPUT69), .A3(new_n387), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n396), .A2(new_n397), .A3(new_n386), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT68), .B(G127gat), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n390), .B1(new_n399), .B2(G134gat), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n392), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n382), .A2(new_n401), .ZN(new_n402));
  AND2_X1   g201(.A1(new_n357), .A2(new_n368), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n374), .A2(new_n378), .A3(new_n360), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n403), .A2(KEYINPUT25), .A3(new_n367), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n369), .A2(new_n370), .ZN(new_n406));
  AND3_X1   g205(.A1(new_n350), .A2(new_n351), .A3(new_n349), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n352), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n405), .A2(new_n406), .B1(new_n408), .B2(new_n348), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n398), .A2(new_n400), .ZN(new_n410));
  INV_X1    g209(.A(new_n392), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n402), .A2(new_n413), .A3(G227gat), .A4(G233gat), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT32), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n415), .B1(new_n419), .B2(KEYINPUT33), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n415), .A2(KEYINPUT33), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n414), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT70), .B1(new_n423), .B2(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT70), .ZN(new_n425));
  AOI211_X1 g224(.A(new_n425), .B(new_n418), .C1(new_n414), .C2(new_n422), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n421), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n402), .A2(new_n413), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT34), .ZN(new_n429));
  NAND2_X1  g228(.A1(G227gat), .A2(G233gat), .ZN(new_n430));
  AND3_X1   g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n433), .B(new_n421), .C1(new_n424), .C2(new_n426), .ZN(new_n436));
  AND3_X1   g235(.A1(new_n435), .A2(KEYINPUT36), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT36), .B1(new_n435), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(G22gat), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT73), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT72), .ZN(new_n442));
  INV_X1    g241(.A(G204gat), .ZN(new_n443));
  NAND2_X1  g242(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(KEYINPUT71), .A2(G197gat), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n443), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT71), .ZN(new_n448));
  INV_X1    g247(.A(G197gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n450), .A2(G204gat), .A3(new_n444), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n447), .A2(new_n451), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n442), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  AOI211_X1 g254(.A(KEYINPUT72), .B(new_n453), .C1(new_n447), .C2(new_n451), .ZN(new_n456));
  XNOR2_X1  g255(.A(G211gat), .B(G218gat), .ZN(new_n457));
  NOR3_X1   g256(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n457), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n445), .A2(new_n446), .A3(new_n443), .ZN(new_n460));
  AOI21_X1  g259(.A(G204gat), .B1(new_n450), .B2(new_n444), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n454), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT72), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n452), .A2(new_n442), .A3(new_n454), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n441), .B1(new_n458), .B2(new_n465), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n457), .B1(new_n455), .B2(new_n456), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n463), .A2(new_n459), .A3(new_n464), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT73), .ZN(new_n469));
  NAND2_X1  g268(.A1(G155gat), .A2(G162gat), .ZN(new_n470));
  INV_X1    g269(.A(G155gat), .ZN(new_n471));
  INV_X1    g270(.A(G162gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  XNOR2_X1  g272(.A(G141gat), .B(G148gat), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n470), .B(new_n473), .C1(new_n474), .C2(KEYINPUT2), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT3), .ZN(new_n476));
  INV_X1    g275(.A(G141gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(G148gat), .ZN(new_n478));
  INV_X1    g277(.A(G148gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n479), .A2(G141gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n473), .A2(new_n470), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n470), .A2(KEYINPUT2), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n475), .A2(new_n476), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT29), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n466), .A2(new_n469), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n475), .A2(new_n484), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT29), .B1(new_n467), .B2(new_n468), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n489), .B1(new_n490), .B2(KEYINPUT3), .ZN(new_n491));
  INV_X1    g290(.A(G228gat), .ZN(new_n492));
  INV_X1    g291(.A(G233gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n488), .A2(new_n491), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n467), .A2(new_n468), .A3(new_n487), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n440), .B(new_n495), .C1(new_n497), .C2(new_n494), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  XNOR2_X1  g299(.A(G78gat), .B(G106gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT31), .B(G50gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n501), .B(new_n502), .ZN(new_n503));
  INV_X1    g302(.A(new_n495), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n494), .B1(new_n491), .B2(new_n496), .ZN(new_n505));
  OAI21_X1  g304(.A(G22gat), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n500), .A2(new_n503), .B1(new_n498), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n506), .A2(new_n498), .A3(KEYINPUT82), .A4(new_n503), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT75), .ZN(new_n511));
  NAND2_X1  g310(.A1(G226gat), .A2(G233gat), .ZN(new_n512));
  OAI211_X1 g311(.A(new_n355), .B(new_n512), .C1(new_n371), .C2(new_n381), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT29), .B1(G226gat), .B2(G233gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n409), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT74), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n515), .A2(new_n516), .A3(new_n469), .A4(new_n466), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n467), .A2(new_n468), .ZN(new_n518));
  OAI211_X1 g317(.A(new_n518), .B(new_n513), .C1(new_n409), .C2(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  AND3_X1   g319(.A1(new_n467), .A2(new_n468), .A3(KEYINPUT73), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT73), .B1(new_n467), .B2(new_n468), .ZN(new_n522));
  NOR2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n516), .B1(new_n523), .B2(new_n515), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n511), .B1(new_n520), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n515), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n466), .A2(new_n469), .ZN(new_n527));
  OAI21_X1  g326(.A(KEYINPUT74), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n528), .A2(KEYINPUT75), .A3(new_n517), .A4(new_n519), .ZN(new_n529));
  XNOR2_X1  g328(.A(G8gat), .B(G36gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(G64gat), .B(G92gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n529), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT76), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT76), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n525), .A2(new_n529), .A3(new_n536), .A4(new_n533), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n528), .A2(new_n517), .A3(new_n519), .A4(new_n532), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n520), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(KEYINPUT30), .A3(new_n528), .A4(new_n532), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n538), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g345(.A(G1gat), .B(G29gat), .Z(new_n547));
  XNOR2_X1  g346(.A(G57gat), .B(G85gat), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n489), .A2(KEYINPUT3), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n412), .A2(new_n553), .A3(new_n485), .ZN(new_n554));
  NAND2_X1  g353(.A1(G225gat), .A2(G233gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n556), .A2(KEYINPUT5), .ZN(new_n557));
  AND3_X1   g356(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n482), .B1(new_n483), .B2(new_n481), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT4), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n401), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n401), .B2(new_n560), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n554), .B(new_n557), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT5), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n554), .A2(new_n555), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT77), .ZN(new_n569));
  AOI211_X1 g368(.A(new_n569), .B(new_n561), .C1(new_n401), .C2(new_n560), .ZN(new_n570));
  NOR2_X1   g369(.A1(new_n568), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n564), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n569), .A3(new_n562), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n567), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n412), .A2(new_n489), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n401), .A2(new_n560), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n556), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT78), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n577), .A2(KEYINPUT78), .A3(new_n556), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n566), .B1(new_n574), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT83), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n552), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NOR3_X1   g384(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT77), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n576), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n587), .A2(new_n555), .A3(new_n554), .ZN(new_n588));
  OAI21_X1  g387(.A(KEYINPUT5), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT78), .B1(new_n577), .B2(new_n556), .ZN(new_n590));
  AOI211_X1 g389(.A(new_n579), .B(new_n555), .C1(new_n575), .C2(new_n576), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n565), .B1(new_n589), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(KEYINPUT83), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n585), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n554), .B1(new_n563), .B2(new_n564), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(new_n556), .ZN(new_n597));
  OAI211_X1 g396(.A(new_n597), .B(KEYINPUT39), .C1(new_n556), .C2(new_n577), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n598), .B(new_n551), .C1(KEYINPUT39), .C2(new_n597), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n599), .A2(KEYINPUT40), .ZN(new_n600));
  OR2_X1    g399(.A1(new_n599), .A2(KEYINPUT40), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n595), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n510), .B1(new_n546), .B2(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(KEYINPUT85), .B(KEYINPUT37), .ZN(new_n604));
  NAND4_X1  g403(.A1(new_n528), .A2(new_n517), .A3(new_n519), .A4(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(KEYINPUT86), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT86), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n542), .A2(new_n607), .A3(new_n528), .A4(new_n604), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n525), .A2(new_n529), .A3(KEYINPUT37), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n533), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT38), .ZN(new_n612));
  INV_X1    g411(.A(new_n539), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n532), .B1(new_n606), .B2(new_n608), .ZN(new_n614));
  INV_X1    g413(.A(KEYINPUT37), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n615), .B1(new_n523), .B2(new_n526), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n515), .A2(new_n518), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT38), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n613), .B1(new_n614), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n593), .A2(new_n552), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT6), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n551), .B(new_n565), .C1(new_n589), .C2(new_n592), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n623), .A2(new_n621), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n551), .B1(new_n593), .B2(KEYINPUT83), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n583), .A2(new_n584), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n622), .B1(new_n627), .B2(KEYINPUT84), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT84), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n595), .B2(new_n624), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n612), .A2(new_n619), .A3(new_n628), .A4(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n439), .B1(new_n603), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT80), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n620), .A2(new_n633), .A3(new_n621), .A4(new_n623), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n593), .B(new_n552), .C1(KEYINPUT80), .C2(KEYINPUT6), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AND4_X1   g435(.A1(KEYINPUT81), .A2(new_n538), .A3(new_n636), .A4(new_n545), .ZN(new_n637));
  AOI21_X1  g436(.A(new_n544), .B1(new_n535), .B2(new_n537), .ZN(new_n638));
  AOI21_X1  g437(.A(KEYINPUT81), .B1(new_n638), .B2(new_n636), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n510), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT87), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n500), .A2(new_n503), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n506), .A2(new_n498), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n645), .A2(new_n508), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n435), .A2(new_n436), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n646), .A2(new_n638), .A3(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT35), .ZN(new_n650));
  AOI21_X1  g449(.A(KEYINPUT6), .B1(new_n583), .B2(new_n551), .ZN(new_n651));
  OAI211_X1 g450(.A(KEYINPUT84), .B(new_n651), .C1(new_n585), .C2(new_n594), .ZN(new_n652));
  INV_X1    g451(.A(new_n622), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n625), .A2(new_n626), .ZN(new_n655));
  AOI21_X1  g454(.A(KEYINPUT84), .B1(new_n655), .B2(new_n651), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n650), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n642), .B1(new_n649), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT35), .B1(new_n628), .B2(new_n630), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n647), .B1(new_n645), .B2(new_n508), .ZN(new_n660));
  NAND4_X1  g459(.A1(new_n659), .A2(KEYINPUT87), .A3(new_n638), .A4(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n648), .ZN(new_n662));
  NOR3_X1   g461(.A1(new_n637), .A2(new_n639), .A3(new_n662), .ZN(new_n663));
  OAI211_X1 g462(.A(new_n658), .B(new_n661), .C1(new_n663), .C2(new_n650), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n338), .B1(new_n641), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n311), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n636), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n546), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT42), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT102), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AND2_X1   g476(.A1(new_n675), .A2(new_n676), .ZN(new_n678));
  AND2_X1   g477(.A1(new_n671), .A2(G8gat), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n673), .B1(new_n679), .B2(new_n674), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n677), .B1(new_n678), .B2(new_n680), .ZN(G1325gat));
  XNOR2_X1  g480(.A(new_n439), .B(KEYINPUT103), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(G15gat), .B1(new_n666), .B2(new_n683), .ZN(new_n684));
  OR2_X1    g483(.A1(new_n647), .A2(G15gat), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n684), .B1(new_n666), .B2(new_n685), .ZN(G1326gat));
  NOR2_X1   g485(.A1(new_n666), .A2(new_n646), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT104), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  XOR2_X1   g489(.A(KEYINPUT106), .B(KEYINPUT44), .Z(new_n691));
  AOI211_X1 g490(.A(new_n251), .B(new_n691), .C1(new_n664), .C2(new_n641), .ZN(new_n692));
  NOR2_X1   g491(.A1(KEYINPUT106), .A2(KEYINPUT44), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n637), .A2(new_n639), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n650), .B1(new_n694), .B2(new_n660), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n658), .A2(new_n661), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n641), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n693), .B1(new_n697), .B2(new_n285), .ZN(new_n698));
  OR2_X1    g497(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n309), .A2(new_n286), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n330), .A2(new_n335), .ZN(new_n701));
  INV_X1    g500(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n700), .A2(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g504(.A(G29gat), .B1(new_n705), .B2(new_n636), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n700), .A2(new_n251), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n665), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n708), .A2(G29gat), .A3(new_n636), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT105), .B(KEYINPUT45), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n706), .A2(new_n711), .ZN(G1328gat));
  NAND2_X1  g511(.A1(new_n546), .A2(new_n204), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT107), .ZN(new_n714));
  OAI22_X1  g513(.A1(new_n708), .A2(new_n713), .B1(new_n714), .B2(KEYINPUT46), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(KEYINPUT46), .ZN(new_n716));
  XOR2_X1   g515(.A(new_n715), .B(new_n716), .Z(new_n717));
  OAI21_X1  g516(.A(G36gat), .B1(new_n705), .B2(new_n638), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(G1329gat));
  NOR3_X1   g518(.A1(new_n708), .A2(G43gat), .A3(new_n647), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n682), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n721), .B2(G43gat), .ZN(new_n722));
  AOI21_X1  g521(.A(new_n209), .B1(new_n704), .B2(new_n439), .ZN(new_n723));
  INV_X1    g522(.A(new_n720), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(KEYINPUT47), .ZN(new_n725));
  OAI22_X1  g524(.A1(new_n722), .A2(KEYINPUT47), .B1(new_n723), .B2(new_n725), .ZN(G1330gat));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  INV_X1    g526(.A(new_n211), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n728), .B1(new_n704), .B2(new_n510), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n708), .A2(new_n211), .A3(new_n646), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n727), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT48), .ZN(G1331gat));
  NOR3_X1   g531(.A1(new_n288), .A2(new_n309), .A3(new_n701), .ZN(new_n733));
  AND2_X1   g532(.A1(new_n733), .A2(new_n697), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n668), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n546), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT49), .B(G64gat), .Z(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n737), .B2(new_n739), .ZN(G1333gat));
  AOI21_X1  g539(.A(G71gat), .B1(new_n734), .B2(new_n648), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n682), .A2(G71gat), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n741), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n510), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g545(.A1(new_n701), .A2(new_n282), .ZN(new_n747));
  INV_X1    g546(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n748), .A2(new_n309), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n699), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(G85gat), .B1(new_n750), .B2(new_n636), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT51), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n697), .A2(KEYINPUT109), .A3(new_n285), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n747), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n251), .B1(new_n664), .B2(new_n641), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(KEYINPUT109), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n752), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n697), .A2(new_n285), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n760), .A2(KEYINPUT51), .A3(new_n747), .A4(new_n753), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n757), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n310), .A2(new_n230), .A3(new_n668), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n751), .B1(new_n762), .B2(new_n763), .ZN(G1336gat));
  OAI21_X1  g563(.A(G92gat), .B1(new_n750), .B2(new_n638), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NOR3_X1   g565(.A1(new_n309), .A2(G92gat), .A3(new_n638), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n765), .B(new_n766), .C1(new_n762), .C2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n757), .A2(new_n761), .A3(KEYINPUT111), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT111), .ZN(new_n771));
  OAI211_X1 g570(.A(new_n771), .B(new_n752), .C1(new_n754), .C2(new_n756), .ZN(new_n772));
  XOR2_X1   g571(.A(new_n767), .B(KEYINPUT110), .Z(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n774), .A2(new_n765), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n769), .B1(new_n775), .B2(new_n766), .ZN(G1337gat));
  OAI21_X1  g575(.A(G99gat), .B1(new_n750), .B2(new_n683), .ZN(new_n777));
  OR3_X1    g576(.A1(new_n309), .A2(G99gat), .A3(new_n647), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n777), .B1(new_n762), .B2(new_n778), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(KEYINPUT112), .ZN(G1338gat));
  OAI211_X1 g579(.A(new_n510), .B(new_n749), .C1(new_n692), .C2(new_n698), .ZN(new_n781));
  AOI21_X1  g580(.A(KEYINPUT53), .B1(new_n781), .B2(G106gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n309), .A2(G106gat), .A3(new_n646), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n782), .B1(new_n762), .B2(new_n784), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT113), .ZN(new_n786));
  AND3_X1   g585(.A1(new_n781), .A2(new_n786), .A3(G106gat), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n786), .B1(new_n781), .B2(G106gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g588(.A(new_n783), .B(KEYINPUT114), .Z(new_n790));
  NAND3_X1  g589(.A1(new_n770), .A2(new_n772), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT115), .B1(new_n792), .B2(KEYINPUT53), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT115), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT53), .ZN(new_n795));
  AOI211_X1 g594(.A(new_n794), .B(new_n795), .C1(new_n789), .C2(new_n791), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n785), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  OAI211_X1 g598(.A(KEYINPUT116), .B(new_n785), .C1(new_n793), .C2(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n322), .A2(new_n323), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n325), .A2(new_n326), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n315), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n335), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n805), .B1(new_n307), .B2(new_n308), .ZN(new_n806));
  OR2_X1    g605(.A1(new_n293), .A2(new_n294), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n293), .A2(new_n294), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n807), .A2(KEYINPUT54), .A3(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT117), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n809), .B(new_n810), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT54), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n300), .B1(new_n295), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT55), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT118), .ZN(new_n817));
  XNOR2_X1  g616(.A(new_n816), .B(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n811), .A2(KEYINPUT55), .A3(new_n813), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n302), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n806), .B1(new_n821), .B2(new_n702), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n822), .A2(new_n251), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n818), .A2(new_n805), .A3(new_n285), .A4(new_n820), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n282), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n288), .A2(new_n701), .A3(new_n310), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR3_X1   g626(.A1(new_n827), .A2(new_n636), .A3(new_n649), .ZN(new_n828));
  AOI21_X1  g627(.A(G113gat), .B1(new_n828), .B2(new_n701), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n338), .A2(new_n383), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(G1340gat));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n310), .ZN(new_n832));
  XOR2_X1   g631(.A(KEYINPUT119), .B(G120gat), .Z(new_n833));
  XNOR2_X1  g632(.A(new_n832), .B(new_n833), .ZN(G1341gat));
  NAND2_X1  g633(.A1(new_n828), .A2(new_n282), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(new_n399), .ZN(G1342gat));
  INV_X1    g635(.A(G134gat), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n828), .A2(new_n837), .A3(new_n285), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(KEYINPUT56), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n837), .B1(new_n828), .B2(new_n285), .ZN(new_n841));
  OR3_X1    g640(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(G1343gat));
  NOR3_X1   g641(.A1(new_n439), .A2(new_n636), .A3(new_n546), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT120), .Z(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  XOR2_X1   g644(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n827), .B2(new_n646), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n820), .B(new_n816), .C1(new_n336), .C2(new_n337), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n285), .B1(new_n848), .B2(new_n806), .ZN(new_n849));
  INV_X1    g648(.A(new_n824), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n286), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  OAI211_X1 g651(.A(KEYINPUT57), .B(new_n510), .C1(new_n852), .C2(new_n826), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n845), .B1(new_n847), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n701), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n827), .A2(new_n636), .ZN(new_n856));
  AND4_X1   g655(.A1(new_n638), .A2(new_n856), .A3(new_n510), .A4(new_n683), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n338), .A2(G141gat), .ZN(new_n858));
  AOI22_X1  g657(.A1(new_n855), .A2(G141gat), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n857), .A2(new_n858), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n860), .ZN(new_n862));
  INV_X1    g661(.A(new_n338), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n477), .B1(new_n854), .B2(new_n863), .ZN(new_n864));
  OAI22_X1  g663(.A1(new_n859), .A2(new_n860), .B1(new_n862), .B2(new_n864), .ZN(G1344gat));
  NAND3_X1  g664(.A1(new_n857), .A2(new_n479), .A3(new_n310), .ZN(new_n866));
  INV_X1    g665(.A(new_n846), .ZN(new_n867));
  OAI211_X1 g666(.A(new_n510), .B(new_n867), .C1(new_n825), .C2(new_n826), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n311), .A2(new_n338), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n646), .B1(new_n851), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n868), .B1(new_n870), .B2(KEYINPUT57), .ZN(new_n871));
  INV_X1    g670(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n309), .B1(new_n845), .B2(KEYINPUT122), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(KEYINPUT122), .B2(new_n845), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT59), .B(G148gat), .C1(new_n872), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n479), .B1(new_n854), .B2(new_n310), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n866), .B(new_n875), .C1(new_n876), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g676(.A(G155gat), .B1(new_n857), .B2(new_n282), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n282), .A2(G155gat), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT123), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n878), .B1(new_n854), .B2(new_n880), .ZN(G1346gat));
  AOI21_X1  g680(.A(G162gat), .B1(new_n857), .B2(new_n285), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n251), .A2(new_n472), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n882), .B1(new_n854), .B2(new_n883), .ZN(G1347gat));
  NOR2_X1   g683(.A1(new_n827), .A2(new_n668), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n662), .A2(new_n638), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n344), .A3(new_n338), .ZN(new_n888));
  INV_X1    g687(.A(new_n887), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n701), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n888), .B1(new_n344), .B2(new_n890), .ZN(G1348gat));
  NOR2_X1   g690(.A1(new_n887), .A2(new_n309), .ZN(new_n892));
  XNOR2_X1  g691(.A(new_n892), .B(new_n345), .ZN(G1349gat));
  NAND3_X1  g692(.A1(new_n885), .A2(new_n282), .A3(new_n886), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n361), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n351), .B2(new_n894), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n897));
  XNOR2_X1  g696(.A(new_n896), .B(new_n897), .ZN(G1350gat));
  NAND3_X1  g697(.A1(new_n885), .A2(new_n285), .A3(new_n886), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G190gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT124), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT124), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n899), .A2(new_n902), .A3(G190gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n901), .A2(KEYINPUT61), .A3(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT61), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n900), .A2(KEYINPUT124), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n889), .A2(new_n350), .A3(new_n285), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n904), .A2(new_n906), .A3(new_n907), .ZN(G1351gat));
  NOR3_X1   g707(.A1(new_n682), .A2(new_n638), .A3(new_n646), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n885), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g709(.A(G197gat), .B1(new_n910), .B2(new_n701), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n638), .A2(new_n668), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n683), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n871), .A2(KEYINPUT125), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n868), .B(new_n915), .C1(new_n870), .C2(KEYINPUT57), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n913), .B1(new_n914), .B2(new_n916), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n338), .A2(new_n449), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n911), .B1(new_n917), .B2(new_n918), .ZN(G1352gat));
  XOR2_X1   g718(.A(KEYINPUT126), .B(G204gat), .Z(new_n920));
  NOR2_X1   g719(.A1(new_n309), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n910), .A2(new_n921), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT62), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n914), .A2(new_n916), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT127), .ZN(new_n926));
  INV_X1    g725(.A(new_n913), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n925), .A2(new_n926), .A3(new_n310), .A4(new_n927), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(new_n920), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n926), .B1(new_n917), .B2(new_n310), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n924), .B1(new_n929), .B2(new_n930), .ZN(G1353gat));
  INV_X1    g730(.A(G211gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n910), .A2(new_n932), .A3(new_n282), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n913), .A2(new_n286), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n932), .B1(new_n871), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g734(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G1354gat));
  INV_X1    g737(.A(G218gat), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n910), .A2(new_n939), .A3(new_n285), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n917), .A2(new_n285), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n941), .B2(new_n939), .ZN(G1355gat));
endmodule


