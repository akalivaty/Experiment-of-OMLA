//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 1 0 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n444, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n457, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n493, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n536, new_n538, new_n540, new_n541, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n601, new_n602,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n847, new_n848, new_n849, new_n850,
    new_n851, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  XNOR2_X1  g004(.A(KEYINPUT65), .B(G1083), .ZN(G367));
  XNOR2_X1  g005(.A(KEYINPUT66), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  XNOR2_X1  g013(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT68), .ZN(G259));
  XNOR2_X1  g020(.A(KEYINPUT69), .B(G452), .ZN(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT70), .ZN(G217));
  NAND4_X1  g027(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT2), .Z(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n456));
  INV_X1    g031(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n455), .A2(new_n457), .ZN(G325));
  XOR2_X1   g033(.A(G325), .B(KEYINPUT71), .Z(G261));
  AOI22_X1  g034(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n457), .ZN(G319));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g040(.A1(new_n465), .A2(G2105), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n461), .A2(G2105), .ZN(new_n467));
  AOI22_X1  g042(.A1(new_n466), .A2(G137), .B1(G101), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G125), .ZN(new_n470));
  OAI21_X1  g045(.A(new_n469), .B1(new_n465), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n468), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n465), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n466), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n477), .A2(new_n478), .A3(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(new_n462), .A2(new_n464), .ZN(new_n482));
  AND2_X1   g057(.A1(KEYINPUT72), .A2(G138), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n482), .A2(KEYINPUT4), .A3(new_n475), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n482), .A2(G126), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n475), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n462), .A2(new_n464), .A3(new_n483), .A4(new_n475), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n484), .A2(new_n485), .A3(new_n487), .A4(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G164));
  NAND2_X1  g067(.A1(KEYINPUT73), .A2(KEYINPUT5), .ZN(new_n493));
  INV_X1    g068(.A(G543), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND3_X1  g070(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  AOI22_X1  g072(.A1(new_n497), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  XNOR2_X1  g076(.A(KEYINPUT6), .B(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G543), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(KEYINPUT6), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(G651), .ZN(new_n506));
  AND3_X1   g081(.A1(KEYINPUT73), .A2(KEYINPUT5), .A3(G543), .ZN(new_n507));
  AOI21_X1  g082(.A(G543), .B1(KEYINPUT73), .B2(KEYINPUT5), .ZN(new_n508));
  OAI211_X1 g083(.A(new_n504), .B(new_n506), .C1(new_n507), .C2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT74), .B(G88), .ZN(new_n510));
  OAI22_X1  g085(.A1(new_n501), .A2(new_n503), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n500), .A2(new_n511), .ZN(G166));
  INV_X1    g087(.A(new_n509), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G89), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT75), .B(KEYINPUT7), .ZN(new_n515));
  AND3_X1   g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  XNOR2_X1  g091(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n504), .A2(new_n506), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n518), .A2(new_n494), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n519), .A2(G51), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n497), .A2(G63), .A3(G651), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n514), .A2(new_n517), .A3(new_n520), .A4(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n497), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n499), .ZN(new_n525));
  INV_X1    g100(.A(G52), .ZN(new_n526));
  INV_X1    g101(.A(G90), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n526), .A2(new_n503), .B1(new_n509), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  NAND4_X1  g104(.A1(new_n504), .A2(new_n506), .A3(G43), .A4(G543), .ZN(new_n530));
  INV_X1    g105(.A(G81), .ZN(new_n531));
  OAI21_X1  g106(.A(new_n530), .B1(new_n509), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g107(.A(G56), .B1(new_n507), .B2(new_n508), .ZN(new_n533));
  NAND2_X1  g108(.A1(G68), .A2(G543), .ZN(new_n534));
  AOI21_X1  g109(.A(new_n499), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n532), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G860), .ZN(G153));
  AND3_X1   g112(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G36), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n538), .A2(new_n541), .ZN(G188));
  NAND4_X1  g117(.A1(new_n504), .A2(new_n506), .A3(G53), .A4(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(KEYINPUT9), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT9), .ZN(new_n545));
  NAND4_X1  g120(.A1(new_n502), .A2(new_n545), .A3(G53), .A4(G543), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n497), .A2(G91), .A3(new_n502), .ZN(new_n548));
  INV_X1    g123(.A(G65), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n549), .B1(new_n495), .B2(new_n496), .ZN(new_n550));
  INV_X1    g125(.A(G78), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n551), .A2(new_n494), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n547), .A2(new_n548), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(KEYINPUT76), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g131(.A1(new_n547), .A2(KEYINPUT76), .A3(new_n553), .A4(new_n548), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(G299));
  INV_X1    g133(.A(G171), .ZN(G301));
  INV_X1    g134(.A(G166), .ZN(G303));
  NAND2_X1  g135(.A1(new_n513), .A2(G87), .ZN(new_n561));
  OAI21_X1  g136(.A(G651), .B1(new_n497), .B2(G74), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n519), .A2(G49), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n561), .A2(new_n562), .A3(new_n563), .ZN(G288));
  INV_X1    g139(.A(G48), .ZN(new_n565));
  INV_X1    g140(.A(G86), .ZN(new_n566));
  OAI22_X1  g141(.A1(new_n565), .A2(new_n503), .B1(new_n509), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n497), .A2(G61), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n499), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n568), .A2(new_n572), .ZN(G305));
  AOI22_X1  g148(.A1(new_n497), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n574), .A2(new_n499), .ZN(new_n575));
  INV_X1    g150(.A(G47), .ZN(new_n576));
  INV_X1    g151(.A(G85), .ZN(new_n577));
  OAI22_X1  g152(.A1(new_n576), .A2(new_n503), .B1(new_n509), .B2(new_n577), .ZN(new_n578));
  NOR2_X1   g153(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(G301), .A2(G868), .ZN(new_n581));
  INV_X1    g156(.A(G66), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n495), .B2(new_n496), .ZN(new_n583));
  NAND2_X1  g158(.A1(G79), .A2(G543), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT77), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n507), .A2(new_n508), .ZN(new_n588));
  OAI211_X1 g163(.A(new_n587), .B(new_n584), .C1(new_n588), .C2(new_n582), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n589), .A3(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  INV_X1    g166(.A(G92), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n509), .B2(new_n592), .ZN(new_n593));
  NAND4_X1  g168(.A1(new_n497), .A2(KEYINPUT10), .A3(new_n502), .A4(G92), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n519), .A2(G54), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n590), .A2(new_n595), .A3(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n581), .B1(G868), .B2(new_n598), .ZN(G321));
  XOR2_X1   g174(.A(G321), .B(KEYINPUT78), .Z(G284));
  NAND2_X1  g175(.A1(G286), .A2(G868), .ZN(new_n601));
  INV_X1    g176(.A(G299), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G297));
  OAI21_X1  g178(.A(new_n601), .B1(new_n602), .B2(G868), .ZN(G280));
  NOR2_X1   g179(.A1(new_n597), .A2(G559), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n598), .B2(G860), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT79), .Z(G148));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(new_n597), .B2(G559), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  NOR3_X1   g185(.A1(new_n597), .A2(new_n608), .A3(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(G868), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n612), .B1(G868), .B2(new_n536), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n476), .A2(G123), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n466), .A2(G135), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n475), .A2(G111), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n615), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  OR2_X1    g194(.A1(new_n619), .A2(KEYINPUT82), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(KEYINPUT82), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XOR2_X1   g197(.A(new_n622), .B(G2096), .Z(new_n623));
  NAND2_X1  g198(.A1(new_n482), .A2(new_n467), .ZN(new_n624));
  XOR2_X1   g199(.A(new_n624), .B(KEYINPUT12), .Z(new_n625));
  XOR2_X1   g200(.A(KEYINPUT81), .B(KEYINPUT13), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(G2100), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n625), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n623), .A2(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT84), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n634), .A2(G2438), .ZN(new_n635));
  OR2_X1    g210(.A1(new_n634), .A2(G2438), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n636), .A2(new_n635), .ZN(new_n638));
  INV_X1    g213(.A(KEYINPUT84), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n632), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n637), .A2(new_n641), .A3(KEYINPUT14), .ZN(new_n642));
  XOR2_X1   g217(.A(KEYINPUT83), .B(KEYINPUT16), .Z(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2443), .B(G2446), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(new_n646), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n643), .ZN(new_n649));
  NAND4_X1  g224(.A1(new_n637), .A2(new_n641), .A3(KEYINPUT14), .A4(new_n649), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n648), .A3(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  AOI21_X1  g227(.A(new_n648), .B1(new_n644), .B2(new_n650), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n631), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n653), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n655), .A2(new_n630), .A3(new_n651), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n654), .A2(new_n656), .A3(G14), .ZN(new_n657));
  INV_X1    g232(.A(KEYINPUT85), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g234(.A1(new_n654), .A2(new_n656), .A3(KEYINPUT85), .A4(G14), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XOR2_X1   g238(.A(G2067), .B(G2678), .Z(new_n664));
  XNOR2_X1  g239(.A(G2084), .B(G2090), .ZN(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n663), .B1(new_n666), .B2(KEYINPUT18), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT87), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT17), .ZN(new_n670));
  AOI22_X1  g245(.A1(new_n664), .A2(new_n665), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  OAI211_X1 g246(.A(new_n666), .B(new_n671), .C1(new_n669), .C2(new_n670), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n668), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G2096), .B(G2100), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(G227));
  XNOR2_X1  g253(.A(G1971), .B(G1976), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1956), .B(G2474), .Z(new_n682));
  XOR2_X1   g257(.A(G1961), .B(G1966), .Z(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT20), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n682), .A2(new_n683), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n681), .A2(new_n687), .ZN(new_n688));
  OR3_X1    g263(.A1(new_n681), .A2(new_n684), .A3(new_n687), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n686), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1991), .B(G1996), .ZN(new_n693));
  INV_X1    g268(.A(G1981), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n696), .ZN(G229));
  XNOR2_X1  g272(.A(KEYINPUT90), .B(G16), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G24), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n579), .B2(new_n699), .ZN(new_n701));
  INV_X1    g276(.A(G1986), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(G25), .A2(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n476), .A2(G119), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n466), .A2(G131), .ZN(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n475), .A2(G107), .ZN(new_n708));
  OAI211_X1 g283(.A(new_n705), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT89), .Z(new_n710));
  AOI21_X1  g285(.A(new_n704), .B1(new_n710), .B2(G29), .ZN(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT35), .B(G1991), .ZN(new_n712));
  INV_X1    g287(.A(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n711), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n699), .A2(G22), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G166), .B2(new_n699), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(G1971), .ZN(new_n717));
  OR2_X1    g292(.A1(G16), .A2(G23), .ZN(new_n718));
  INV_X1    g293(.A(G16), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(G288), .B2(new_n719), .ZN(new_n720));
  XOR2_X1   g295(.A(KEYINPUT33), .B(G1976), .Z(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n720), .A2(new_n722), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n717), .A2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n719), .A2(G6), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n727), .B1(G305), .B2(G16), .ZN(new_n728));
  XOR2_X1   g303(.A(KEYINPUT91), .B(G1981), .Z(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT32), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n728), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(new_n731), .ZN(new_n732));
  AOI21_X1  g307(.A(KEYINPUT34), .B1(new_n726), .B2(new_n732), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n716), .A2(G1971), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n716), .A2(G1971), .ZN(new_n735));
  NAND4_X1  g310(.A1(new_n734), .A2(new_n735), .A3(new_n723), .A4(new_n724), .ZN(new_n736));
  INV_X1    g311(.A(KEYINPUT34), .ZN(new_n737));
  NOR3_X1   g312(.A1(new_n736), .A2(new_n731), .A3(new_n737), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n703), .B(new_n714), .C1(new_n733), .C2(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n739), .A2(KEYINPUT36), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n726), .A2(new_n732), .A3(KEYINPUT34), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n737), .B1(new_n736), .B2(new_n731), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT36), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n743), .A2(new_n744), .A3(new_n703), .A4(new_n714), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n740), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g321(.A1(G16), .A2(G21), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n747), .B1(G168), .B2(G16), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n748), .A2(G1966), .ZN(new_n749));
  AND2_X1   g324(.A1(new_n748), .A2(G1966), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  NAND2_X1  g326(.A1(G171), .A2(G16), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G5), .B2(G16), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n749), .B(new_n750), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  OR2_X1    g329(.A1(G29), .A2(G32), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT27), .B(G1996), .Z(new_n756));
  NAND2_X1  g331(.A1(new_n466), .A2(G141), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n476), .A2(G129), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n467), .A2(G105), .ZN(new_n759));
  NAND3_X1  g334(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT26), .Z(new_n761));
  NAND4_X1  g336(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT96), .ZN(new_n763));
  AOI22_X1  g338(.A1(G129), .A2(new_n476), .B1(new_n466), .B2(G141), .ZN(new_n764));
  INV_X1    g339(.A(KEYINPUT96), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n764), .A2(new_n765), .A3(new_n759), .A4(new_n761), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  INV_X1    g342(.A(G29), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n755), .B(new_n756), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(G28), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(G28), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n771), .A2(new_n772), .A3(new_n768), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT95), .B(KEYINPUT25), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n467), .A2(G103), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(G115), .A2(G2104), .ZN(new_n777));
  INV_X1    g352(.A(G127), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n465), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G2105), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n466), .A2(G139), .ZN(new_n781));
  AND3_X1   g356(.A1(new_n776), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n782), .A2(G29), .ZN(new_n783));
  NOR2_X1   g358(.A1(G29), .A2(G33), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n783), .A2(G2072), .A3(new_n785), .ZN(new_n786));
  NAND3_X1  g361(.A1(new_n620), .A2(G29), .A3(new_n621), .ZN(new_n787));
  NAND4_X1  g362(.A1(new_n769), .A2(new_n773), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n699), .A2(G20), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT99), .B(KEYINPUT23), .Z(new_n790));
  XOR2_X1   g365(.A(new_n789), .B(new_n790), .Z(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OAI211_X1 g367(.A(G1956), .B(new_n792), .C1(new_n602), .C2(new_n719), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n792), .B1(new_n602), .B2(new_n719), .ZN(new_n794));
  INV_X1    g369(.A(G1956), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n788), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n798), .A2(new_n768), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G160), .B2(new_n768), .ZN(new_n801));
  XOR2_X1   g376(.A(new_n801), .B(G2084), .Z(new_n802));
  NOR2_X1   g377(.A1(G29), .A2(G35), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n803), .B1(G162), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT29), .B(G2090), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n755), .B1(new_n767), .B2(new_n768), .ZN(new_n807));
  INV_X1    g382(.A(new_n756), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n754), .A2(new_n797), .A3(new_n802), .A4(new_n809), .ZN(new_n810));
  AOI21_X1  g385(.A(G2072), .B1(new_n783), .B2(new_n785), .ZN(new_n811));
  INV_X1    g386(.A(G11), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n811), .B1(KEYINPUT31), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(KEYINPUT31), .B2(new_n812), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n753), .A2(new_n751), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n699), .A2(G19), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n536), .B2(new_n699), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(G1341), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n768), .A2(G27), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G164), .B2(new_n768), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT98), .ZN(new_n823));
  INV_X1    g398(.A(G2078), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR4_X1   g400(.A1(new_n810), .A2(new_n814), .A3(new_n820), .A4(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n719), .A2(G4), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n598), .B2(new_n719), .ZN(new_n828));
  INV_X1    g403(.A(G1348), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n823), .A2(new_n824), .ZN(new_n831));
  NAND4_X1  g406(.A1(new_n746), .A2(new_n826), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n768), .A2(G26), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(G116), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(G2105), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT92), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n476), .A2(G128), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n466), .A2(G140), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n835), .B1(new_n842), .B2(G29), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT94), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(G2067), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n832), .A2(new_n845), .ZN(G311));
  AND3_X1   g421(.A1(new_n746), .A2(new_n831), .A3(new_n826), .ZN(new_n847));
  INV_X1    g422(.A(new_n845), .ZN(new_n848));
  NAND4_X1  g423(.A1(new_n847), .A2(KEYINPUT100), .A3(new_n848), .A4(new_n830), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n850), .B1(new_n832), .B2(new_n845), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G150));
  NAND3_X1  g427(.A1(new_n502), .A2(G55), .A3(G543), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n497), .A2(G93), .A3(new_n502), .ZN(new_n854));
  NAND2_X1  g429(.A1(G80), .A2(G543), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n497), .B2(G67), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n853), .B(new_n854), .C1(new_n857), .C2(new_n499), .ZN(new_n858));
  XNOR2_X1  g433(.A(KEYINPUT105), .B(G860), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  XOR2_X1   g435(.A(new_n860), .B(KEYINPUT37), .Z(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n854), .A2(new_n853), .ZN(new_n863));
  OAI21_X1  g438(.A(G67), .B1(new_n507), .B2(new_n508), .ZN(new_n864));
  AOI21_X1  g439(.A(new_n499), .B1(new_n864), .B2(new_n855), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n497), .A2(G81), .A3(new_n502), .ZN(new_n867));
  INV_X1    g442(.A(new_n534), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n497), .B2(G56), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n530), .B(new_n867), .C1(new_n869), .C2(new_n499), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n862), .B1(new_n866), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n536), .A2(new_n858), .A3(KEYINPUT102), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g448(.A(KEYINPUT103), .B1(new_n536), .B2(new_n858), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT103), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n866), .A2(new_n875), .A3(new_n870), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n873), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT39), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n598), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT104), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n879), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(KEYINPUT101), .B(KEYINPUT38), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n882), .B(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n861), .B1(new_n884), .B2(new_n859), .ZN(G145));
  XNOR2_X1  g460(.A(new_n622), .B(new_n473), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT107), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n767), .B(new_n887), .ZN(new_n888));
  XOR2_X1   g463(.A(new_n782), .B(new_n842), .Z(new_n889));
  OR2_X1    g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g465(.A1(G130), .A2(new_n476), .B1(new_n466), .B2(G142), .ZN(new_n891));
  OAI21_X1  g466(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n475), .A2(G118), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT106), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n891), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(new_n709), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n625), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n888), .A2(new_n889), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n890), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(new_n897), .B1(new_n890), .B2(new_n898), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n886), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n901), .ZN(new_n903));
  INV_X1    g478(.A(new_n886), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n903), .A2(new_n899), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n902), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g481(.A(G164), .B(G162), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(G37), .ZN(new_n909));
  INV_X1    g484(.A(new_n907), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n902), .A2(new_n905), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n908), .A2(new_n909), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n912), .A2(KEYINPUT40), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT40), .ZN(new_n914));
  NAND4_X1  g489(.A1(new_n908), .A2(new_n914), .A3(new_n909), .A4(new_n911), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n915), .ZN(G395));
  INV_X1    g491(.A(new_n611), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n609), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n918), .B1(new_n917), .B2(new_n609), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n878), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n921), .ZN(new_n923));
  INV_X1    g498(.A(new_n878), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n923), .A2(new_n924), .A3(new_n919), .ZN(new_n925));
  NOR2_X1   g500(.A1(G299), .A2(new_n597), .ZN(new_n926));
  AND2_X1   g501(.A1(new_n590), .A2(new_n596), .ZN(new_n927));
  AOI22_X1  g502(.A1(new_n927), .A2(new_n595), .B1(new_n556), .B2(new_n557), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(new_n929), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n922), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(G299), .A2(new_n597), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT41), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n927), .A2(new_n556), .A3(new_n557), .A4(new_n595), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OR2_X1    g510(.A1(new_n935), .A2(KEYINPUT109), .ZN(new_n936));
  OAI21_X1  g511(.A(KEYINPUT41), .B1(new_n926), .B2(new_n928), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n937), .A2(KEYINPUT109), .A3(new_n935), .ZN(new_n938));
  AOI22_X1  g513(.A1(new_n922), .A2(new_n925), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  XOR2_X1   g514(.A(G305), .B(KEYINPUT110), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(G166), .B(G288), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n942), .A2(G290), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(G290), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n941), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  OR2_X1    g520(.A1(new_n942), .A2(G290), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n942), .A2(G290), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n946), .A2(new_n940), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT42), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n949), .B1(new_n945), .B2(new_n948), .ZN(new_n951));
  OAI22_X1  g526(.A1(new_n931), .A2(new_n939), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n950), .A2(new_n951), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n922), .A2(new_n925), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n938), .A2(new_n936), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n922), .A2(new_n925), .A3(new_n930), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n952), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(G868), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n866), .A2(G868), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n960), .A2(new_n962), .ZN(G295));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  AOI21_X1  g539(.A(new_n964), .B1(new_n960), .B2(new_n962), .ZN(new_n965));
  AOI211_X1 g540(.A(KEYINPUT111), .B(new_n961), .C1(new_n959), .C2(G868), .ZN(new_n966));
  NOR2_X1   g541(.A1(new_n965), .A2(new_n966), .ZN(G331));
  AND3_X1   g542(.A1(new_n873), .A2(new_n877), .A3(G301), .ZN(new_n968));
  AOI21_X1  g543(.A(G301), .B1(new_n873), .B2(new_n877), .ZN(new_n969));
  OAI21_X1  g544(.A(G286), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n878), .A2(G171), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n873), .A2(new_n877), .A3(G301), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(G168), .A3(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n970), .A2(new_n973), .A3(new_n929), .ZN(new_n974));
  AND2_X1   g549(.A1(new_n970), .A2(new_n973), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n974), .B1(new_n975), .B2(new_n955), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n945), .A2(new_n948), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT112), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n909), .ZN(new_n981));
  NOR3_X1   g556(.A1(new_n968), .A2(new_n969), .A3(G286), .ZN(new_n982));
  AOI21_X1  g557(.A(G168), .B1(new_n971), .B2(new_n972), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n936), .B(new_n938), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n977), .B1(new_n984), .B2(new_n974), .ZN(new_n985));
  OAI21_X1  g560(.A(KEYINPUT112), .B1(new_n985), .B2(G37), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n984), .A2(new_n977), .A3(new_n974), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n981), .A2(new_n986), .A3(KEYINPUT43), .A4(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT44), .ZN(new_n989));
  INV_X1    g564(.A(new_n974), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n970), .A2(new_n973), .B1(new_n935), .B2(new_n937), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n978), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n992), .A2(new_n987), .A3(new_n909), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT43), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n988), .A2(new_n989), .A3(new_n995), .ZN(new_n996));
  NOR2_X1   g571(.A1(new_n993), .A2(new_n994), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n981), .A2(new_n986), .A3(new_n987), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n998), .B2(new_n994), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n996), .B1(new_n999), .B2(new_n989), .ZN(G397));
  INV_X1    g575(.A(G1384), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n491), .A2(new_n1001), .ZN(new_n1002));
  XNOR2_X1  g577(.A(new_n1002), .B(KEYINPUT113), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(KEYINPUT45), .ZN(new_n1004));
  XNOR2_X1  g579(.A(KEYINPUT114), .B(G40), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n468), .A2(new_n472), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1004), .A2(new_n1008), .ZN(new_n1009));
  NOR3_X1   g584(.A1(new_n1009), .A2(new_n702), .A3(new_n579), .ZN(new_n1010));
  NOR3_X1   g585(.A1(new_n1009), .A2(G1986), .A3(G290), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g587(.A(new_n1012), .B(KEYINPUT115), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1009), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n767), .A2(G1996), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n842), .B(G2067), .ZN(new_n1016));
  INV_X1    g591(.A(G1996), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n763), .B2(new_n766), .ZN(new_n1018));
  NOR3_X1   g593(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1014), .A2(KEYINPUT116), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT116), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n1009), .B2(new_n1019), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n709), .B(new_n712), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1024), .B1(new_n1014), .B2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1013), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT45), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1002), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n491), .A2(KEYINPUT45), .A3(new_n1001), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1029), .A2(new_n1008), .A3(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT117), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT117), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n1029), .A2(new_n1033), .A3(new_n1008), .A4(new_n1030), .ZN(new_n1034));
  AOI21_X1  g609(.A(G1971), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1007), .B1(new_n1002), .B2(KEYINPUT50), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n491), .A2(new_n1037), .A3(new_n1001), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1036), .A2(new_n1038), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1039), .A2(G2090), .ZN(new_n1040));
  OAI21_X1  g615(.A(G8), .B1(new_n1035), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(G303), .A2(G8), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1042), .B(KEYINPUT55), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1041), .A2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1043), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1038), .A2(KEYINPUT118), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n491), .A2(new_n1047), .A3(new_n1037), .A4(new_n1001), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1036), .A2(new_n1046), .A3(new_n1048), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1049), .A2(G2090), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1045), .B(G8), .C1(new_n1035), .C2(new_n1050), .ZN(new_n1051));
  NOR3_X1   g626(.A1(new_n567), .A2(new_n571), .A3(G1981), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT119), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT49), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n568), .A2(new_n572), .A3(new_n694), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT49), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(KEYINPUT119), .A3(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(G305), .A2(G1981), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1002), .A2(new_n1007), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1054), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1061), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(G1976), .ZN(new_n1067));
  OAI221_X1 g642(.A(G8), .B1(G288), .B2(new_n1067), .C1(new_n1002), .C2(new_n1007), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT52), .ZN(new_n1069));
  INV_X1    g644(.A(G288), .ZN(new_n1070));
  NOR2_X1   g645(.A1(new_n1070), .A2(G1976), .ZN(new_n1071));
  OR3_X1    g646(.A1(new_n1068), .A2(KEYINPUT52), .A3(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1066), .A2(new_n1069), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1966), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1031), .A2(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(G2084), .B2(new_n1049), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1076), .A2(G8), .A3(G168), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1044), .A2(new_n1051), .A3(new_n1073), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT63), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(G8), .B1(new_n1035), .B2(new_n1050), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1079), .B1(new_n1081), .B2(new_n1043), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1082), .A2(new_n1051), .A3(new_n1073), .A4(new_n1077), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1080), .A2(new_n1083), .ZN(new_n1084));
  AND3_X1   g659(.A1(new_n1044), .A2(new_n1051), .A3(new_n1073), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT51), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1086), .B1(new_n1076), .B2(G286), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1075), .B(G168), .C1(G2084), .C2(new_n1049), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1086), .B1(new_n1088), .B2(G8), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT62), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1091), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT62), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(new_n1094), .C1(new_n1089), .C2(new_n1087), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1032), .A2(new_n824), .A3(new_n1034), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT53), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1096), .A2(new_n1097), .B1(new_n751), .B2(new_n1049), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1031), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1099), .A2(KEYINPUT53), .A3(new_n824), .ZN(new_n1100));
  AOI21_X1  g675(.A(G301), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  NAND4_X1  g676(.A1(new_n1085), .A2(new_n1092), .A3(new_n1095), .A4(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1051), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1066), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1104), .A2(new_n1055), .ZN(new_n1105));
  AOI22_X1  g680(.A1(new_n1103), .A2(new_n1073), .B1(new_n1105), .B2(new_n1064), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1084), .A2(new_n1102), .A3(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1049), .A2(new_n829), .ZN(new_n1108));
  INV_X1    g683(.A(G2067), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1062), .A2(new_n1109), .ZN(new_n1110));
  OR2_X1    g685(.A1(new_n597), .A2(KEYINPUT123), .ZN(new_n1111));
  NAND4_X1  g686(.A1(new_n1108), .A2(new_n1110), .A3(KEYINPUT60), .A4(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n597), .A2(KEYINPUT123), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1049), .A2(new_n829), .B1(new_n1062), .B2(new_n1109), .ZN(new_n1116));
  OR2_X1    g691(.A1(new_n1116), .A2(KEYINPUT60), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1116), .A2(KEYINPUT60), .A3(new_n1113), .A4(new_n1111), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1115), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT61), .ZN(new_n1120));
  XNOR2_X1  g695(.A(KEYINPUT56), .B(G2072), .ZN(new_n1121));
  AOI22_X1  g696(.A1(new_n1099), .A2(new_n1121), .B1(new_n1039), .B2(new_n795), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT57), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n554), .A2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1124), .A2(KEYINPUT121), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n1126));
  NOR3_X1   g701(.A1(new_n554), .A2(new_n1126), .A3(new_n1123), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n553), .A2(new_n548), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT120), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n553), .A2(KEYINPUT120), .A3(new_n548), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n1130), .A2(new_n547), .A3(new_n1131), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1125), .A2(new_n1127), .B1(new_n1132), .B2(KEYINPUT57), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n1120), .B1(new_n1122), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1039), .A2(new_n795), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1029), .A2(new_n1008), .A3(new_n1030), .A4(new_n1121), .ZN(new_n1136));
  AND4_X1   g711(.A1(new_n1120), .A2(new_n1135), .A3(new_n1133), .A4(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT58), .B(G1341), .Z(new_n1139));
  OAI21_X1  g714(.A(new_n1139), .B1(new_n1002), .B2(new_n1007), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  OAI211_X1 g717(.A(KEYINPUT122), .B(new_n1139), .C1(new_n1002), .C2(new_n1007), .ZN(new_n1143));
  OAI211_X1 g718(.A(new_n1142), .B(new_n1143), .C1(new_n1031), .C2(G1996), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1144), .A2(KEYINPUT59), .A3(new_n536), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT59), .B1(new_n1144), .B2(new_n536), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1119), .A2(new_n1138), .A3(new_n1147), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1122), .A2(new_n1133), .ZN(new_n1150));
  INV_X1    g725(.A(new_n1116), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1150), .A2(new_n598), .A3(new_n1151), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n1148), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1093), .B1(new_n1089), .B2(new_n1087), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1098), .A2(new_n1100), .ZN(new_n1155));
  XNOR2_X1  g730(.A(G171), .B(KEYINPUT54), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(G160), .A2(G40), .ZN(new_n1159));
  XNOR2_X1  g734(.A(new_n1159), .B(KEYINPUT124), .ZN(new_n1160));
  OR2_X1    g735(.A1(KEYINPUT125), .A2(G2078), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1097), .B1(KEYINPUT125), .B2(G2078), .ZN(new_n1162));
  NAND4_X1  g737(.A1(new_n1160), .A2(new_n1030), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1098), .B(new_n1156), .C1(new_n1163), .C2(new_n1004), .ZN(new_n1164));
  NAND4_X1  g739(.A1(new_n1085), .A2(new_n1154), .A3(new_n1158), .A4(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1027), .B1(new_n1107), .B2(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1021), .A2(new_n1023), .A3(new_n713), .A4(new_n710), .ZN(new_n1168));
  OR2_X1    g743(.A1(new_n842), .A2(G2067), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT126), .ZN(new_n1171));
  INV_X1    g746(.A(KEYINPUT126), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1168), .A2(new_n1172), .A3(new_n1169), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1171), .A2(new_n1014), .A3(new_n1173), .ZN(new_n1174));
  XOR2_X1   g749(.A(new_n1011), .B(KEYINPUT48), .Z(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1026), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1014), .B1(new_n767), .B2(new_n1016), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1014), .A2(KEYINPUT46), .A3(new_n1017), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT46), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1179), .B1(new_n1009), .B2(G1996), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1177), .A2(new_n1178), .A3(new_n1180), .ZN(new_n1181));
  XNOR2_X1  g756(.A(new_n1181), .B(KEYINPUT47), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1174), .A2(new_n1176), .A3(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1167), .A2(new_n1183), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g759(.A1(new_n661), .A2(G319), .A3(new_n677), .ZN(new_n1186));
  NAND2_X1  g760(.A1(new_n1186), .A2(KEYINPUT127), .ZN(new_n1187));
  INV_X1    g761(.A(KEYINPUT127), .ZN(new_n1188));
  NAND4_X1  g762(.A1(new_n661), .A2(new_n1188), .A3(G319), .A4(new_n677), .ZN(new_n1189));
  AOI21_X1  g763(.A(G229), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AND4_X1   g764(.A1(new_n912), .A2(new_n1190), .A3(new_n995), .A4(new_n988), .ZN(G308));
  NAND4_X1  g765(.A1(new_n912), .A2(new_n1190), .A3(new_n995), .A4(new_n988), .ZN(G225));
endmodule


