//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950;
  INV_X1    g000(.A(G902), .ZN(new_n187));
  INV_X1    g001(.A(G237), .ZN(new_n188));
  INV_X1    g002(.A(G953), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n188), .A2(new_n189), .A3(G214), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  NAND2_X1  g006(.A1(KEYINPUT18), .A2(G131), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n192), .B(new_n193), .ZN(new_n194));
  XNOR2_X1  g008(.A(G125), .B(G140), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  AND2_X1   g011(.A1(KEYINPUT79), .A2(G125), .ZN(new_n198));
  NOR2_X1   g012(.A1(KEYINPUT79), .A2(G125), .ZN(new_n199));
  OAI21_X1  g013(.A(G140), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  NOR2_X1   g014(.A1(G125), .A2(G140), .ZN(new_n201));
  INV_X1    g015(.A(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(new_n203), .B2(new_n196), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n194), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT66), .B(G131), .ZN(new_n206));
  XNOR2_X1  g020(.A(new_n192), .B(new_n206), .ZN(new_n207));
  OR2_X1    g021(.A1(new_n207), .A2(KEYINPUT17), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n192), .A2(KEYINPUT17), .A3(new_n206), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n211), .B1(new_n200), .B2(new_n202), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n198), .A2(new_n199), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n213), .A2(KEYINPUT16), .A3(G140), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n196), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT79), .B(G125), .ZN(new_n217));
  INV_X1    g031(.A(G140), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n211), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n201), .B1(new_n217), .B2(G140), .ZN(new_n220));
  OAI211_X1 g034(.A(G146), .B(new_n219), .C1(new_n220), .C2(new_n211), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n215), .A2(new_n216), .A3(new_n221), .ZN(new_n222));
  OAI211_X1 g036(.A(KEYINPUT80), .B(new_n196), .C1(new_n212), .C2(new_n214), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n210), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT92), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n208), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI211_X1 g040(.A(KEYINPUT92), .B(new_n210), .C1(new_n222), .C2(new_n223), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n205), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G113), .B(G122), .ZN(new_n229));
  INV_X1    g043(.A(G104), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n229), .B(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n228), .A2(new_n232), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n231), .B(new_n205), .C1(new_n226), .C2(new_n227), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n187), .B1(new_n233), .B2(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G475), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n203), .A2(KEYINPUT19), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n195), .A2(KEYINPUT19), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(KEYINPUT91), .B1(new_n240), .B2(G146), .ZN(new_n241));
  INV_X1    g055(.A(KEYINPUT91), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n242), .B(new_n196), .C1(new_n238), .C2(new_n239), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n241), .A2(new_n207), .A3(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n221), .B(KEYINPUT81), .ZN(new_n245));
  INV_X1    g059(.A(new_n245), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n205), .B1(new_n244), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n247), .A2(new_n232), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n234), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT93), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT20), .ZN(new_n252));
  NOR2_X1   g066(.A1(G475), .A2(G902), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n251), .A2(new_n252), .B1(new_n249), .B2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n249), .A2(KEYINPUT93), .A3(new_n252), .A4(new_n253), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n237), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT94), .ZN(new_n258));
  NAND2_X1  g072(.A1(G234), .A2(G237), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(G952), .A3(new_n189), .ZN(new_n260));
  XOR2_X1   g074(.A(new_n260), .B(KEYINPUT97), .Z(new_n261));
  AND3_X1   g075(.A1(new_n259), .A2(G902), .A3(G953), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT21), .B(G898), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n249), .A2(new_n253), .ZN(new_n267));
  AOI21_X1  g081(.A(KEYINPUT93), .B1(new_n234), .B2(new_n248), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n267), .B1(KEYINPUT20), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n255), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT94), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n237), .ZN(new_n272));
  XNOR2_X1  g086(.A(G116), .B(G122), .ZN(new_n273));
  XNOR2_X1  g087(.A(new_n273), .B(G107), .ZN(new_n274));
  XNOR2_X1  g088(.A(G128), .B(G143), .ZN(new_n275));
  INV_X1    g089(.A(G134), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OR2_X1    g091(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G128), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n279), .A2(KEYINPUT13), .A3(G143), .ZN(new_n280));
  AOI211_X1 g094(.A(new_n276), .B(new_n280), .C1(KEYINPUT13), .C2(new_n275), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n275), .A2(new_n276), .ZN(new_n282));
  OAI21_X1  g096(.A(KEYINPUT95), .B1(new_n277), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G107), .ZN(new_n284));
  INV_X1    g098(.A(G116), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n285), .A2(G122), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n286), .B2(KEYINPUT14), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT14), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n273), .A2(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n287), .A2(new_n289), .B1(new_n284), .B2(new_n273), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  NOR3_X1   g105(.A1(new_n277), .A2(new_n282), .A3(KEYINPUT95), .ZN(new_n292));
  OAI22_X1  g106(.A1(new_n278), .A2(new_n281), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(G217), .A3(new_n189), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n293), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT96), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n293), .A2(new_n296), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n293), .A2(KEYINPUT96), .A3(new_n296), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(G902), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n303), .B(new_n305), .ZN(new_n306));
  NAND4_X1  g120(.A1(new_n258), .A2(new_n266), .A3(new_n272), .A4(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G221), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n309), .B1(new_n295), .B2(new_n187), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G110), .B(G140), .ZN(new_n312));
  AND2_X1   g126(.A1(new_n189), .A2(G227), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n312), .B(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT10), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT1), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n196), .A2(G143), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n191), .A2(G146), .ZN(new_n318));
  AND4_X1   g132(.A1(new_n316), .A2(new_n317), .A3(new_n318), .A4(G128), .ZN(new_n319));
  OAI21_X1  g133(.A(KEYINPUT1), .B1(new_n191), .B2(G146), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n320), .A2(G128), .B1(new_n317), .B2(new_n318), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g136(.A(KEYINPUT3), .B1(new_n230), .B2(G107), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(new_n284), .A3(G104), .ZN(new_n325));
  INV_X1    g139(.A(G101), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n230), .A2(G107), .ZN(new_n327));
  NAND4_X1  g141(.A1(new_n323), .A2(new_n325), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n230), .A2(G107), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n284), .A2(G104), .ZN(new_n330));
  OAI21_X1  g144(.A(G101), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n315), .B1(new_n322), .B2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n320), .A2(G128), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n317), .A2(new_n318), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G143), .B(G146), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G128), .A3(new_n320), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n339), .A2(KEYINPUT10), .A3(new_n331), .A4(new_n328), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n333), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n323), .A2(new_n325), .A3(new_n327), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(G101), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n343), .A2(KEYINPUT4), .A3(new_n328), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n335), .A2(KEYINPUT65), .A3(KEYINPUT0), .A4(G128), .ZN(new_n345));
  NAND2_X1  g159(.A1(KEYINPUT0), .A2(G128), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT65), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n346), .B1(new_n337), .B2(new_n347), .ZN(new_n348));
  OR3_X1    g162(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n335), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n345), .A2(new_n348), .A3(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT4), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n342), .A2(new_n353), .A3(G101), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT86), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT86), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n344), .A2(new_n352), .A3(new_n357), .A4(new_n354), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n341), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT69), .ZN(new_n360));
  INV_X1    g174(.A(G131), .ZN(new_n361));
  INV_X1    g175(.A(G137), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT11), .B1(new_n362), .B2(G134), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(G134), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(KEYINPUT11), .A3(G134), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n361), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT11), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n368), .B1(new_n276), .B2(G137), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n276), .A2(G137), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n366), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n371), .A2(new_n206), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n360), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n206), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(new_n365), .A3(new_n366), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(G131), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(KEYINPUT69), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  AND2_X1   g192(.A1(new_n359), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n359), .A2(new_n378), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n314), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n314), .B1(new_n359), .B2(new_n378), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n322), .B(new_n332), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n375), .A2(new_n376), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n383), .A2(KEYINPUT12), .A3(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(new_n339), .B(new_n332), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n378), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n385), .B1(new_n387), .B2(KEYINPUT12), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n388), .ZN(new_n389));
  AOI211_X1 g203(.A(G469), .B(G902), .C1(new_n381), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n359), .A2(new_n378), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n388), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(new_n314), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n382), .B1(new_n378), .B2(new_n359), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(new_n394), .A3(G469), .ZN(new_n395));
  INV_X1    g209(.A(G469), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n396), .A2(new_n187), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n311), .B1(new_n390), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n400), .A2(KEYINPUT87), .ZN(new_n401));
  OAI21_X1  g215(.A(G214), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n352), .A2(new_n217), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n404), .B1(new_n217), .B2(new_n322), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n189), .A2(G224), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n405), .B1(KEYINPUT7), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G119), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G116), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n285), .A2(G119), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n409), .A2(new_n410), .A3(KEYINPUT5), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n411), .B(G113), .C1(KEYINPUT5), .C2(new_n409), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n409), .A2(new_n410), .ZN(new_n413));
  XNOR2_X1  g227(.A(KEYINPUT2), .B(G113), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n412), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n415), .B(new_n332), .ZN(new_n416));
  XNOR2_X1  g230(.A(G110), .B(G122), .ZN(new_n417));
  XNOR2_X1  g231(.A(new_n417), .B(KEYINPUT8), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n407), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n406), .ZN(new_n420));
  OR2_X1    g234(.A1(new_n420), .A2(KEYINPUT89), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT7), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n422), .B1(new_n420), .B2(KEYINPUT89), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n405), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT90), .ZN(new_n425));
  OR2_X1    g239(.A1(new_n415), .A2(new_n332), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n413), .A2(KEYINPUT68), .ZN(new_n427));
  INV_X1    g241(.A(new_n414), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT68), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n344), .A3(new_n354), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n417), .A3(new_n432), .ZN(new_n433));
  OR2_X1    g247(.A1(new_n424), .A2(KEYINPUT90), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n419), .A2(new_n425), .A3(new_n433), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n426), .A2(new_n432), .ZN(new_n436));
  INV_X1    g250(.A(new_n417), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n438), .A2(KEYINPUT6), .A3(new_n433), .ZN(new_n439));
  XNOR2_X1  g253(.A(new_n406), .B(KEYINPUT88), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n405), .B(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT6), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n436), .A2(new_n442), .A3(new_n437), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n435), .A2(new_n187), .A3(new_n444), .ZN(new_n445));
  OAI21_X1  g259(.A(G210), .B1(G237), .B2(G902), .ZN(new_n446));
  INV_X1    g260(.A(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n435), .A2(new_n444), .A3(new_n187), .A4(new_n446), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n403), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n381), .A2(new_n389), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n451), .A2(new_n396), .A3(new_n187), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n398), .A3(new_n395), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT87), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n311), .ZN(new_n455));
  AND3_X1   g269(.A1(new_n401), .A2(new_n450), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n308), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(G472), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT73), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT71), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n413), .A2(new_n414), .A3(KEYINPUT68), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n414), .B1(KEYINPUT68), .B2(new_n413), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n429), .A2(KEYINPUT71), .A3(new_n430), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n362), .A2(G134), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n465), .A2(new_n370), .A3(KEYINPUT67), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT67), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n361), .B1(new_n364), .B2(new_n467), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n336), .A2(new_n338), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  AOI22_X1  g283(.A1(new_n463), .A2(new_n464), .B1(new_n469), .B2(new_n375), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n373), .A2(new_n352), .A3(new_n377), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT28), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n459), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI211_X1 g288(.A(KEYINPUT73), .B(KEYINPUT28), .C1(new_n470), .C2(new_n471), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  XOR2_X1   g290(.A(KEYINPUT72), .B(KEYINPUT27), .Z(new_n477));
  NAND3_X1  g291(.A1(new_n188), .A2(new_n189), .A3(G210), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XNOR2_X1  g293(.A(KEYINPUT26), .B(G101), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT29), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n471), .A2(KEYINPUT70), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n469), .A2(new_n375), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT70), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n373), .A2(new_n486), .A3(new_n377), .A4(new_n352), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n463), .A2(new_n464), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n484), .A2(new_n470), .A3(new_n487), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n476), .B(new_n483), .C1(new_n492), .C2(new_n473), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n493), .A2(KEYINPUT76), .A3(new_n187), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT76), .B1(new_n493), .B2(new_n187), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n384), .A2(new_n352), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n485), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(new_n431), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n491), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n500), .A2(KEYINPUT28), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n476), .ZN(new_n502));
  INV_X1    g316(.A(new_n481), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(KEYINPUT29), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT75), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n498), .A2(KEYINPUT30), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n507), .B1(new_n488), .B2(KEYINPUT30), .ZN(new_n508));
  INV_X1    g322(.A(new_n431), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n491), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n506), .B1(new_n511), .B2(new_n481), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n510), .A2(KEYINPUT75), .A3(new_n503), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n505), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n458), .B1(new_n496), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(G472), .A2(G902), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT74), .ZN(new_n519));
  OAI211_X1 g333(.A(new_n481), .B(new_n491), .C1(new_n508), .C2(new_n509), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT31), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n502), .A2(new_n503), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n520), .A2(KEYINPUT31), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n520), .A2(KEYINPUT31), .B1(new_n502), .B2(new_n503), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n488), .A2(KEYINPUT30), .ZN(new_n527));
  INV_X1    g341(.A(new_n507), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n431), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT31), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n481), .A4(new_n491), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n526), .A2(KEYINPUT74), .A3(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n518), .B1(new_n525), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AND4_X1   g350(.A1(KEYINPUT74), .A2(new_n532), .A3(new_n521), .A4(new_n522), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT74), .B1(new_n526), .B2(new_n532), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n535), .B(new_n517), .C1(new_n537), .C2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n516), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT85), .ZN(new_n542));
  XOR2_X1   g356(.A(G119), .B(G128), .Z(new_n543));
  XNOR2_X1  g357(.A(new_n543), .B(KEYINPUT77), .ZN(new_n544));
  XOR2_X1   g358(.A(KEYINPUT24), .B(G110), .Z(new_n545));
  INV_X1    g359(.A(KEYINPUT78), .ZN(new_n546));
  OAI211_X1 g360(.A(G119), .B(new_n279), .C1(new_n546), .C2(KEYINPUT23), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT23), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n548), .B1(new_n408), .B2(G128), .ZN(new_n549));
  OAI21_X1  g363(.A(KEYINPUT78), .B1(new_n408), .B2(G128), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI22_X1  g365(.A1(new_n544), .A2(new_n545), .B1(G110), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n245), .A2(new_n197), .A3(new_n552), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n544), .A2(new_n545), .B1(G110), .B2(new_n551), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n222), .A2(new_n554), .A3(new_n223), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  XNOR2_X1  g370(.A(KEYINPUT22), .B(G137), .ZN(new_n557));
  INV_X1    g371(.A(G234), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n309), .A2(new_n558), .A3(G953), .ZN(new_n559));
  XOR2_X1   g373(.A(new_n557), .B(new_n559), .Z(new_n560));
  INV_X1    g374(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n556), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n553), .A2(new_n555), .A3(new_n560), .ZN(new_n563));
  OAI21_X1  g377(.A(G217), .B1(new_n558), .B2(G902), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(new_n187), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n565), .B(KEYINPUT83), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n562), .A2(new_n563), .A3(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT84), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n568), .B(new_n569), .ZN(new_n570));
  AND3_X1   g384(.A1(new_n553), .A2(new_n555), .A3(new_n560), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n560), .B1(new_n553), .B2(new_n555), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(KEYINPUT25), .B1(new_n573), .B2(new_n187), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n564), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT25), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n562), .A2(new_n563), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n577), .B1(new_n578), .B2(G902), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n573), .A2(KEYINPUT25), .A3(new_n187), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT82), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n570), .B1(new_n576), .B2(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n541), .A2(new_n542), .A3(new_n582), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n517), .B1(new_n537), .B2(new_n538), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT32), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n515), .B1(new_n585), .B2(new_n539), .ZN(new_n586));
  INV_X1    g400(.A(new_n582), .ZN(new_n587));
  OAI21_X1  g401(.A(KEYINPUT85), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n457), .B1(new_n583), .B2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(new_n326), .ZN(G3));
  OAI21_X1  g404(.A(new_n187), .B1(new_n537), .B2(new_n538), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n584), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n401), .A2(new_n455), .A3(new_n582), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT98), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT99), .B(G478), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n303), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n302), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT33), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n293), .B2(new_n296), .ZN(new_n601));
  AOI22_X1  g415(.A1(new_n599), .A2(new_n600), .B1(new_n297), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n304), .A2(G902), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n450), .A2(new_n266), .ZN(new_n605));
  AOI211_X1 g419(.A(new_n604), .B(new_n605), .C1(new_n258), .C2(new_n272), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n596), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(KEYINPUT100), .ZN(new_n608));
  XOR2_X1   g422(.A(KEYINPUT34), .B(G104), .Z(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G6));
  INV_X1    g424(.A(new_n605), .ZN(new_n611));
  INV_X1    g425(.A(new_n306), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n267), .B(KEYINPUT20), .ZN(new_n613));
  AND4_X1   g427(.A1(new_n237), .A2(new_n611), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n596), .A2(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT35), .B(G107), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G9));
  AOI21_X1  g431(.A(G902), .B1(new_n525), .B2(new_n533), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n618), .A2(new_n458), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n534), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n576), .A2(new_n581), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n561), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n556), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n567), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n308), .A2(new_n620), .A3(new_n456), .A4(new_n625), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT37), .B(G110), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G12));
  INV_X1    g442(.A(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n585), .A2(new_n539), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n629), .B1(new_n630), .B2(new_n516), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n262), .A2(new_n632), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n261), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  AND4_X1   g449(.A1(new_n237), .A2(new_n612), .A3(new_n613), .A4(new_n635), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n636), .A2(new_n456), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  NAND2_X1  g453(.A1(new_n448), .A2(new_n449), .ZN(new_n640));
  XOR2_X1   g454(.A(new_n640), .B(KEYINPUT38), .Z(new_n641));
  AND2_X1   g455(.A1(new_n401), .A2(new_n455), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n634), .B(KEYINPUT39), .Z(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT103), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT103), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n645), .A2(KEYINPUT40), .A3(new_n646), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n641), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g465(.A(G902), .B1(new_n492), .B2(new_n503), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n510), .A2(new_n481), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n630), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT101), .Z(new_n657));
  INV_X1    g471(.A(new_n272), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n271), .B1(new_n270), .B2(new_n237), .ZN(new_n659));
  OAI21_X1  g473(.A(new_n612), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n660), .A2(new_n403), .A3(new_n625), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(KEYINPUT102), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n651), .A2(new_n657), .A3(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(G143), .ZN(G45));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n541), .A2(new_n625), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n258), .A2(new_n272), .ZN(new_n667));
  INV_X1    g481(.A(new_n604), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n456), .A2(new_n667), .A3(new_n668), .A4(new_n635), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n665), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n669), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n671), .A2(new_n631), .A3(KEYINPUT104), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n670), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  NAND2_X1  g488(.A1(new_n451), .A2(new_n187), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n675), .A2(KEYINPUT105), .A3(G469), .ZN(new_n676));
  NAND2_X1  g490(.A1(KEYINPUT105), .A2(G469), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n451), .A2(new_n187), .A3(new_n677), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(new_n311), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n541), .A2(new_n606), .A3(new_n582), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(KEYINPUT41), .B(G113), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n541), .A2(new_n614), .A3(new_n582), .A4(new_n681), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n450), .A3(new_n311), .ZN(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n541), .A2(new_n308), .A3(new_n625), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G119), .ZN(G21));
  NAND2_X1  g504(.A1(new_n660), .A2(KEYINPUT108), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT108), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n667), .A2(new_n692), .A3(new_n612), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n680), .A2(new_n605), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n691), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n476), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n473), .B1(new_n490), .B2(new_n491), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n503), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT106), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n521), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(new_n532), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n700), .B1(new_n521), .B2(new_n699), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n517), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI211_X1 g518(.A(new_n704), .B(new_n582), .C1(new_n618), .C2(new_n458), .ZN(new_n705));
  XOR2_X1   g519(.A(new_n705), .B(KEYINPUT107), .Z(new_n706));
  NAND2_X1  g520(.A1(new_n696), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G122), .ZN(G24));
  OAI211_X1 g522(.A(new_n704), .B(new_n625), .C1(new_n618), .C2(new_n458), .ZN(new_n709));
  INV_X1    g523(.A(KEYINPUT109), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n592), .A2(KEYINPUT109), .A3(new_n625), .A4(new_n704), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND4_X1   g527(.A1(new_n667), .A2(new_n688), .A3(new_n668), .A4(new_n635), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  AOI211_X1 g530(.A(new_n604), .B(new_n634), .C1(new_n258), .C2(new_n272), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n640), .A2(new_n403), .ZN(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n400), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n541), .A2(new_n717), .A3(new_n582), .A4(new_n720), .ZN(new_n721));
  NOR2_X1   g535(.A1(KEYINPUT110), .A2(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n586), .A2(new_n587), .ZN(new_n724));
  INV_X1    g538(.A(new_n722), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n717), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G131), .ZN(G33));
  NAND4_X1  g542(.A1(new_n541), .A2(new_n582), .A3(new_n636), .A4(new_n720), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT111), .B(G134), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G36));
  NAND2_X1  g545(.A1(new_n593), .A2(new_n625), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(KEYINPUT115), .ZN(new_n733));
  INV_X1    g547(.A(new_n667), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n668), .ZN(new_n735));
  NAND2_X1  g549(.A1(KEYINPUT114), .A2(KEYINPUT43), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(KEYINPUT114), .B(KEYINPUT43), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n668), .A3(new_n738), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n733), .A2(new_n740), .ZN(new_n741));
  OR2_X1    g555(.A1(new_n741), .A2(KEYINPUT44), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n741), .A2(KEYINPUT44), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n393), .A2(new_n394), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT45), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(KEYINPUT112), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n396), .B1(new_n744), .B2(new_n745), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g563(.A(KEYINPUT113), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n747), .A2(KEYINPUT113), .A3(new_n748), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n397), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AND2_X1   g567(.A1(new_n753), .A2(KEYINPUT46), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n452), .B1(new_n753), .B2(KEYINPUT46), .ZN(new_n755));
  OAI211_X1 g569(.A(new_n311), .B(new_n643), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n719), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n742), .A2(new_n743), .A3(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  NAND4_X1  g573(.A1(new_n717), .A2(new_n586), .A3(new_n587), .A4(new_n718), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n311), .B1(new_n754), .B2(new_n755), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT47), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g577(.A(KEYINPUT47), .B(new_n311), .C1(new_n754), .C2(new_n755), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n760), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(new_n218), .ZN(G42));
  INV_X1    g580(.A(new_n679), .ZN(new_n767));
  OR2_X1    g581(.A1(new_n767), .A2(KEYINPUT49), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n587), .A2(new_n403), .A3(new_n310), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(KEYINPUT49), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n768), .A2(new_n769), .A3(new_n641), .A4(new_n770), .ZN(new_n771));
  OR3_X1    g585(.A1(new_n657), .A2(new_n735), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n261), .B1(new_n737), .B2(new_n739), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n773), .A2(new_n706), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n641), .A2(new_n403), .A3(new_n681), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT50), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n774), .A2(KEYINPUT50), .A3(new_n775), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n681), .A2(new_n718), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(KEYINPUT117), .ZN(new_n782));
  INV_X1    g596(.A(new_n261), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n783), .A3(new_n582), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT118), .ZN(new_n785));
  OR3_X1    g599(.A1(new_n657), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n785), .B1(new_n657), .B2(new_n784), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n786), .A2(new_n734), .A3(new_n604), .A4(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n773), .A2(new_n713), .A3(new_n782), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n780), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n763), .B(new_n764), .C1(new_n311), .C2(new_n767), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n791), .A2(new_n718), .A3(new_n774), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT116), .ZN(new_n793));
  OAI211_X1 g607(.A(new_n790), .B(new_n792), .C1(new_n793), .C2(KEYINPUT51), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n780), .A2(new_n788), .A3(new_n792), .A4(new_n789), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n780), .A2(new_n788), .A3(new_n793), .A4(new_n789), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n786), .A2(new_n667), .A3(new_n668), .A4(new_n787), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n773), .A2(new_n724), .A3(new_n782), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT48), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n189), .A2(G952), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n774), .B2(new_n688), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT119), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT119), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n794), .A2(new_n798), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g623(.A1(new_n713), .A2(new_n714), .B1(new_n631), .B2(new_n637), .ZN(new_n810));
  OR3_X1    g624(.A1(new_n625), .A2(new_n400), .A3(new_n634), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n811), .B1(new_n630), .B2(new_n655), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n812), .A2(new_n450), .A3(new_n691), .A4(new_n693), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT104), .B1(new_n671), .B2(new_n631), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n669), .A2(new_n586), .A3(new_n665), .A4(new_n629), .ZN(new_n815));
  OAI211_X1 g629(.A(new_n810), .B(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(KEYINPUT52), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT52), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n673), .A2(new_n818), .A3(new_n810), .A4(new_n813), .ZN(new_n819));
  XNOR2_X1  g633(.A(new_n705), .B(KEYINPUT107), .ZN(new_n820));
  OAI211_X1 g634(.A(new_n682), .B(new_n685), .C1(new_n820), .C2(new_n695), .ZN(new_n821));
  NOR4_X1   g635(.A1(new_n619), .A2(new_n594), .A3(new_n534), .A4(new_n605), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n658), .A2(new_n659), .A3(new_n612), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n668), .B1(new_n258), .B2(new_n272), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n826), .A2(new_n626), .A3(new_n689), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n821), .A2(new_n827), .A3(new_n589), .ZN(new_n828));
  AND4_X1   g642(.A1(new_n667), .A2(new_n720), .A3(new_n668), .A4(new_n635), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n713), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n613), .A2(new_n635), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n306), .A2(new_n237), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n719), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n541), .A2(new_n833), .A3(new_n642), .A4(new_n625), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n830), .A2(new_n729), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n835), .B1(new_n726), .B2(new_n723), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n817), .A2(new_n819), .A3(new_n828), .A4(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n826), .A2(new_n626), .A3(new_n689), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n583), .A2(new_n588), .ZN(new_n841));
  INV_X1    g655(.A(new_n457), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n682), .A2(new_n685), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n840), .A2(new_n843), .A3(new_n707), .A4(new_n844), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n834), .A2(new_n729), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n727), .A2(new_n830), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n848), .A2(KEYINPUT53), .A3(new_n819), .A4(new_n817), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n839), .A2(new_n849), .A3(KEYINPUT54), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT54), .B1(new_n839), .B2(new_n849), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n809), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(G952), .A2(G953), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n772), .B1(new_n854), .B2(new_n855), .ZN(G75));
  AOI21_X1  g670(.A(new_n187), .B1(new_n839), .B2(new_n849), .ZN(new_n857));
  AOI21_X1  g671(.A(KEYINPUT56), .B1(new_n857), .B2(G210), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n439), .A2(new_n443), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n859), .B(new_n441), .ZN(new_n860));
  XNOR2_X1  g674(.A(new_n860), .B(KEYINPUT55), .ZN(new_n861));
  NOR2_X1   g675(.A1(KEYINPUT120), .A2(KEYINPUT56), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n858), .A2(new_n863), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n189), .A2(G952), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n864), .A2(new_n865), .A3(new_n866), .ZN(G51));
  NAND2_X1  g681(.A1(new_n839), .A2(new_n849), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT54), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n397), .B(KEYINPUT57), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n850), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT121), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n870), .A2(KEYINPUT121), .A3(new_n850), .A4(new_n871), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n874), .A2(new_n451), .A3(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n857), .A2(new_n751), .A3(new_n752), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n866), .B1(new_n876), .B2(new_n877), .ZN(G54));
  NAND3_X1  g692(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .ZN(new_n879));
  INV_X1    g693(.A(new_n249), .ZN(new_n880));
  OR3_X1    g694(.A1(new_n879), .A2(KEYINPUT122), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g695(.A(KEYINPUT122), .B1(new_n879), .B2(new_n880), .ZN(new_n882));
  AOI21_X1  g696(.A(new_n866), .B1(new_n879), .B2(new_n880), .ZN(new_n883));
  AND3_X1   g697(.A1(new_n881), .A2(new_n882), .A3(new_n883), .ZN(G60));
  INV_X1    g698(.A(new_n866), .ZN(new_n885));
  NAND2_X1  g699(.A1(G478), .A2(G902), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT59), .Z(new_n887));
  NOR3_X1   g701(.A1(new_n851), .A2(new_n852), .A3(new_n887), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n885), .B1(new_n888), .B2(new_n602), .ZN(new_n889));
  INV_X1    g703(.A(new_n887), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n853), .A2(new_n602), .A3(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT123), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n888), .A2(new_n893), .A3(new_n602), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n889), .B1(new_n892), .B2(new_n894), .ZN(G63));
  NAND2_X1  g709(.A1(G217), .A2(G902), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT60), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n868), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n623), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n885), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  XNOR2_X1  g715(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n902));
  INV_X1    g716(.A(new_n898), .ZN(new_n903));
  XNOR2_X1  g717(.A(new_n578), .B(KEYINPUT124), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n901), .B(new_n902), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(new_n902), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n903), .A2(new_n904), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n906), .B1(new_n907), .B2(new_n900), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n905), .A2(new_n908), .ZN(G66));
  INV_X1    g723(.A(new_n263), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n189), .B1(new_n910), .B2(G224), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n911), .B1(new_n845), .B2(new_n189), .ZN(new_n912));
  INV_X1    g726(.A(G898), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n859), .B1(new_n913), .B2(G953), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n912), .B(new_n914), .ZN(G69));
  XNOR2_X1  g729(.A(new_n508), .B(new_n240), .ZN(new_n916));
  INV_X1    g730(.A(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n663), .A2(new_n673), .A3(new_n810), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NOR4_X1   g734(.A1(new_n647), .A2(new_n823), .A3(new_n719), .A4(new_n824), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n765), .B1(new_n841), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n663), .A2(new_n673), .A3(new_n810), .A4(new_n923), .ZN(new_n924));
  AND4_X1   g738(.A1(new_n758), .A2(new_n920), .A3(new_n922), .A4(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n917), .B1(new_n925), .B2(G953), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n189), .B1(G227), .B2(G900), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT127), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n691), .A2(new_n450), .A3(new_n693), .ZN(new_n931));
  NOR4_X1   g745(.A1(new_n756), .A2(new_n586), .A3(new_n587), .A4(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n729), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n765), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n727), .A2(new_n673), .A3(new_n810), .ZN(new_n935));
  NAND4_X1  g749(.A1(new_n934), .A2(new_n758), .A3(new_n189), .A4(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n917), .B1(G900), .B2(G953), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n936), .A2(new_n937), .B1(new_n928), .B2(new_n927), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n926), .A2(new_n930), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n930), .B1(new_n926), .B2(new_n938), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n939), .A2(new_n940), .ZN(G72));
  NAND2_X1  g755(.A1(new_n925), .A2(new_n828), .ZN(new_n942));
  NAND2_X1  g756(.A1(G472), .A2(G902), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n943), .B(KEYINPUT63), .Z(new_n944));
  AOI21_X1  g758(.A(new_n653), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n934), .A2(new_n758), .A3(new_n935), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n944), .B1(new_n946), .B2(new_n845), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n947), .A2(new_n503), .A3(new_n511), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n512), .A2(new_n513), .A3(new_n520), .ZN(new_n949));
  AND3_X1   g763(.A1(new_n868), .A2(new_n944), .A3(new_n949), .ZN(new_n950));
  NOR4_X1   g764(.A1(new_n945), .A2(new_n948), .A3(new_n866), .A4(new_n950), .ZN(G57));
endmodule


