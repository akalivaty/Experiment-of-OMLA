

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753;

  XNOR2_X1 U365 ( .A(n560), .B(n559), .ZN(n589) );
  AND2_X1 U366 ( .A1(n393), .A2(n391), .ZN(n390) );
  AND2_X1 U367 ( .A1(n633), .A2(n634), .ZN(n516) );
  XNOR2_X1 U368 ( .A(n596), .B(KEYINPUT38), .ZN(n687) );
  NAND2_X1 U369 ( .A1(n582), .A2(n687), .ZN(n560) );
  INV_X1 U370 ( .A(G953), .ZN(n746) );
  AND2_X2 U371 ( .A1(n384), .A2(n597), .ZN(n744) );
  NOR2_X1 U372 ( .A1(n751), .A2(n753), .ZN(n561) );
  XNOR2_X1 U373 ( .A(n367), .B(n428), .ZN(n464) );
  XNOR2_X2 U374 ( .A(n483), .B(KEYINPUT4), .ZN(n735) );
  OR2_X1 U375 ( .A1(n640), .A2(G902), .ZN(n465) );
  NAND2_X1 U376 ( .A1(n377), .A2(n380), .ZN(n751) );
  XNOR2_X1 U377 ( .A(n363), .B(n548), .ZN(n709) );
  XNOR2_X1 U378 ( .A(n457), .B(n456), .ZN(n695) );
  OR2_X1 U379 ( .A1(n653), .A2(G902), .ZN(n434) );
  XNOR2_X1 U380 ( .A(n399), .B(G146), .ZN(n442) );
  BUF_X1 U381 ( .A(n471), .Z(n343) );
  XNOR2_X2 U382 ( .A(n386), .B(n385), .ZN(n517) );
  NOR2_X2 U383 ( .A1(n558), .A2(n557), .ZN(n582) );
  XOR2_X1 U384 ( .A(KEYINPUT8), .B(KEYINPUT68), .Z(n437) );
  XOR2_X1 U385 ( .A(KEYINPUT70), .B(G131), .Z(n427) );
  XNOR2_X1 U386 ( .A(n547), .B(KEYINPUT105), .ZN(n684) );
  INV_X1 U387 ( .A(n670), .ZN(n372) );
  OR2_X1 U388 ( .A1(n686), .A2(n392), .ZN(n391) );
  NAND2_X1 U389 ( .A1(n389), .A2(n388), .ZN(n387) );
  AND2_X1 U390 ( .A1(n686), .A2(n392), .ZN(n388) );
  XNOR2_X1 U391 ( .A(n702), .B(n374), .ZN(n466) );
  INV_X1 U392 ( .A(KEYINPUT6), .ZN(n374) );
  XOR2_X1 U393 ( .A(G119), .B(G128), .Z(n394) );
  NAND2_X1 U394 ( .A1(n357), .A2(n356), .ZN(n563) );
  NAND2_X1 U395 ( .A1(n544), .A2(KEYINPUT28), .ZN(n356) );
  AND2_X1 U396 ( .A1(n360), .A2(n358), .ZN(n357) );
  AND2_X1 U397 ( .A1(n359), .A2(n546), .ZN(n358) );
  INV_X1 U398 ( .A(KEYINPUT40), .ZN(n383) );
  NAND2_X1 U399 ( .A1(n670), .A2(n383), .ZN(n381) );
  XNOR2_X1 U400 ( .A(n421), .B(n420), .ZN(n422) );
  INV_X1 U401 ( .A(KEYINPUT81), .ZN(n368) );
  INV_X1 U402 ( .A(G128), .ZN(n397) );
  INV_X1 U403 ( .A(G125), .ZN(n399) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n384) );
  INV_X1 U405 ( .A(KEYINPUT48), .ZN(n353) );
  NAND2_X1 U406 ( .A1(n588), .A2(n395), .ZN(n354) );
  NAND2_X1 U407 ( .A1(n566), .A2(KEYINPUT28), .ZN(n359) );
  NAND2_X1 U408 ( .A1(n362), .A2(n361), .ZN(n360) );
  NOR2_X1 U409 ( .A1(n566), .A2(KEYINPUT28), .ZN(n361) );
  XNOR2_X1 U410 ( .A(n545), .B(n435), .ZN(n508) );
  XNOR2_X1 U411 ( .A(G116), .B(G113), .ZN(n404) );
  XOR2_X1 U412 ( .A(G119), .B(KEYINPUT3), .Z(n405) );
  XNOR2_X1 U413 ( .A(G110), .B(G107), .ZN(n406) );
  BUF_X1 U414 ( .A(n682), .Z(n693) );
  NAND2_X1 U415 ( .A1(n684), .A2(n685), .ZN(n363) );
  AND2_X1 U416 ( .A1(n466), .A2(n372), .ZN(n570) );
  NOR2_X1 U417 ( .A1(n563), .A2(n345), .ZN(n575) );
  XNOR2_X1 U418 ( .A(n702), .B(n512), .ZN(n554) );
  BUF_X1 U419 ( .A(n702), .Z(n355) );
  BUF_X1 U420 ( .A(n508), .Z(n592) );
  INV_X1 U421 ( .A(n466), .ZN(n373) );
  INV_X1 U422 ( .A(KEYINPUT22), .ZN(n376) );
  XNOR2_X1 U423 ( .A(n448), .B(n447), .ZN(n645) );
  BUF_X1 U424 ( .A(n638), .Z(n650) );
  NAND2_X1 U425 ( .A1(n379), .A2(n378), .ZN(n377) );
  AND2_X1 U426 ( .A1(n382), .A2(n381), .ZN(n380) );
  NOR2_X1 U427 ( .A1(n670), .A2(n383), .ZN(n378) );
  INV_X1 U428 ( .A(KEYINPUT35), .ZN(n385) );
  AND2_X1 U429 ( .A1(n677), .A2(G478), .ZN(n344) );
  AND2_X1 U430 ( .A1(n390), .A2(n387), .ZN(n345) );
  AND2_X1 U431 ( .A1(n597), .A2(KEYINPUT2), .ZN(n346) );
  NOR2_X1 U432 ( .A1(n550), .A2(n355), .ZN(n347) );
  AND2_X1 U433 ( .A1(n531), .A2(n373), .ZN(n348) );
  AND2_X1 U434 ( .A1(n513), .A2(n554), .ZN(n349) );
  AND2_X1 U435 ( .A1(n510), .A2(n373), .ZN(n350) );
  AND2_X1 U436 ( .A1(n604), .A2(n744), .ZN(n351) );
  NAND2_X1 U437 ( .A1(n370), .A2(n744), .ZN(n369) );
  XNOR2_X1 U438 ( .A(n371), .B(n537), .ZN(n370) );
  NAND2_X1 U439 ( .A1(n390), .A2(n387), .ZN(n562) );
  XNOR2_X1 U440 ( .A(n736), .B(n396), .ZN(n447) );
  XNOR2_X1 U441 ( .A(n369), .B(n368), .ZN(n601) );
  XNOR2_X1 U442 ( .A(n352), .B(n472), .ZN(n365) );
  NAND2_X1 U443 ( .A1(n471), .A2(n366), .ZN(n352) );
  XNOR2_X1 U444 ( .A(n521), .B(KEYINPUT88), .ZN(n471) );
  BUF_X2 U445 ( .A(n572), .Z(n596) );
  INV_X1 U446 ( .A(n544), .ZN(n362) );
  NOR2_X1 U447 ( .A1(n709), .A2(n563), .ZN(n549) );
  OR2_X2 U448 ( .A1(n615), .A2(n536), .ZN(n364) );
  XNOR2_X2 U449 ( .A(n364), .B(n412), .ZN(n572) );
  NAND2_X1 U450 ( .A1(n365), .A2(n584), .ZN(n386) );
  INV_X1 U451 ( .A(n682), .ZN(n366) );
  XNOR2_X1 U452 ( .A(n367), .B(n403), .ZN(n409) );
  XNOR2_X2 U453 ( .A(n735), .B(G101), .ZN(n367) );
  NAND2_X1 U454 ( .A1(n603), .A2(n536), .ZN(n371) );
  AND2_X2 U455 ( .A1(n606), .A2(n677), .ZN(n638) );
  AND2_X1 U456 ( .A1(n606), .A2(n344), .ZN(n610) );
  NAND2_X1 U457 ( .A1(n375), .A2(n349), .ZN(n515) );
  NAND2_X1 U458 ( .A1(n375), .A2(n350), .ZN(n511) );
  NAND2_X1 U459 ( .A1(n375), .A2(n348), .ZN(n632) );
  XNOR2_X2 U460 ( .A(n507), .B(n376), .ZN(n375) );
  XNOR2_X2 U461 ( .A(n398), .B(n397), .ZN(n483) );
  NAND2_X1 U462 ( .A1(n589), .A2(n383), .ZN(n382) );
  INV_X1 U463 ( .A(n589), .ZN(n379) );
  NAND2_X1 U464 ( .A1(n384), .A2(n346), .ZN(n602) );
  INV_X1 U465 ( .A(n517), .ZN(n636) );
  NAND2_X1 U466 ( .A1(n343), .A2(n347), .ZN(n520) );
  INV_X1 U467 ( .A(n572), .ZN(n389) );
  INV_X1 U468 ( .A(n414), .ZN(n392) );
  NAND2_X1 U469 ( .A1(n572), .A2(n414), .ZN(n393) );
  NAND2_X1 U470 ( .A1(n562), .A2(n422), .ZN(n425) );
  NOR2_X1 U471 ( .A1(n587), .A2(n586), .ZN(n395) );
  XOR2_X1 U472 ( .A(n446), .B(n445), .Z(n396) );
  INV_X1 U473 ( .A(n667), .ZN(n586) );
  INV_X1 U474 ( .A(KEYINPUT39), .ZN(n559) );
  INV_X1 U475 ( .A(KEYINPUT120), .ZN(n613) );
  XNOR2_X2 U476 ( .A(G143), .B(KEYINPUT64), .ZN(n398) );
  XNOR2_X1 U477 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n401) );
  NAND2_X1 U478 ( .A1(n746), .A2(G224), .ZN(n400) );
  XNOR2_X1 U479 ( .A(n401), .B(n400), .ZN(n402) );
  XNOR2_X1 U480 ( .A(n442), .B(n402), .ZN(n403) );
  XNOR2_X1 U481 ( .A(n405), .B(n404), .ZN(n462) );
  XNOR2_X1 U482 ( .A(n406), .B(G104), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n462), .B(n429), .ZN(n408) );
  XOR2_X1 U484 ( .A(KEYINPUT16), .B(G122), .Z(n407) );
  XNOR2_X1 U485 ( .A(n408), .B(n407), .ZN(n728) );
  XNOR2_X1 U486 ( .A(n409), .B(n728), .ZN(n615) );
  XNOR2_X1 U487 ( .A(G902), .B(KEYINPUT15), .ZN(n599) );
  INV_X1 U488 ( .A(n599), .ZN(n536) );
  INV_X1 U489 ( .A(G902), .ZN(n500) );
  INV_X1 U490 ( .A(G237), .ZN(n410) );
  NAND2_X1 U491 ( .A1(n500), .A2(n410), .ZN(n413) );
  NAND2_X1 U492 ( .A1(n413), .A2(G210), .ZN(n411) );
  XNOR2_X1 U493 ( .A(n411), .B(KEYINPUT86), .ZN(n412) );
  NAND2_X1 U494 ( .A1(n413), .A2(G214), .ZN(n686) );
  XNOR2_X1 U495 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n414) );
  XOR2_X1 U496 ( .A(KEYINPUT75), .B(KEYINPUT14), .Z(n416) );
  NAND2_X1 U497 ( .A1(G234), .A2(G237), .ZN(n415) );
  XNOR2_X1 U498 ( .A(n416), .B(n415), .ZN(n417) );
  NAND2_X1 U499 ( .A1(G952), .A2(n417), .ZN(n716) );
  NOR2_X1 U500 ( .A1(G953), .A2(n716), .ZN(n541) );
  AND2_X1 U501 ( .A1(G953), .A2(n417), .ZN(n418) );
  NAND2_X1 U502 ( .A1(G902), .A2(n418), .ZN(n538) );
  NOR2_X1 U503 ( .A1(G898), .A2(n538), .ZN(n419) );
  OR2_X1 U504 ( .A1(n541), .A2(n419), .ZN(n421) );
  INV_X1 U505 ( .A(KEYINPUT87), .ZN(n420) );
  INV_X1 U506 ( .A(KEYINPUT84), .ZN(n423) );
  XNOR2_X1 U507 ( .A(n423), .B(KEYINPUT0), .ZN(n424) );
  XNOR2_X2 U508 ( .A(n425), .B(n424), .ZN(n521) );
  XNOR2_X1 U509 ( .A(G137), .B(G134), .ZN(n426) );
  XNOR2_X1 U510 ( .A(n427), .B(n426), .ZN(n737) );
  XNOR2_X1 U511 ( .A(G146), .B(n737), .ZN(n428) );
  XOR2_X1 U512 ( .A(G140), .B(n429), .Z(n431) );
  NAND2_X1 U513 ( .A1(G227), .A2(n746), .ZN(n430) );
  XNOR2_X1 U514 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U515 ( .A(n464), .B(n432), .ZN(n653) );
  XOR2_X1 U516 ( .A(KEYINPUT72), .B(G469), .Z(n433) );
  XNOR2_X2 U517 ( .A(n434), .B(n433), .ZN(n545) );
  XNOR2_X1 U518 ( .A(KEYINPUT65), .B(KEYINPUT1), .ZN(n435) );
  NAND2_X1 U519 ( .A1(G234), .A2(n746), .ZN(n436) );
  XNOR2_X1 U520 ( .A(n437), .B(n436), .ZN(n438) );
  XNOR2_X1 U521 ( .A(KEYINPUT80), .B(n438), .ZN(n484) );
  NAND2_X1 U522 ( .A1(G221), .A2(n484), .ZN(n441) );
  XOR2_X1 U523 ( .A(G110), .B(G137), .Z(n439) );
  XNOR2_X1 U524 ( .A(n439), .B(n394), .ZN(n440) );
  XNOR2_X1 U525 ( .A(n441), .B(n440), .ZN(n448) );
  XOR2_X1 U526 ( .A(KEYINPUT69), .B(KEYINPUT10), .Z(n444) );
  XNOR2_X1 U527 ( .A(n442), .B(G140), .ZN(n443) );
  XNOR2_X1 U528 ( .A(n444), .B(n443), .ZN(n736) );
  XOR2_X1 U529 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n446) );
  XNOR2_X1 U530 ( .A(KEYINPUT73), .B(KEYINPUT24), .ZN(n445) );
  NAND2_X1 U531 ( .A1(n645), .A2(n500), .ZN(n453) );
  NAND2_X1 U532 ( .A1(n599), .A2(G234), .ZN(n449) );
  XNOR2_X1 U533 ( .A(n449), .B(KEYINPUT20), .ZN(n454) );
  NAND2_X1 U534 ( .A1(G217), .A2(n454), .ZN(n451) );
  INV_X1 U535 ( .A(KEYINPUT25), .ZN(n450) );
  XNOR2_X1 U536 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U537 ( .A(n453), .B(n452), .ZN(n509) );
  NAND2_X1 U538 ( .A1(G221), .A2(n454), .ZN(n455) );
  XNOR2_X1 U539 ( .A(n455), .B(KEYINPUT21), .ZN(n699) );
  INV_X1 U540 ( .A(n699), .ZN(n505) );
  NAND2_X1 U541 ( .A1(n509), .A2(n505), .ZN(n457) );
  INV_X1 U542 ( .A(KEYINPUT67), .ZN(n456) );
  INV_X1 U543 ( .A(n695), .ZN(n458) );
  NAND2_X1 U544 ( .A1(n508), .A2(n458), .ZN(n523) );
  INV_X1 U545 ( .A(n523), .ZN(n467) );
  XOR2_X1 U546 ( .A(KEYINPUT76), .B(KEYINPUT5), .Z(n460) );
  NOR2_X1 U547 ( .A1(G953), .A2(G237), .ZN(n489) );
  NAND2_X1 U548 ( .A1(n489), .A2(G210), .ZN(n459) );
  XNOR2_X1 U549 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U550 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U551 ( .A(n464), .B(n463), .ZN(n640) );
  XNOR2_X2 U552 ( .A(n465), .B(G472), .ZN(n702) );
  NAND2_X1 U553 ( .A1(n467), .A2(n466), .ZN(n470) );
  INV_X1 U554 ( .A(KEYINPUT102), .ZN(n468) );
  XNOR2_X1 U555 ( .A(n468), .B(KEYINPUT33), .ZN(n469) );
  XNOR2_X1 U556 ( .A(n470), .B(n469), .ZN(n682) );
  INV_X1 U557 ( .A(KEYINPUT34), .ZN(n472) );
  XOR2_X1 U558 ( .A(KEYINPUT97), .B(KEYINPUT96), .Z(n474) );
  XNOR2_X1 U559 ( .A(KEYINPUT9), .B(KEYINPUT94), .ZN(n473) );
  XNOR2_X1 U560 ( .A(n474), .B(n473), .ZN(n478) );
  XOR2_X1 U561 ( .A(KEYINPUT93), .B(KEYINPUT7), .Z(n476) );
  XNOR2_X1 U562 ( .A(KEYINPUT98), .B(KEYINPUT95), .ZN(n475) );
  XNOR2_X1 U563 ( .A(n476), .B(n475), .ZN(n477) );
  XNOR2_X1 U564 ( .A(n478), .B(n477), .ZN(n482) );
  XOR2_X1 U565 ( .A(G122), .B(G107), .Z(n480) );
  XNOR2_X1 U566 ( .A(G116), .B(G134), .ZN(n479) );
  XNOR2_X1 U567 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U568 ( .A(n482), .B(n481), .ZN(n487) );
  NAND2_X1 U569 ( .A1(n484), .A2(G217), .ZN(n485) );
  XNOR2_X1 U570 ( .A(n483), .B(n485), .ZN(n486) );
  XNOR2_X1 U571 ( .A(n487), .B(n486), .ZN(n608) );
  NAND2_X1 U572 ( .A1(n608), .A2(n500), .ZN(n488) );
  INV_X1 U573 ( .A(G478), .ZN(n607) );
  XNOR2_X1 U574 ( .A(n488), .B(n607), .ZN(n528) );
  INV_X1 U575 ( .A(n528), .ZN(n503) );
  XOR2_X1 U576 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n491) );
  NAND2_X1 U577 ( .A1(G214), .A2(n489), .ZN(n490) );
  XNOR2_X1 U578 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U579 ( .A(n492), .B(G122), .Z(n498) );
  XOR2_X1 U580 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n494) );
  XNOR2_X1 U581 ( .A(G131), .B(G104), .ZN(n493) );
  XNOR2_X1 U582 ( .A(n494), .B(n493), .ZN(n496) );
  XOR2_X1 U583 ( .A(G113), .B(G143), .Z(n495) );
  XNOR2_X1 U584 ( .A(n496), .B(n495), .ZN(n497) );
  XNOR2_X1 U585 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U586 ( .A(n736), .B(n499), .ZN(n626) );
  NAND2_X1 U587 ( .A1(n626), .A2(n500), .ZN(n502) );
  XOR2_X1 U588 ( .A(KEYINPUT13), .B(G475), .Z(n501) );
  XNOR2_X1 U589 ( .A(n502), .B(n501), .ZN(n529) );
  AND2_X1 U590 ( .A1(n503), .A2(n529), .ZN(n584) );
  INV_X1 U591 ( .A(n529), .ZN(n504) );
  AND2_X1 U592 ( .A1(n504), .A2(n528), .ZN(n685) );
  AND2_X1 U593 ( .A1(n685), .A2(n505), .ZN(n506) );
  NAND2_X1 U594 ( .A1(n521), .A2(n506), .ZN(n507) );
  BUF_X1 U595 ( .A(n509), .Z(n566) );
  XNOR2_X1 U596 ( .A(n566), .B(KEYINPUT99), .ZN(n698) );
  AND2_X1 U597 ( .A1(n592), .A2(n698), .ZN(n510) );
  XNOR2_X1 U598 ( .A(n511), .B(KEYINPUT32), .ZN(n633) );
  NOR2_X1 U599 ( .A1(n592), .A2(n566), .ZN(n513) );
  INV_X1 U600 ( .A(KEYINPUT100), .ZN(n512) );
  INV_X1 U601 ( .A(KEYINPUT101), .ZN(n514) );
  XNOR2_X1 U602 ( .A(n515), .B(n514), .ZN(n634) );
  NAND2_X1 U603 ( .A1(n517), .A2(n516), .ZN(n519) );
  INV_X1 U604 ( .A(KEYINPUT44), .ZN(n518) );
  XNOR2_X1 U605 ( .A(n519), .B(n518), .ZN(n534) );
  OR2_X1 U606 ( .A1(n695), .A2(n545), .ZN(n550) );
  XNOR2_X1 U607 ( .A(n520), .B(KEYINPUT90), .ZN(n658) );
  BUF_X1 U608 ( .A(n521), .Z(n525) );
  INV_X1 U609 ( .A(n355), .ZN(n522) );
  OR2_X1 U610 ( .A1(n523), .A2(n522), .ZN(n705) );
  INV_X1 U611 ( .A(n705), .ZN(n524) );
  NAND2_X1 U612 ( .A1(n525), .A2(n524), .ZN(n527) );
  INV_X1 U613 ( .A(KEYINPUT31), .ZN(n526) );
  XNOR2_X1 U614 ( .A(n527), .B(n526), .ZN(n672) );
  NAND2_X1 U615 ( .A1(n658), .A2(n672), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n529), .A2(n528), .ZN(n670) );
  OR2_X1 U617 ( .A1(n529), .A2(n528), .ZN(n673) );
  NAND2_X1 U618 ( .A1(n670), .A2(n673), .ZN(n683) );
  NAND2_X1 U619 ( .A1(n530), .A2(n683), .ZN(n532) );
  NOR2_X1 U620 ( .A1(n592), .A2(n698), .ZN(n531) );
  AND2_X1 U621 ( .A1(n532), .A2(n632), .ZN(n533) );
  NAND2_X1 U622 ( .A1(n534), .A2(n533), .ZN(n535) );
  XNOR2_X1 U623 ( .A(n535), .B(KEYINPUT45), .ZN(n603) );
  INV_X1 U624 ( .A(KEYINPUT82), .ZN(n537) );
  XOR2_X1 U625 ( .A(KEYINPUT103), .B(n538), .Z(n539) );
  NOR2_X1 U626 ( .A1(G900), .A2(n539), .ZN(n540) );
  NOR2_X1 U627 ( .A1(n541), .A2(n540), .ZN(n542) );
  XOR2_X1 U628 ( .A(KEYINPUT77), .B(n542), .Z(n551) );
  NOR2_X1 U629 ( .A1(n551), .A2(n699), .ZN(n543) );
  XNOR2_X1 U630 ( .A(n543), .B(KEYINPUT71), .ZN(n569) );
  OR2_X1 U631 ( .A1(n569), .A2(n554), .ZN(n544) );
  INV_X1 U632 ( .A(n545), .ZN(n546) );
  XOR2_X1 U633 ( .A(KEYINPUT41), .B(KEYINPUT106), .Z(n548) );
  NAND2_X1 U634 ( .A1(n687), .A2(n686), .ZN(n547) );
  XNOR2_X1 U635 ( .A(n549), .B(KEYINPUT42), .ZN(n753) );
  INV_X1 U636 ( .A(n550), .ZN(n553) );
  INV_X1 U637 ( .A(n551), .ZN(n552) );
  NAND2_X1 U638 ( .A1(n553), .A2(n552), .ZN(n558) );
  INV_X1 U639 ( .A(n554), .ZN(n555) );
  NAND2_X1 U640 ( .A1(n555), .A2(n686), .ZN(n556) );
  XNOR2_X1 U641 ( .A(n556), .B(KEYINPUT30), .ZN(n557) );
  XNOR2_X1 U642 ( .A(n561), .B(KEYINPUT46), .ZN(n588) );
  AND2_X1 U643 ( .A1(n683), .A2(KEYINPUT74), .ZN(n564) );
  NAND2_X1 U644 ( .A1(n575), .A2(n564), .ZN(n565) );
  NAND2_X1 U645 ( .A1(n565), .A2(KEYINPUT47), .ZN(n581) );
  INV_X1 U646 ( .A(n592), .ZN(n696) );
  INV_X1 U647 ( .A(n566), .ZN(n567) );
  NAND2_X1 U648 ( .A1(n567), .A2(n686), .ZN(n568) );
  NOR2_X1 U649 ( .A1(n569), .A2(n568), .ZN(n571) );
  NAND2_X1 U650 ( .A1(n571), .A2(n570), .ZN(n593) );
  NOR2_X1 U651 ( .A1(n593), .A2(n596), .ZN(n573) );
  XOR2_X1 U652 ( .A(KEYINPUT36), .B(n573), .Z(n574) );
  NOR2_X1 U653 ( .A1(n696), .A2(n574), .ZN(n675) );
  INV_X1 U654 ( .A(n575), .ZN(n668) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(n683), .ZN(n577) );
  INV_X1 U656 ( .A(KEYINPUT47), .ZN(n576) );
  NAND2_X1 U657 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U658 ( .A1(n668), .A2(n578), .ZN(n579) );
  NOR2_X1 U659 ( .A1(n675), .A2(n579), .ZN(n580) );
  NAND2_X1 U660 ( .A1(n581), .A2(n580), .ZN(n587) );
  NAND2_X1 U661 ( .A1(n582), .A2(n389), .ZN(n583) );
  XOR2_X1 U662 ( .A(KEYINPUT104), .B(n583), .Z(n585) );
  NAND2_X1 U663 ( .A1(n585), .A2(n584), .ZN(n667) );
  NOR2_X1 U664 ( .A1(n589), .A2(n673), .ZN(n591) );
  INV_X1 U665 ( .A(KEYINPUT107), .ZN(n590) );
  XNOR2_X1 U666 ( .A(n591), .B(n590), .ZN(n750) );
  OR2_X1 U667 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U668 ( .A(KEYINPUT43), .B(n594), .ZN(n595) );
  AND2_X1 U669 ( .A1(n596), .A2(n595), .ZN(n637) );
  NOR2_X1 U670 ( .A1(n750), .A2(n637), .ZN(n597) );
  INV_X1 U671 ( .A(KEYINPUT2), .ZN(n598) );
  OR2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n601), .A2(n600), .ZN(n606) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT83), .ZN(n605) );
  BUF_X1 U675 ( .A(n603), .Z(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n677) );
  XNOR2_X1 U677 ( .A(n608), .B(KEYINPUT119), .ZN(n609) );
  XNOR2_X1 U678 ( .A(n610), .B(n609), .ZN(n612) );
  INV_X1 U679 ( .A(G952), .ZN(n611) );
  NAND2_X1 U680 ( .A1(n611), .A2(G953), .ZN(n648) );
  NAND2_X1 U681 ( .A1(n612), .A2(n648), .ZN(n614) );
  XNOR2_X1 U682 ( .A(n614), .B(n613), .ZN(G63) );
  NAND2_X1 U683 ( .A1(n638), .A2(G210), .ZN(n621) );
  BUF_X1 U684 ( .A(n615), .Z(n616) );
  XOR2_X1 U685 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n618) );
  XNOR2_X1 U686 ( .A(KEYINPUT55), .B(KEYINPUT78), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n618), .B(n617), .ZN(n619) );
  XNOR2_X1 U688 ( .A(n616), .B(n619), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n621), .B(n620), .ZN(n622) );
  NAND2_X1 U690 ( .A1(n622), .A2(n648), .ZN(n624) );
  INV_X1 U691 ( .A(KEYINPUT56), .ZN(n623) );
  XNOR2_X1 U692 ( .A(n624), .B(n623), .ZN(G51) );
  NAND2_X1 U693 ( .A1(n638), .A2(G475), .ZN(n628) );
  XNOR2_X1 U694 ( .A(KEYINPUT85), .B(KEYINPUT59), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U696 ( .A(n628), .B(n627), .ZN(n629) );
  NAND2_X1 U697 ( .A1(n629), .A2(n648), .ZN(n631) );
  INV_X1 U698 ( .A(KEYINPUT60), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n631), .B(n630), .ZN(G60) );
  XNOR2_X1 U700 ( .A(n632), .B(G101), .ZN(G3) );
  XNOR2_X1 U701 ( .A(n633), .B(G119), .ZN(G21) );
  XNOR2_X1 U702 ( .A(n634), .B(G110), .ZN(G12) );
  NOR2_X1 U703 ( .A1(n658), .A2(n670), .ZN(n635) );
  XOR2_X1 U704 ( .A(G104), .B(n635), .Z(G6) );
  XOR2_X1 U705 ( .A(n636), .B(G122), .Z(G24) );
  XOR2_X1 U706 ( .A(n637), .B(G140), .Z(G42) );
  NAND2_X1 U707 ( .A1(n638), .A2(G472), .ZN(n642) );
  XOR2_X1 U708 ( .A(KEYINPUT108), .B(KEYINPUT62), .Z(n639) );
  XNOR2_X1 U709 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U710 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U711 ( .A1(n643), .A2(n648), .ZN(n644) );
  XNOR2_X1 U712 ( .A(n644), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U713 ( .A1(n650), .A2(G217), .ZN(n647) );
  XNOR2_X1 U714 ( .A(n645), .B(KEYINPUT121), .ZN(n646) );
  XNOR2_X1 U715 ( .A(n647), .B(n646), .ZN(n649) );
  INV_X1 U716 ( .A(n648), .ZN(n656) );
  NOR2_X1 U717 ( .A1(n649), .A2(n656), .ZN(G66) );
  NAND2_X1 U718 ( .A1(n650), .A2(G469), .ZN(n655) );
  XOR2_X1 U719 ( .A(KEYINPUT118), .B(KEYINPUT57), .Z(n651) );
  XNOR2_X1 U720 ( .A(n651), .B(KEYINPUT58), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(n654) );
  XNOR2_X1 U722 ( .A(n655), .B(n654), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n657), .A2(n656), .ZN(G54) );
  NOR2_X1 U724 ( .A1(n658), .A2(n673), .ZN(n660) );
  XNOR2_X1 U725 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n659) );
  XNOR2_X1 U726 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U727 ( .A(G107), .B(n661), .ZN(G9) );
  NOR2_X1 U728 ( .A1(n668), .A2(n673), .ZN(n665) );
  XOR2_X1 U729 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n663) );
  XNOR2_X1 U730 ( .A(G128), .B(KEYINPUT29), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(n664), .ZN(G30) );
  XOR2_X1 U733 ( .A(G143), .B(KEYINPUT111), .Z(n666) );
  XNOR2_X1 U734 ( .A(n667), .B(n666), .ZN(G45) );
  NOR2_X1 U735 ( .A1(n668), .A2(n670), .ZN(n669) );
  XOR2_X1 U736 ( .A(G146), .B(n669), .Z(G48) );
  NOR2_X1 U737 ( .A1(n670), .A2(n672), .ZN(n671) );
  XOR2_X1 U738 ( .A(G113), .B(n671), .Z(G15) );
  NOR2_X1 U739 ( .A1(n673), .A2(n672), .ZN(n674) );
  XOR2_X1 U740 ( .A(G116), .B(n674), .Z(G18) );
  XNOR2_X1 U741 ( .A(G125), .B(n675), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n676), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U743 ( .A(KEYINPUT116), .B(KEYINPUT53), .Z(n723) );
  INV_X1 U744 ( .A(n677), .ZN(n680) );
  XOR2_X1 U745 ( .A(KEYINPUT79), .B(KEYINPUT2), .Z(n678) );
  NOR2_X1 U746 ( .A1(n351), .A2(n678), .ZN(n679) );
  NOR2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U748 ( .A1(G953), .A2(n681), .ZN(n721) );
  NOR2_X1 U749 ( .A1(n693), .A2(n709), .ZN(n719) );
  XOR2_X1 U750 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n715) );
  AND2_X1 U751 ( .A1(n684), .A2(n683), .ZN(n691) );
  INV_X1 U752 ( .A(n685), .ZN(n689) );
  NOR2_X1 U753 ( .A1(n687), .A2(n686), .ZN(n688) );
  NOR2_X1 U754 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U755 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U756 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U757 ( .A(KEYINPUT113), .B(n694), .Z(n712) );
  NAND2_X1 U758 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U759 ( .A(n697), .B(KEYINPUT50), .ZN(n704) );
  NAND2_X1 U760 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U761 ( .A(KEYINPUT49), .B(n700), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n355), .A2(n701), .ZN(n703) );
  NAND2_X1 U763 ( .A1(n704), .A2(n703), .ZN(n706) );
  NAND2_X1 U764 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U765 ( .A(KEYINPUT51), .B(n707), .ZN(n708) );
  NOR2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U767 ( .A(KEYINPUT112), .B(n710), .ZN(n711) );
  NOR2_X1 U768 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U769 ( .A(n713), .B(KEYINPUT52), .ZN(n714) );
  XNOR2_X1 U770 ( .A(n715), .B(n714), .ZN(n717) );
  NOR2_X1 U771 ( .A1(n717), .A2(n716), .ZN(n718) );
  NOR2_X1 U772 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XNOR2_X1 U774 ( .A(n723), .B(n722), .ZN(G75) );
  NAND2_X1 U775 ( .A1(n604), .A2(n746), .ZN(n727) );
  NAND2_X1 U776 ( .A1(G953), .A2(G224), .ZN(n724) );
  XNOR2_X1 U777 ( .A(KEYINPUT61), .B(n724), .ZN(n725) );
  NAND2_X1 U778 ( .A1(n725), .A2(G898), .ZN(n726) );
  NAND2_X1 U779 ( .A1(n727), .A2(n726), .ZN(n733) );
  XNOR2_X1 U780 ( .A(G101), .B(n728), .ZN(n729) );
  XNOR2_X1 U781 ( .A(n729), .B(KEYINPUT122), .ZN(n731) );
  NOR2_X1 U782 ( .A1(G898), .A2(n746), .ZN(n730) );
  NOR2_X1 U783 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U784 ( .A(n733), .B(n732), .ZN(n734) );
  XOR2_X1 U785 ( .A(KEYINPUT123), .B(n734), .Z(G69) );
  XNOR2_X1 U786 ( .A(n737), .B(n736), .ZN(n738) );
  XNOR2_X1 U787 ( .A(n738), .B(KEYINPUT124), .ZN(n739) );
  XNOR2_X1 U788 ( .A(n735), .B(n739), .ZN(n743) );
  XNOR2_X1 U789 ( .A(n743), .B(G227), .ZN(n740) );
  NAND2_X1 U790 ( .A1(n740), .A2(G900), .ZN(n741) );
  NAND2_X1 U791 ( .A1(G953), .A2(n741), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n742), .B(KEYINPUT126), .ZN(n749) );
  XOR2_X1 U793 ( .A(KEYINPUT125), .B(n743), .Z(n745) );
  XOR2_X1 U794 ( .A(n745), .B(n744), .Z(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n749), .A2(n748), .ZN(G72) );
  XOR2_X1 U797 ( .A(G134), .B(n750), .Z(G36) );
  XNOR2_X1 U798 ( .A(G131), .B(KEYINPUT127), .ZN(n752) );
  XNOR2_X1 U799 ( .A(n752), .B(n751), .ZN(G33) );
  XOR2_X1 U800 ( .A(n753), .B(G137), .Z(G39) );
endmodule

