//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 1 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1217, new_n1218, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1277, new_n1278;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G77), .ZN(new_n202));
  AND2_X1   g0002(.A1(new_n201), .A2(new_n202), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(G257), .ZN(new_n209));
  INV_X1    g0009(.A(G264), .ZN(new_n210));
  AOI211_X1 g0010(.A(new_n205), .B(new_n208), .C1(new_n209), .C2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G1), .A2(G13), .ZN(new_n213));
  INV_X1    g0013(.A(KEYINPUT64), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g0015(.A1(KEYINPUT64), .A2(G1), .A3(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G20), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(G50), .B1(G58), .B2(G68), .ZN(new_n221));
  INV_X1    g0021(.A(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n211), .A2(KEYINPUT0), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n212), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT65), .Z(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G68), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  INV_X1    g0029(.A(G87), .ZN(new_n230));
  OAI221_X1 g0030(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n205), .ZN(new_n231));
  AOI22_X1  g0031(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n232));
  INV_X1    g0032(.A(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G107), .ZN(new_n234));
  OAI221_X1 g0034(.A(new_n232), .B1(new_n202), .B2(new_n233), .C1(new_n234), .C2(new_n210), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n206), .B1(new_n231), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(KEYINPUT1), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n226), .A2(new_n237), .ZN(G361));
  XOR2_X1   g0038(.A(G238), .B(G244), .Z(new_n239));
  XNOR2_X1  g0039(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G226), .B(G232), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n228), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n250), .B(new_n256), .ZN(G351));
  NAND2_X1  g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G1), .A3(G13), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n259), .A2(G274), .ZN(new_n260));
  INV_X1    g0060(.A(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n213), .B1(G33), .B2(G41), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n263), .ZN(new_n266));
  AND2_X1   g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n268), .A2(G1698), .ZN(new_n271));
  INV_X1    g0071(.A(G223), .ZN(new_n272));
  OAI221_X1 g0072(.A(new_n270), .B1(new_n202), .B2(new_n268), .C1(new_n271), .C2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n217), .A2(new_n258), .ZN(new_n274));
  INV_X1    g0074(.A(new_n274), .ZN(new_n275));
  AOI211_X1 g0075(.A(new_n264), .B(new_n267), .C1(new_n273), .C2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n215), .A2(new_n216), .A3(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n219), .A2(new_n279), .A3(KEYINPUT67), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT67), .ZN(new_n281));
  OAI21_X1  g0081(.A(new_n281), .B1(G20), .B2(G33), .ZN(new_n282));
  AND2_X1   g0082(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g0085(.A(KEYINPUT8), .B(G58), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n219), .A2(G33), .ZN(new_n287));
  OAI22_X1  g0087(.A1(new_n286), .A2(new_n287), .B1(new_n219), .B2(new_n201), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n278), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G1), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n290), .A2(G13), .A3(G20), .ZN(new_n291));
  NAND4_X1  g0091(.A1(new_n215), .A2(new_n291), .A3(new_n216), .A4(new_n277), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n219), .A2(G1), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(G50), .A3(new_n295), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n289), .B(new_n296), .C1(G50), .C2(new_n291), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT9), .ZN(new_n298));
  AOI22_X1  g0098(.A1(new_n276), .A2(G190), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G200), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n299), .B1(new_n298), .B2(new_n297), .C1(new_n300), .C2(new_n276), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT10), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT70), .B(KEYINPUT10), .Z(new_n303));
  OAI211_X1 g0103(.A(new_n302), .B(KEYINPUT71), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  OR3_X1    g0104(.A1(new_n301), .A2(KEYINPUT71), .A3(new_n303), .ZN(new_n305));
  AND2_X1   g0105(.A1(KEYINPUT68), .A2(G179), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT68), .A2(G179), .ZN(new_n307));
  NOR2_X1   g0107(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n276), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n297), .C1(G169), .C2(new_n276), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n304), .A2(new_n305), .A3(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n264), .B1(G244), .B2(new_n266), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n313));
  OAI221_X1 g0113(.A(new_n313), .B1(new_n234), .B2(new_n268), .C1(new_n271), .C2(new_n229), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(new_n275), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  INV_X1    g0116(.A(G169), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n278), .ZN(new_n319));
  XOR2_X1   g0119(.A(new_n286), .B(KEYINPUT69), .Z(new_n320));
  INV_X1    g0120(.A(new_n283), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  XOR2_X1   g0122(.A(KEYINPUT15), .B(G87), .Z(new_n323));
  INV_X1    g0123(.A(new_n287), .ZN(new_n324));
  AOI22_X1  g0124(.A1(new_n323), .A2(new_n324), .B1(G20), .B2(G77), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n319), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n294), .A2(new_n202), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n292), .B1(G77), .B2(new_n291), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n318), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n308), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n316), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n326), .A2(new_n329), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n316), .A2(G200), .ZN(new_n336));
  INV_X1    g0136(.A(G190), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n316), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n334), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n311), .A2(new_n339), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n324), .A2(G77), .B1(G20), .B2(new_n228), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT73), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n342), .B1(new_n321), .B2(G50), .ZN(new_n343));
  NOR3_X1   g0143(.A1(new_n283), .A2(KEYINPUT73), .A3(new_n251), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n341), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n345), .A2(KEYINPUT11), .A3(new_n278), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n292), .A2(new_n228), .A3(new_n294), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT74), .ZN(new_n348));
  OAI22_X1  g0148(.A1(new_n291), .A2(G68), .B1(new_n348), .B2(KEYINPUT12), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT12), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(KEYINPUT74), .B2(new_n350), .ZN(new_n351));
  OAI211_X1 g0151(.A(new_n348), .B(KEYINPUT12), .C1(new_n291), .C2(G68), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n346), .A2(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT11), .B1(new_n345), .B2(new_n278), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT14), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n268), .A2(G232), .A3(G1698), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n268), .A2(G226), .A3(new_n269), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT72), .A4(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n364), .A2(new_n275), .A3(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT13), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n264), .B1(G238), .B2(new_n266), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n367), .B1(new_n366), .B2(new_n368), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n358), .B(G169), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n366), .A2(new_n368), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(KEYINPUT13), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n366), .A2(new_n367), .A3(new_n368), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(G179), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n373), .A2(new_n374), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n358), .B1(new_n377), .B2(G169), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n357), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(G200), .B1(new_n369), .B2(new_n370), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n373), .A2(G190), .A3(new_n374), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(new_n356), .ZN(new_n382));
  INV_X1    g0182(.A(G58), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n228), .ZN(new_n384));
  NOR2_X1   g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  OAI21_X1  g0185(.A(G20), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(G159), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n386), .B1(new_n283), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT7), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n389), .B1(new_n268), .B2(G20), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n279), .A2(KEYINPUT3), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G33), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(KEYINPUT7), .A3(new_n219), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n388), .B1(G68), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n319), .B1(new_n397), .B2(KEYINPUT16), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT16), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n228), .B1(new_n390), .B2(new_n395), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n400), .B2(new_n388), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(KEYINPUT75), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT75), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n403), .B(new_n399), .C1(new_n400), .C2(new_n388), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n398), .A2(new_n402), .A3(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n286), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n295), .ZN(new_n407));
  XNOR2_X1  g0207(.A(new_n407), .B(KEYINPUT76), .ZN(new_n408));
  INV_X1    g0208(.A(new_n291), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n408), .A2(new_n293), .B1(new_n409), .B2(new_n286), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n405), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n391), .A2(new_n393), .A3(G226), .A4(G1698), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n391), .A2(new_n393), .A3(G223), .A4(new_n269), .ZN(new_n413));
  OAI211_X1 g0213(.A(new_n412), .B(new_n413), .C1(new_n279), .C2(new_n230), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(new_n275), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n266), .A2(G232), .B1(new_n260), .B2(new_n263), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n415), .A2(new_n416), .A3(new_n331), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n317), .B1(new_n415), .B2(new_n416), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n411), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n419), .B1(new_n405), .B2(new_n410), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n422), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n415), .A2(new_n416), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n300), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n428), .B1(G190), .B2(new_n427), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n405), .A2(new_n429), .A3(new_n410), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT17), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n405), .A2(new_n429), .A3(KEYINPUT17), .A4(new_n410), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT77), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(KEYINPUT77), .A3(new_n433), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n426), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n340), .A2(new_n379), .A3(new_n382), .A4(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n262), .A2(G1), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n441), .A2(new_n205), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n259), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT78), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT78), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n290), .A2(G45), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n259), .A2(new_n445), .A3(G250), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(KEYINPUT79), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n259), .A2(G274), .A3(new_n441), .ZN(new_n449));
  NAND4_X1  g0249(.A1(new_n444), .A2(new_n447), .A3(new_n448), .A4(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n449), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n445), .B1(new_n442), .B2(new_n259), .ZN(new_n452));
  OAI21_X1  g0252(.A(KEYINPUT79), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n450), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n233), .A2(new_n269), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n268), .A2(new_n455), .B1(G33), .B2(G116), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n268), .A2(G238), .A3(new_n269), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n274), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n308), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n460), .A2(KEYINPUT80), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n458), .B1(new_n450), .B2(new_n453), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT80), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n462), .A2(new_n463), .A3(new_n308), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n461), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n323), .A2(new_n291), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT19), .ZN(new_n467));
  OAI21_X1  g0267(.A(new_n219), .B1(new_n361), .B2(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(G97), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n230), .A2(new_n469), .A3(new_n234), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n391), .A2(new_n393), .A3(new_n219), .A4(G68), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n467), .B1(new_n287), .B2(new_n469), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT81), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n319), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT81), .A4(new_n473), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n466), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n292), .B1(new_n290), .B2(G33), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(new_n323), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT82), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n478), .A2(KEYINPUT82), .A3(new_n480), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n454), .A2(new_n459), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n317), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n465), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n391), .A2(new_n393), .A3(G244), .A4(new_n269), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT4), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n269), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n493));
  NAND2_X1  g0293(.A1(G33), .A2(G283), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n493), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(new_n275), .ZN(new_n496));
  XNOR2_X1  g0296(.A(KEYINPUT5), .B(G41), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n497), .A2(new_n259), .A3(G274), .A4(new_n441), .ZN(new_n498));
  AND2_X1   g0298(.A1(KEYINPUT5), .A2(G41), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT5), .A2(G41), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n441), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n259), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n498), .B1(new_n502), .B2(new_n209), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n496), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT6), .ZN(new_n507));
  NOR3_X1   g0307(.A1(new_n507), .A2(new_n469), .A3(G107), .ZN(new_n508));
  XNOR2_X1  g0308(.A(G97), .B(G107), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  OAI22_X1  g0310(.A1(new_n510), .A2(new_n219), .B1(new_n202), .B2(new_n283), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n234), .B1(new_n390), .B2(new_n395), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n278), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n291), .A2(G97), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n514), .B1(new_n479), .B2(G97), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n503), .B1(new_n495), .B2(new_n275), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G190), .ZN(new_n517));
  NAND4_X1  g0317(.A1(new_n506), .A2(new_n513), .A3(new_n515), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n505), .A2(new_n317), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n513), .A2(new_n515), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n308), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n486), .A2(G200), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n479), .A2(G87), .ZN(new_n525));
  AND2_X1   g0325(.A1(new_n478), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n462), .A2(G190), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n524), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  AND3_X1   g0328(.A1(new_n488), .A2(new_n523), .A3(new_n528), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n391), .A2(new_n393), .A3(new_n219), .A4(G87), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT22), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT22), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n268), .A2(new_n532), .A3(new_n219), .A4(G87), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(G116), .ZN(new_n535));
  NOR3_X1   g0335(.A1(new_n279), .A2(new_n535), .A3(G20), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT23), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(G20), .B2(new_n234), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n219), .A2(KEYINPUT23), .A3(G107), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n541));
  NOR4_X1   g0341(.A1(new_n536), .A2(new_n538), .A3(new_n539), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n543));
  INV_X1    g0343(.A(new_n543), .ZN(new_n544));
  AND3_X1   g0344(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g0345(.A(new_n544), .B1(new_n534), .B2(new_n542), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n278), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n409), .A2(new_n234), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT25), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n549), .B1(G107), .B2(new_n479), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n547), .A2(new_n550), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n391), .A2(new_n393), .A3(G250), .A4(new_n269), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT85), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT85), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n268), .A2(new_n554), .A3(G250), .A4(new_n269), .ZN(new_n555));
  XNOR2_X1  g0355(.A(KEYINPUT86), .B(G294), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G33), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n268), .A2(G257), .A3(G1698), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n553), .A2(new_n555), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(new_n275), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n501), .A2(G264), .A3(new_n259), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(new_n498), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n564), .A2(KEYINPUT87), .A3(G169), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n562), .B1(new_n559), .B2(new_n275), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G179), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g0368(.A(KEYINPUT87), .B1(new_n564), .B2(G169), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n551), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n268), .A2(G264), .A3(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n394), .A2(G303), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n391), .A2(new_n393), .A3(G257), .A4(new_n269), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n265), .B1(new_n441), .B2(new_n497), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n574), .A2(new_n275), .B1(G270), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n317), .B1(new_n576), .B2(new_n498), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n479), .A2(G116), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n409), .A2(new_n535), .ZN(new_n579));
  AOI21_X1  g0379(.A(G20), .B1(G33), .B2(G283), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n279), .A2(G97), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n580), .A2(new_n581), .B1(G20), .B2(new_n535), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n582), .A2(new_n278), .A3(KEYINPUT20), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT20), .B1(new_n582), .B2(new_n278), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n578), .B(new_n579), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n577), .A2(KEYINPUT21), .A3(new_n586), .ZN(new_n587));
  NAND4_X1  g0387(.A1(new_n586), .A2(G179), .A3(new_n498), .A4(new_n576), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT21), .B1(new_n577), .B2(new_n586), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT83), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n574), .A2(new_n275), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n575), .A2(G270), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(G190), .A3(new_n498), .A4(new_n594), .ZN(new_n595));
  OR2_X1    g0395(.A1(new_n584), .A2(new_n585), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n595), .A2(new_n578), .A3(new_n596), .A4(new_n579), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n300), .B1(new_n576), .B2(new_n498), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n592), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(new_n598), .ZN(new_n600));
  INV_X1    g0400(.A(new_n586), .ZN(new_n601));
  NAND4_X1  g0401(.A1(new_n600), .A2(new_n601), .A3(KEYINPUT83), .A4(new_n595), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n599), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n566), .A2(new_n337), .ZN(new_n604));
  OAI211_X1 g0404(.A(new_n604), .B(KEYINPUT88), .C1(G200), .C2(new_n566), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT88), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n564), .A2(new_n606), .A3(new_n300), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n605), .A2(new_n547), .A3(new_n550), .A4(new_n607), .ZN(new_n608));
  AND4_X1   g0408(.A1(new_n570), .A2(new_n591), .A3(new_n603), .A4(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n440), .A2(new_n529), .A3(new_n609), .ZN(G372));
  NAND2_X1  g0410(.A1(new_n382), .A2(new_n333), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n436), .A2(new_n437), .B1(new_n379), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n422), .A2(KEYINPUT91), .A3(new_n425), .ZN(new_n613));
  INV_X1    g0413(.A(KEYINPUT91), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n423), .A2(new_n424), .ZN(new_n615));
  AOI211_X1 g0415(.A(KEYINPUT18), .B(new_n419), .C1(new_n405), .C2(new_n410), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n304), .B(new_n305), .C1(new_n612), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n310), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT89), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n476), .A2(new_n477), .ZN(new_n623));
  INV_X1    g0423(.A(new_n466), .ZN(new_n624));
  AND4_X1   g0424(.A1(KEYINPUT82), .A2(new_n623), .A3(new_n624), .A4(new_n480), .ZN(new_n625));
  AOI21_X1  g0425(.A(KEYINPUT82), .B1(new_n478), .B2(new_n480), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n460), .B1(G169), .B2(new_n462), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n622), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AOI211_X1 g0429(.A(new_n331), .B(new_n458), .C1(new_n450), .C2(new_n453), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n630), .B1(new_n317), .B2(new_n486), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n485), .A2(new_n631), .A3(KEYINPUT89), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n528), .B1(new_n627), .B2(new_n628), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n607), .A2(new_n547), .A3(new_n550), .ZN(new_n635));
  OAI21_X1  g0435(.A(KEYINPUT88), .B1(new_n566), .B2(G200), .ZN(new_n636));
  AOI211_X1 g0436(.A(G190), .B(new_n562), .C1(new_n559), .C2(new_n275), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n522), .B(new_n518), .C1(new_n635), .C2(new_n638), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n634), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n591), .A2(new_n570), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n633), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT26), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n634), .B2(new_n522), .ZN(new_n644));
  INV_X1    g0444(.A(new_n522), .ZN(new_n645));
  XNOR2_X1  g0445(.A(KEYINPUT90), .B(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n488), .A2(new_n528), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n644), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n621), .B1(new_n440), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n651), .B(KEYINPUT92), .ZN(G369));
  NAND2_X1  g0452(.A1(new_n591), .A2(new_n603), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n290), .A2(new_n219), .A3(G13), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  INV_X1    g0456(.A(G213), .ZN(new_n657));
  NOR3_X1   g0457(.A1(new_n655), .A2(new_n656), .A3(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n658), .A2(G343), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n586), .A2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT93), .Z(new_n662));
  AND2_X1   g0462(.A1(new_n653), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g0463(.A1(new_n662), .A2(new_n590), .A3(new_n589), .ZN(new_n664));
  OR3_X1    g0464(.A1(new_n663), .A2(KEYINPUT94), .A3(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(KEYINPUT94), .B1(new_n663), .B2(new_n664), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND2_X1   g0469(.A1(new_n570), .A2(new_n608), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n551), .A2(new_n660), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n570), .B2(new_n659), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n669), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n570), .A2(new_n660), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n591), .A2(new_n660), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n674), .A2(new_n677), .ZN(G399));
  NOR2_X1   g0478(.A1(new_n208), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n470), .A2(G116), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(G1), .A3(new_n681), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n682), .B1(new_n221), .B2(new_n680), .ZN(new_n683));
  XOR2_X1   g0483(.A(KEYINPUT95), .B(KEYINPUT28), .Z(new_n684));
  XNOR2_X1  g0484(.A(new_n683), .B(new_n684), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n454), .A2(new_n516), .A3(new_n459), .A4(new_n576), .ZN(new_n686));
  INV_X1    g0486(.A(KEYINPUT30), .ZN(new_n687));
  NOR3_X1   g0487(.A1(new_n686), .A2(new_n687), .A3(new_n567), .ZN(new_n688));
  AND3_X1   g0488(.A1(new_n454), .A2(new_n459), .A3(new_n576), .ZN(new_n689));
  INV_X1    g0489(.A(new_n567), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n689), .A2(KEYINPUT96), .A3(new_n690), .A4(new_n516), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT96), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n692), .B1(new_n686), .B2(new_n567), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n687), .A3(new_n693), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n516), .A2(new_n566), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n576), .A2(new_n498), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(new_n486), .A3(new_n308), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT97), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n688), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n694), .A2(KEYINPUT97), .A3(new_n697), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n609), .A2(new_n529), .A3(new_n659), .ZN(new_n704));
  INV_X1    g0504(.A(new_n688), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n694), .A2(new_n705), .A3(new_n697), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(new_n660), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT31), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(KEYINPUT98), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT98), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n711), .B1(new_n707), .B2(new_n708), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n703), .B(new_n704), .C1(new_n710), .C2(new_n712), .ZN(new_n713));
  AND2_X1   g0513(.A1(new_n713), .A2(G330), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n634), .A2(new_n522), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n488), .A2(new_n528), .A3(new_n645), .ZN(new_n716));
  AOI22_X1  g0516(.A1(new_n715), .A2(KEYINPUT26), .B1(new_n716), .B2(new_n646), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n629), .A2(new_n632), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n485), .A2(new_n631), .ZN(new_n719));
  NAND4_X1  g0519(.A1(new_n523), .A2(new_n719), .A3(new_n528), .A4(new_n608), .ZN(new_n720));
  AND2_X1   g0520(.A1(new_n591), .A2(new_n570), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n718), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n659), .B1(new_n717), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n660), .B1(new_n642), .B2(new_n649), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT29), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n724), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n714), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n685), .B1(new_n729), .B2(G1), .ZN(G364));
  INV_X1    g0530(.A(G13), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(G20), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n290), .B1(new_n732), .B2(G45), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n679), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n669), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n667), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(G330), .B2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G13), .A2(G33), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n740), .A2(G20), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n735), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n208), .A2(new_n394), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n745), .A2(G355), .B1(new_n535), .B2(new_n208), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n256), .A2(new_n262), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n208), .A2(new_n268), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n748), .B1(G45), .B2(new_n221), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n747), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n218), .B1(G20), .B2(new_n317), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(new_n741), .ZN(new_n752));
  AOI21_X1  g0552(.A(new_n744), .B1(new_n750), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n300), .A2(G179), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n219), .A2(G190), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G179), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  AOI22_X1  g0560(.A1(G283), .A2(new_n757), .B1(new_n760), .B2(G329), .ZN(new_n761));
  INV_X1    g0561(.A(G303), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n219), .A2(new_n337), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(new_n754), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n761), .B(new_n394), .C1(new_n762), .C2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n331), .A2(new_n300), .A3(new_n763), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(G322), .ZN(new_n768));
  INV_X1    g0568(.A(G311), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n331), .A2(new_n300), .A3(new_n755), .ZN(new_n770));
  INV_X1    g0570(.A(G326), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n219), .A2(new_n300), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n331), .A2(G190), .A3(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n768), .B1(new_n769), .B2(new_n770), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n219), .B1(new_n758), .B2(G190), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n765), .B(new_n774), .C1(new_n556), .C2(new_n776), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n331), .A2(new_n337), .A3(new_n772), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT100), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n778), .A2(new_n779), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  XNOR2_X1  g0583(.A(KEYINPUT33), .B(G317), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n783), .A2(G68), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n764), .A2(new_n230), .ZN(new_n787));
  OR3_X1    g0587(.A1(new_n787), .A2(KEYINPUT99), .A3(new_n394), .ZN(new_n788));
  OAI21_X1  g0588(.A(KEYINPUT99), .B1(new_n787), .B2(new_n394), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n788), .B(new_n789), .C1(new_n251), .C2(new_n773), .ZN(new_n790));
  OAI22_X1  g0590(.A1(new_n756), .A2(new_n234), .B1(new_n775), .B2(new_n469), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n760), .A2(G159), .ZN(new_n792));
  XNOR2_X1  g0592(.A(new_n792), .B(KEYINPUT32), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n383), .A2(new_n766), .B1(new_n770), .B2(new_n202), .ZN(new_n794));
  NOR4_X1   g0594(.A1(new_n790), .A2(new_n791), .A3(new_n793), .A4(new_n794), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n777), .A2(new_n785), .B1(new_n786), .B2(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(new_n751), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n753), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n738), .B1(new_n743), .B2(new_n798), .ZN(G396));
  OAI21_X1  g0599(.A(new_n338), .B1(new_n335), .B2(new_n659), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n334), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n333), .A2(new_n659), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n725), .B(new_n803), .ZN(new_n804));
  OR2_X1    g0604(.A1(new_n714), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n714), .A2(new_n804), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n805), .A2(new_n744), .A3(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n773), .ZN(new_n808));
  INV_X1    g0608(.A(new_n770), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n808), .B1(new_n809), .B2(G159), .ZN(new_n810));
  XOR2_X1   g0610(.A(KEYINPUT102), .B(G143), .Z(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n766), .B2(new_n811), .C1(new_n782), .C2(new_n284), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT34), .ZN(new_n814));
  INV_X1    g0614(.A(G132), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n268), .B1(new_n759), .B2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT103), .Z(new_n817));
  INV_X1    g0617(.A(new_n764), .ZN(new_n818));
  AOI22_X1  g0618(.A1(G50), .A2(new_n818), .B1(new_n757), .B2(G68), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n819), .B1(new_n383), .B2(new_n775), .ZN(new_n820));
  NOR3_X1   g0620(.A1(new_n814), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g0621(.A(new_n821), .B1(KEYINPUT34), .B2(new_n813), .ZN(new_n822));
  INV_X1    g0622(.A(G283), .ZN(new_n823));
  OAI22_X1  g0623(.A1(new_n782), .A2(new_n823), .B1(new_n535), .B2(new_n770), .ZN(new_n824));
  OR2_X1    g0624(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(KEYINPUT101), .ZN(new_n826));
  INV_X1    g0626(.A(G294), .ZN(new_n827));
  OAI22_X1  g0627(.A1(new_n827), .A2(new_n766), .B1(new_n773), .B2(new_n762), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n268), .B1(new_n760), .B2(G311), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n756), .A2(new_n230), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n829), .B(new_n831), .C1(new_n234), .C2(new_n764), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n828), .B(new_n832), .C1(G97), .C2(new_n776), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n825), .A2(new_n826), .A3(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n797), .B1(new_n822), .B2(new_n834), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n751), .A2(new_n739), .ZN(new_n836));
  AOI211_X1 g0636(.A(new_n744), .B(new_n835), .C1(new_n202), .C2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT104), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n837), .A2(new_n838), .B1(new_n739), .B2(new_n803), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n839), .B1(new_n838), .B2(new_n837), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n807), .A2(new_n840), .ZN(G384));
  NOR2_X1   g0641(.A1(new_n732), .A2(new_n290), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT37), .ZN(new_n843));
  AND2_X1   g0643(.A1(new_n398), .A2(new_n401), .ZN(new_n844));
  INV_X1    g0644(.A(new_n410), .ZN(new_n845));
  OAI22_X1  g0645(.A1(new_n844), .A2(new_n845), .B1(new_n420), .B2(new_n658), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n843), .B1(new_n846), .B2(new_n430), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n658), .B(KEYINPUT105), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n405), .B2(new_n410), .ZN(new_n851));
  INV_X1    g0651(.A(new_n851), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n852), .A2(new_n421), .A3(new_n430), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n848), .B1(KEYINPUT37), .B2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n844), .A2(new_n845), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(new_n658), .ZN(new_n856));
  OAI211_X1 g0656(.A(KEYINPUT38), .B(new_n854), .C1(new_n438), .C2(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n857), .A2(KEYINPUT106), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  INV_X1    g0659(.A(new_n434), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n852), .B1(new_n618), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n853), .B(new_n843), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n859), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT39), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n615), .A2(new_n616), .ZN(new_n865));
  AND3_X1   g0665(.A1(new_n432), .A2(KEYINPUT77), .A3(new_n433), .ZN(new_n866));
  AOI21_X1  g0666(.A(KEYINPUT77), .B1(new_n432), .B2(new_n433), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n865), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n856), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT106), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n870), .A2(new_n871), .A3(KEYINPUT38), .A4(new_n854), .ZN(new_n872));
  NAND4_X1  g0672(.A1(new_n858), .A2(new_n863), .A3(new_n864), .A4(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n857), .ZN(new_n874));
  AOI21_X1  g0674(.A(KEYINPUT38), .B1(new_n870), .B2(new_n854), .ZN(new_n875));
  OAI21_X1  g0675(.A(KEYINPUT39), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n369), .A2(new_n370), .ZN(new_n878));
  OAI21_X1  g0678(.A(KEYINPUT14), .B1(new_n878), .B2(new_n317), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n375), .A3(new_n371), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n880), .A2(new_n357), .A3(new_n659), .ZN(new_n881));
  INV_X1    g0681(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n877), .A2(new_n882), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n874), .A2(new_n875), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n802), .ZN(new_n886));
  INV_X1    g0686(.A(new_n803), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n725), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n382), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n357), .B(new_n660), .C1(new_n880), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n357), .A2(new_n660), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n379), .A2(new_n382), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n888), .A2(new_n894), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n885), .A2(new_n895), .B1(new_n619), .B2(new_n850), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n883), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n439), .B1(new_n724), .B2(new_n727), .ZN(new_n898));
  NOR2_X1   g0698(.A1(new_n898), .A2(new_n621), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n897), .B(new_n899), .Z(new_n900));
  INV_X1    g0700(.A(KEYINPUT40), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n706), .A2(KEYINPUT31), .A3(new_n660), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n709), .A2(new_n704), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n803), .B1(new_n890), .B2(new_n892), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n901), .B1(new_n884), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n858), .A2(new_n863), .A3(new_n872), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n905), .A2(new_n901), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AND2_X1   g0709(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n440), .A2(new_n903), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n668), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n910), .B2(new_n911), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n842), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n900), .B2(new_n913), .ZN(new_n915));
  INV_X1    g0715(.A(new_n510), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(KEYINPUT35), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(G116), .A3(new_n220), .A4(new_n918), .ZN(new_n919));
  XNOR2_X1  g0719(.A(new_n919), .B(KEYINPUT36), .ZN(new_n920));
  OAI21_X1  g0720(.A(G77), .B1(new_n383), .B2(new_n228), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n252), .B1(new_n921), .B2(new_n221), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n731), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(new_n920), .A3(new_n923), .ZN(G367));
  AOI211_X1 g0724(.A(new_n741), .B(new_n751), .C1(new_n208), .C2(new_n323), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n246), .A2(new_n748), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n744), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n526), .A2(new_n659), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n719), .A2(new_n528), .A3(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n718), .B2(new_n928), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n284), .A2(new_n766), .B1(new_n773), .B2(new_n811), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(G50), .B2(new_n809), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n268), .B1(new_n764), .B2(new_n383), .ZN(new_n933));
  INV_X1    g0733(.A(G137), .ZN(new_n934));
  OAI22_X1  g0734(.A1(new_n756), .A2(new_n202), .B1(new_n759), .B2(new_n934), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(G68), .C2(new_n776), .ZN(new_n936));
  OAI211_X1 g0736(.A(new_n932), .B(new_n936), .C1(new_n387), .C2(new_n782), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n764), .A2(new_n535), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT46), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n939), .B1(G283), .B2(new_n809), .ZN(new_n940));
  INV_X1    g0740(.A(new_n556), .ZN(new_n941));
  OAI221_X1 g0741(.A(new_n940), .B1(new_n769), .B2(new_n773), .C1(new_n941), .C2(new_n782), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n756), .A2(new_n469), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n268), .B(new_n943), .C1(G317), .C2(new_n760), .ZN(new_n944));
  OR2_X1    g0744(.A1(new_n944), .A2(KEYINPUT108), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n944), .A2(KEYINPUT108), .ZN(new_n946));
  AOI22_X1  g0746(.A1(new_n767), .A2(G303), .B1(G107), .B2(new_n776), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n937), .B1(new_n942), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT47), .Z(new_n950));
  OAI221_X1 g0750(.A(new_n927), .B1(new_n930), .B2(new_n742), .C1(new_n797), .C2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n520), .A2(new_n660), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n523), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n645), .A2(new_n660), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n677), .A2(new_n955), .ZN(new_n956));
  XOR2_X1   g0756(.A(new_n956), .B(KEYINPUT45), .Z(new_n957));
  NOR2_X1   g0757(.A1(new_n677), .A2(new_n955), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT44), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  XOR2_X1   g0760(.A(new_n960), .B(new_n674), .Z(new_n961));
  NAND2_X1  g0761(.A1(new_n670), .A2(new_n676), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n962), .B1(new_n673), .B2(new_n676), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n669), .B(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(new_n729), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n961), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n729), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n679), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n734), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n955), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(new_n962), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT42), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n522), .B1(new_n953), .B2(new_n570), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n659), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n972), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT107), .ZN(new_n976));
  AOI21_X1  g0776(.A(KEYINPUT43), .B1(new_n930), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n976), .B2(new_n930), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n930), .A2(KEYINPUT43), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  OAI21_X1  g0780(.A(new_n980), .B1(new_n978), .B2(new_n975), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n674), .A2(new_n970), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n981), .B(new_n982), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n951), .B1(new_n969), .B2(new_n983), .ZN(G387));
  NAND2_X1  g0784(.A1(new_n964), .A2(new_n734), .ZN(new_n985));
  INV_X1    g0785(.A(new_n681), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n745), .A2(new_n986), .B1(new_n234), .B2(new_n208), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n320), .A2(new_n251), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT50), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n262), .B1(new_n228), .B2(new_n202), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n989), .A2(new_n986), .A3(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n748), .B1(new_n243), .B2(new_n262), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n987), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n744), .B1(new_n993), .B2(new_n752), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n773), .A2(new_n387), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT109), .ZN(new_n996));
  AND2_X1   g0796(.A1(new_n776), .A2(new_n323), .ZN(new_n997));
  OAI22_X1  g0797(.A1(new_n764), .A2(new_n202), .B1(new_n759), .B2(new_n284), .ZN(new_n998));
  NOR4_X1   g0798(.A1(new_n997), .A2(new_n998), .A3(new_n394), .A4(new_n943), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G50), .A2(new_n767), .B1(new_n809), .B2(G68), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n996), .A2(new_n999), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1001), .B1(new_n406), .B2(new_n783), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G317), .A2(new_n767), .B1(new_n808), .B2(G322), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n762), .B2(new_n770), .C1(new_n782), .C2(new_n769), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT48), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n818), .A2(new_n556), .B1(new_n776), .B2(G283), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT49), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n394), .B1(new_n759), .B2(new_n771), .C1(new_n535), .C2(new_n756), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1010), .B2(KEYINPUT49), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1002), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n994), .B1(new_n673), .B2(new_n742), .C1(new_n1014), .C2(new_n797), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n965), .A2(new_n679), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n964), .A2(new_n729), .ZN(new_n1017));
  OAI211_X1 g0817(.A(new_n985), .B(new_n1015), .C1(new_n1016), .C2(new_n1017), .ZN(G393));
  OAI21_X1  g0818(.A(new_n752), .B1(new_n469), .B2(new_n207), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n250), .A2(new_n208), .A3(new_n268), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n735), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n775), .A2(new_n202), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n830), .A2(new_n394), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1023), .B1(new_n228), .B2(new_n764), .C1(new_n759), .C2(new_n811), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1022), .B(new_n1024), .C1(new_n320), .C2(new_n809), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n251), .B2(new_n782), .ZN(new_n1026));
  OAI22_X1  g0826(.A1(new_n284), .A2(new_n773), .B1(new_n766), .B2(new_n387), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT51), .Z(new_n1028));
  NOR2_X1   g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  OR2_X1    g0829(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1029), .A2(KEYINPUT110), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G311), .A2(new_n767), .B1(new_n808), .B2(G317), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT52), .Z(new_n1033));
  AOI22_X1  g0833(.A1(G283), .A2(new_n818), .B1(new_n760), .B2(G322), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n268), .B1(new_n757), .B2(G107), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1034), .B(new_n1035), .C1(new_n535), .C2(new_n775), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G294), .B2(new_n809), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1033), .B(new_n1037), .C1(new_n762), .C2(new_n782), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1030), .A2(new_n1031), .A3(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1021), .B1(new_n1039), .B2(new_n751), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1040), .B1(new_n742), .B2(new_n955), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n961), .B2(new_n733), .ZN(new_n1042));
  AND2_X1   g0842(.A1(new_n966), .A2(new_n679), .ZN(new_n1043));
  AND2_X1   g0843(.A1(new_n961), .A2(new_n965), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1044), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(G390));
  NAND3_X1  g0847(.A1(new_n873), .A2(new_n876), .A3(new_n739), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n836), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n735), .B1(new_n1049), .B2(new_n406), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n469), .A2(new_n770), .B1(new_n773), .B2(new_n823), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(G116), .B2(new_n767), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n756), .A2(new_n228), .B1(new_n759), .B2(new_n827), .ZN(new_n1053));
  NOR4_X1   g0853(.A1(new_n1053), .A2(new_n787), .A3(new_n1022), .A4(new_n268), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(new_n234), .C2(new_n782), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n764), .A2(new_n284), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(KEYINPUT115), .B(KEYINPUT53), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1056), .B(new_n1057), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(G159), .B2(new_n776), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT54), .B(G143), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT113), .Z(new_n1061));
  AOI22_X1  g0861(.A1(new_n1061), .A2(new_n809), .B1(new_n767), .B2(G132), .ZN(new_n1062));
  INV_X1    g0862(.A(G128), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1059), .B(new_n1062), .C1(new_n1063), .C2(new_n773), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n268), .B1(new_n756), .B2(new_n251), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(G125), .B2(new_n760), .ZN(new_n1066));
  XNOR2_X1  g0866(.A(new_n1066), .B(KEYINPUT114), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1067), .B1(new_n934), .B2(new_n782), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1055), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n1050), .B1(new_n1069), .B2(new_n751), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1048), .A2(new_n1070), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n903), .A2(G330), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n1073), .A2(new_n894), .A3(new_n803), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n881), .B1(new_n888), .B2(new_n894), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n873), .A2(new_n1076), .A3(new_n876), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n659), .B(new_n801), .C1(new_n717), .C2(new_n722), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n802), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n893), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n907), .A2(new_n1080), .A3(new_n881), .ZN(new_n1081));
  AOI211_X1 g0881(.A(KEYINPUT111), .B(new_n1075), .C1(new_n1077), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(KEYINPUT111), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n1081), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n1074), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n713), .A2(G330), .A3(new_n887), .A4(new_n893), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1077), .A2(new_n1086), .A3(new_n1081), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1082), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n894), .B1(new_n1073), .B2(new_n803), .ZN(new_n1089));
  NAND4_X1  g0889(.A1(new_n1086), .A2(new_n802), .A3(new_n1078), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n713), .A2(G330), .A3(new_n887), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1074), .B1(new_n1091), .B2(new_n894), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1090), .B1(new_n1092), .B2(new_n888), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n439), .A2(new_n1073), .ZN(new_n1094));
  NOR3_X1   g0894(.A1(new_n898), .A2(new_n621), .A3(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1093), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n680), .B1(new_n1088), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1084), .A2(new_n1074), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(KEYINPUT111), .A3(new_n1087), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n1084), .A2(new_n1083), .A3(new_n1074), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1096), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1072), .B1(new_n1097), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g0904(.A(KEYINPUT112), .B1(new_n1088), .B2(new_n733), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT112), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1101), .A2(new_n1106), .A3(new_n734), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1105), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1104), .A2(new_n1108), .ZN(G378));
  NAND2_X1  g0909(.A1(new_n297), .A2(new_n658), .ZN(new_n1110));
  XOR2_X1   g0910(.A(new_n1110), .B(KEYINPUT55), .Z(new_n1111));
  AND2_X1   g0911(.A1(new_n311), .A2(new_n1111), .ZN(new_n1112));
  NOR2_X1   g0912(.A1(new_n311), .A2(new_n1111), .ZN(new_n1113));
  NOR2_X1   g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  XOR2_X1   g0914(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1115), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1116), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n739), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n735), .B1(new_n1049), .B2(G50), .ZN(new_n1122));
  OAI22_X1  g0922(.A1(new_n234), .A2(new_n766), .B1(new_n773), .B2(new_n535), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1123), .B1(new_n323), .B2(new_n809), .ZN(new_n1124));
  OAI211_X1 g0924(.A(new_n261), .B(new_n394), .C1(new_n756), .C2(new_n383), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n764), .A2(new_n202), .B1(new_n759), .B2(new_n823), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(G68), .C2(new_n776), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1124), .B(new_n1127), .C1(new_n469), .C2(new_n782), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT58), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(G33), .A2(G41), .ZN(new_n1130));
  XNOR2_X1  g0930(.A(new_n1130), .B(KEYINPUT116), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G50), .B1(new_n394), .B2(new_n261), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n1128), .A2(new_n1129), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1131), .B1(G124), .B2(new_n760), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n1061), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1135), .A2(new_n764), .B1(new_n284), .B2(new_n775), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G125), .A2(new_n808), .B1(new_n767), .B2(G128), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1137), .B1(new_n934), .B2(new_n770), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1136), .B(new_n1138), .C1(G132), .C2(new_n783), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT59), .ZN(new_n1140));
  OAI221_X1 g0940(.A(new_n1134), .B1(new_n387), .B2(new_n756), .C1(new_n1139), .C2(new_n1140), .ZN(new_n1141));
  AND2_X1   g0941(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1133), .B1(new_n1129), .B2(new_n1128), .C1(new_n1141), .C2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1122), .B1(new_n1143), .B2(new_n751), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1121), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n870), .A2(new_n854), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n859), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n905), .B1(new_n1147), .B2(new_n857), .ZN(new_n1148));
  OAI21_X1  g0948(.A(G330), .B1(new_n1148), .B2(KEYINPUT40), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n907), .A2(new_n908), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT118), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT118), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n906), .A2(new_n909), .A3(new_n1152), .A4(G330), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1153), .A3(new_n1120), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1119), .A2(new_n906), .A3(G330), .A4(new_n909), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT119), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1154), .A2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n906), .A2(G330), .A3(new_n909), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1119), .B1(new_n1159), .B2(KEYINPUT118), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1160), .A2(new_n1156), .A3(new_n1153), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n897), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1158), .A2(new_n897), .A3(new_n1161), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1145), .B1(new_n1165), .B2(new_n733), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT120), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1096), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1095), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1167), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1170));
  OAI211_X1 g0970(.A(KEYINPUT120), .B(new_n1095), .C1(new_n1088), .C2(new_n1096), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AND3_X1   g0972(.A1(new_n1158), .A2(new_n897), .A3(new_n1161), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1173), .A2(new_n1162), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  NOR3_X1   g0977(.A1(new_n1173), .A2(new_n1162), .A3(new_n1176), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n680), .B1(new_n1178), .B2(new_n1172), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1166), .B1(new_n1177), .B2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(G375));
  INV_X1    g0981(.A(new_n1093), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n1169), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1183), .A2(new_n968), .A3(new_n1096), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n735), .B1(new_n1049), .B2(G68), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n893), .A2(new_n740), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n815), .A2(new_n773), .B1(new_n770), .B2(new_n284), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1187), .B1(G137), .B2(new_n767), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n268), .B1(new_n756), .B2(new_n383), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n764), .A2(new_n387), .B1(new_n759), .B2(new_n1063), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n1189), .B(new_n1190), .C1(G50), .C2(new_n776), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1188), .B(new_n1191), .C1(new_n782), .C2(new_n1135), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n782), .A2(new_n535), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n268), .B1(new_n757), .B2(G77), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1194), .A2(KEYINPUT122), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1195), .B1(G283), .B2(new_n767), .ZN(new_n1196));
  OAI22_X1  g0996(.A1(new_n764), .A2(new_n469), .B1(new_n759), .B2(new_n762), .ZN(new_n1197));
  AOI211_X1 g0997(.A(new_n1197), .B(new_n997), .C1(KEYINPUT122), .C2(new_n1194), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(G294), .A2(new_n808), .B1(new_n809), .B2(G107), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1196), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1192), .B1(new_n1193), .B2(new_n1200), .ZN(new_n1201));
  AOI211_X1 g1001(.A(new_n1185), .B(new_n1186), .C1(new_n751), .C2(new_n1201), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n733), .B(KEYINPUT121), .Z(new_n1203));
  AOI21_X1  g1003(.A(new_n1202), .B1(new_n1093), .B2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1184), .A2(new_n1204), .ZN(G381));
  NAND3_X1  g1005(.A1(new_n1099), .A2(new_n1100), .A3(new_n1096), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1103), .A2(new_n679), .A3(new_n1206), .ZN(new_n1207));
  AND4_X1   g1007(.A1(KEYINPUT124), .A2(new_n1108), .A3(new_n1207), .A4(new_n1071), .ZN(new_n1208));
  AOI21_X1  g1008(.A(KEYINPUT124), .B1(new_n1104), .B2(new_n1108), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(G375), .A2(new_n1211), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1213));
  XOR2_X1   g1013(.A(new_n1213), .B(KEYINPUT123), .Z(new_n1214));
  NOR3_X1   g1014(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(G407));
  NOR2_X1   g1016(.A1(new_n657), .A2(G343), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1212), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(G407), .A2(new_n1218), .A3(G213), .ZN(G409));
  INV_X1    g1019(.A(new_n1217), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1203), .B1(new_n1172), .B2(new_n968), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1145), .B1(new_n1221), .B2(new_n1165), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1180), .A2(G378), .B1(new_n1222), .B2(new_n1210), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1220), .B1(new_n1223), .B2(KEYINPUT125), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1222), .A2(new_n1210), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n1174), .A2(new_n734), .B1(new_n1121), .B2(new_n1144), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1163), .A2(KEYINPUT57), .A3(new_n1164), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n679), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(KEYINPUT57), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1230));
  OAI211_X1 g1030(.A(G378), .B(new_n1226), .C1(new_n1229), .C2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1225), .A2(new_n1231), .A3(KEYINPUT125), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(KEYINPUT127), .B1(new_n1224), .B2(new_n1233), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n807), .A2(KEYINPUT126), .A3(new_n840), .ZN(new_n1235));
  AND2_X1   g1035(.A1(new_n1235), .A2(new_n1204), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1096), .A2(KEYINPUT60), .ZN(new_n1237));
  AND2_X1   g1037(.A1(new_n1237), .A2(new_n1183), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n679), .B1(new_n1237), .B2(new_n1183), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1236), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT126), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n1241), .A3(G384), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(G384), .A2(new_n1241), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1236), .B(new_n1243), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1217), .A2(G2897), .ZN(new_n1246));
  XOR2_X1   g1046(.A(new_n1245), .B(new_n1246), .Z(new_n1247));
  NAND2_X1  g1047(.A1(new_n1225), .A2(new_n1231), .ZN(new_n1248));
  INV_X1    g1048(.A(KEYINPUT125), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT127), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1250), .A2(new_n1251), .A3(new_n1220), .A4(new_n1232), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1234), .A2(new_n1247), .A3(new_n1252), .ZN(new_n1253));
  NAND4_X1  g1053(.A1(new_n1248), .A2(KEYINPUT63), .A3(new_n1220), .A4(new_n1245), .ZN(new_n1254));
  OR2_X1    g1054(.A1(G387), .A2(new_n1046), .ZN(new_n1255));
  XOR2_X1   g1055(.A(G393), .B(G396), .Z(new_n1256));
  NAND2_X1  g1056(.A1(G387), .A2(new_n1046), .ZN(new_n1257));
  AND3_X1   g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1256), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1258), .A2(new_n1259), .A3(KEYINPUT61), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1254), .A2(new_n1260), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT63), .ZN(new_n1262));
  NAND4_X1  g1062(.A1(new_n1250), .A2(new_n1220), .A3(new_n1245), .A4(new_n1232), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1261), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1253), .A2(new_n1264), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1263), .A2(KEYINPUT62), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1247), .B1(new_n1223), .B2(new_n1217), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1245), .ZN(new_n1271));
  AOI211_X1 g1071(.A(new_n1217), .B(new_n1271), .C1(new_n1225), .C2(new_n1231), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT62), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1269), .B(new_n1270), .C1(new_n1272), .C2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1267), .B1(new_n1268), .B2(new_n1274), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1265), .A2(new_n1275), .ZN(G405));
  OAI21_X1  g1076(.A(new_n1231), .B1(new_n1211), .B2(new_n1180), .ZN(new_n1277));
  XNOR2_X1  g1077(.A(new_n1266), .B(new_n1277), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(new_n1278), .B(new_n1271), .ZN(G402));
endmodule


