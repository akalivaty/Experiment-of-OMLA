//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1224, new_n1225,
    new_n1226, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1279, new_n1280, new_n1281,
    new_n1282, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G58), .ZN(new_n205));
  INV_X1    g0005(.A(G232), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT67), .Z(new_n209));
  NAND2_X1  g0009(.A1(G116), .A2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  XOR2_X1   g0011(.A(KEYINPUT65), .B(G77), .Z(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(G244), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n210), .B(new_n211), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  AOI211_X1 g0015(.A(new_n207), .B(new_n209), .C1(new_n215), .C2(KEYINPUT66), .ZN(new_n216));
  INV_X1    g0016(.A(G107), .ZN(new_n217));
  INV_X1    g0017(.A(G264), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n216), .B1(KEYINPUT66), .B2(new_n215), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G20), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT64), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND2_X1  g0026(.A1(G1), .A2(G13), .ZN(new_n227));
  INV_X1    g0027(.A(new_n227), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(G50), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n223), .B(new_n226), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G250), .B(G257), .Z(new_n237));
  XNOR2_X1  g0037(.A(G264), .B(G270), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT68), .B(G107), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G68), .B(G77), .Z(new_n245));
  XNOR2_X1  g0045(.A(G50), .B(G58), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT70), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  OAI21_X1  g0050(.A(new_n249), .B1(new_n220), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g0051(.A1(KEYINPUT70), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n251), .A2(new_n227), .A3(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT76), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT3), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(G33), .A3(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g0061(.A(G20), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G87), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT22), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT22), .A2(G20), .ZN(new_n265));
  AND2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  OAI211_X1 g0066(.A(G87), .B(new_n265), .C1(new_n266), .C2(new_n260), .ZN(new_n267));
  XOR2_X1   g0067(.A(new_n267), .B(KEYINPUT87), .Z(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT24), .ZN(new_n270));
  INV_X1    g0070(.A(G20), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n271), .A2(G33), .A3(G116), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n217), .A2(G20), .ZN(new_n273));
  XOR2_X1   g0073(.A(new_n273), .B(KEYINPUT23), .Z(new_n274));
  NAND4_X1  g0074(.A1(new_n269), .A2(new_n270), .A3(new_n272), .A4(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT22), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n262), .B2(G87), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n267), .B(KEYINPUT87), .ZN(new_n278));
  OAI211_X1 g0078(.A(new_n272), .B(new_n274), .C1(new_n277), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(KEYINPUT24), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n254), .B1(new_n275), .B2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G13), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n282), .A2(G1), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G20), .A3(new_n217), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(KEYINPUT25), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NOR3_X1   g0086(.A1(new_n282), .A2(new_n271), .A3(G1), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n250), .A2(G1), .ZN(new_n288));
  NOR3_X1   g0088(.A1(new_n253), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  OAI22_X1  g0090(.A1(new_n290), .A2(new_n217), .B1(KEYINPUT25), .B2(new_n284), .ZN(new_n291));
  OR3_X1    g0091(.A1(new_n281), .A2(new_n286), .A3(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n259), .A2(new_n261), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  OR2_X1    g0094(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n295));
  NAND2_X1  g0095(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AOI22_X1  g0097(.A1(new_n297), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n298));
  INV_X1    g0098(.A(G294), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n294), .A2(new_n298), .B1(new_n250), .B2(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n227), .B1(G33), .B2(G41), .ZN(new_n301));
  INV_X1    g0101(.A(G45), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  AND2_X1   g0103(.A1(KEYINPUT5), .A2(G41), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT5), .A2(G41), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G41), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n228), .B1(new_n250), .B2(new_n307), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n300), .A2(new_n301), .B1(G264), .B2(new_n309), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n303), .B(G274), .C1(new_n305), .C2(new_n304), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G169), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n310), .A2(G179), .A3(new_n311), .ZN(new_n314));
  AND2_X1   g0114(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT88), .ZN(new_n316));
  AOI21_X1  g0116(.A(KEYINPUT88), .B1(new_n313), .B2(new_n314), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n292), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(G58), .A2(G68), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n271), .B1(new_n202), .B2(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n271), .A2(new_n250), .A3(KEYINPUT71), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT71), .B1(new_n271), .B2(new_n250), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n321), .B1(new_n325), .B2(G159), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT79), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n256), .B2(G33), .ZN(new_n328));
  NOR3_X1   g0128(.A1(new_n250), .A2(KEYINPUT79), .A3(KEYINPUT3), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n257), .A2(new_n250), .A3(new_n258), .ZN(new_n331));
  AOI21_X1  g0131(.A(G20), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NOR3_X1   g0132(.A1(new_n266), .A2(new_n260), .A3(G20), .ZN(new_n333));
  OAI21_X1  g0133(.A(KEYINPUT78), .B1(new_n333), .B2(KEYINPUT7), .ZN(new_n334));
  NAND2_X1  g0134(.A1(KEYINPUT3), .A2(G33), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n261), .A2(new_n271), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT78), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT7), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  AOI22_X1  g0139(.A1(new_n332), .A2(KEYINPUT7), .B1(new_n334), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G68), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n326), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT16), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g0144(.A(KEYINPUT7), .B1(new_n293), .B2(G20), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n259), .A2(new_n338), .A3(new_n271), .A4(new_n261), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(G68), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n326), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT77), .B1(new_n348), .B2(new_n343), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT77), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n347), .A2(new_n350), .A3(KEYINPUT16), .A4(new_n326), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n344), .A2(new_n349), .A3(new_n253), .A4(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G1), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(G41), .B2(G45), .ZN(new_n354));
  INV_X1    g0154(.A(G274), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(new_n308), .A2(new_n354), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(G232), .ZN(new_n359));
  AND2_X1   g0159(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n360));
  NOR2_X1   g0160(.A1(KEYINPUT69), .A2(G1698), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(G223), .ZN(new_n363));
  INV_X1    g0163(.A(G226), .ZN(new_n364));
  INV_X1    g0164(.A(G1698), .ZN(new_n365));
  OAI22_X1  g0165(.A1(new_n362), .A2(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(new_n293), .B1(G33), .B2(G87), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n357), .B(new_n359), .C1(new_n367), .C2(new_n308), .ZN(new_n368));
  INV_X1    g0168(.A(G190), .ZN(new_n369));
  OR2_X1    g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n287), .ZN(new_n371));
  XNOR2_X1  g0171(.A(KEYINPUT8), .B(G58), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n253), .B1(new_n353), .B2(G20), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n373), .B1(new_n374), .B2(new_n372), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n368), .A2(G200), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n352), .A2(new_n370), .A3(new_n375), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(KEYINPUT17), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT17), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n352), .A2(new_n375), .ZN(new_n382));
  INV_X1    g0182(.A(new_n368), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT80), .ZN(new_n384));
  INV_X1    g0184(.A(G179), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g0186(.A(KEYINPUT80), .B1(new_n368), .B2(G179), .ZN(new_n387));
  INV_X1    g0187(.A(G169), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n368), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n386), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n382), .A2(new_n391), .A3(KEYINPUT18), .ZN(new_n392));
  INV_X1    g0192(.A(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(KEYINPUT18), .B1(new_n382), .B2(new_n391), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n379), .B(new_n381), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n266), .A2(new_n260), .ZN(new_n398));
  INV_X1    g0198(.A(new_n398), .ZN(new_n399));
  INV_X1    g0199(.A(G238), .ZN(new_n400));
  OAI221_X1 g0200(.A(new_n399), .B1(new_n400), .B2(new_n365), .C1(new_n362), .C2(new_n206), .ZN(new_n401));
  OAI211_X1 g0201(.A(new_n401), .B(new_n301), .C1(G107), .C2(new_n399), .ZN(new_n402));
  INV_X1    g0202(.A(new_n358), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n357), .C1(new_n214), .C2(new_n403), .ZN(new_n404));
  OR2_X1    g0204(.A1(new_n404), .A2(new_n369), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(G200), .ZN(new_n406));
  XOR2_X1   g0206(.A(KEYINPUT15), .B(G87), .Z(new_n407));
  NAND3_X1  g0207(.A1(new_n407), .A2(new_n271), .A3(G33), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n408), .B1(new_n324), .B2(new_n372), .C1(new_n271), .C2(new_n213), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(new_n253), .B1(G77), .B2(new_n374), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n213), .A2(new_n287), .ZN(new_n411));
  XNOR2_X1  g0211(.A(new_n411), .B(KEYINPUT72), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT73), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(KEYINPUT73), .A3(new_n412), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n405), .A2(new_n406), .A3(new_n415), .A4(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n297), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n398), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G97), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(KEYINPUT74), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT74), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n422), .A2(G33), .A3(G97), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n301), .B1(new_n419), .B2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT13), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n358), .A2(G238), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n357), .ZN(new_n428));
  OAI22_X1  g0228(.A1(new_n362), .A2(new_n364), .B1(new_n206), .B2(new_n365), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n424), .B1(new_n429), .B2(new_n399), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n427), .B(new_n357), .C1(new_n430), .C2(new_n308), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT13), .ZN(new_n432));
  AND2_X1   g0232(.A1(new_n428), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n433), .A2(G190), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n271), .A2(G33), .A3(G77), .ZN(new_n435));
  INV_X1    g0235(.A(G50), .ZN(new_n436));
  OAI221_X1 g0236(.A(new_n435), .B1(new_n271), .B2(G68), .C1(new_n324), .C2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n253), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT11), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n437), .A2(KEYINPUT11), .A3(new_n253), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n374), .A2(G68), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n283), .A2(G20), .A3(new_n341), .ZN(new_n443));
  XNOR2_X1  g0243(.A(new_n443), .B(KEYINPUT12), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n440), .A2(new_n441), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n428), .A2(new_n432), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(G200), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n434), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  OR2_X1    g0249(.A1(new_n404), .A2(G179), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n404), .A2(new_n388), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n450), .A2(new_n413), .A3(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n397), .A2(new_n417), .A3(new_n449), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n374), .A2(G50), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n271), .B1(new_n201), .B2(new_n436), .ZN(new_n455));
  NOR3_X1   g0255(.A1(new_n372), .A2(G20), .A3(new_n250), .ZN(new_n456));
  AOI211_X1 g0256(.A(new_n455), .B(new_n456), .C1(G150), .C2(new_n325), .ZN(new_n457));
  OAI221_X1 g0257(.A(new_n454), .B1(G50), .B2(new_n371), .C1(new_n457), .C2(new_n254), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT9), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n398), .B1(G222), .B2(new_n297), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n363), .B2(new_n365), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n301), .C1(new_n212), .C2(new_n399), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n463), .B(new_n357), .C1(new_n364), .C2(new_n403), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G200), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n458), .A2(new_n459), .ZN(new_n466));
  OR2_X1    g0266(.A1(new_n464), .A2(new_n369), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n460), .A2(new_n465), .A3(new_n466), .A4(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT10), .ZN(new_n469));
  OR2_X1    g0269(.A1(new_n464), .A2(G179), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n464), .A2(new_n388), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(new_n458), .A3(new_n471), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n445), .A2(KEYINPUT75), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n445), .A2(KEYINPUT75), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT14), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n447), .B2(G169), .ZN(new_n477));
  AOI211_X1 g0277(.A(KEYINPUT14), .B(new_n388), .C1(new_n428), .C2(new_n432), .ZN(new_n478));
  NOR2_X1   g0278(.A1(new_n447), .A2(new_n385), .ZN(new_n479));
  NOR3_X1   g0279(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n469), .B(new_n472), .C1(new_n475), .C2(new_n480), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n396), .A2(KEYINPUT81), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n453), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(G257), .ZN(new_n484));
  OAI22_X1  g0284(.A1(new_n362), .A2(new_n484), .B1(new_n218), .B2(new_n365), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(new_n293), .B1(G303), .B2(new_n398), .ZN(new_n486));
  NOR2_X1   g0286(.A1(new_n486), .A2(new_n308), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n487), .B1(G270), .B2(new_n309), .ZN(new_n488));
  INV_X1    g0288(.A(G116), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n489), .A2(G20), .ZN(new_n490));
  NAND2_X1  g0290(.A1(G33), .A2(G283), .ZN(new_n491));
  INV_X1    g0291(.A(G97), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n491), .B(new_n271), .C1(G33), .C2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n253), .A2(new_n490), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT20), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n253), .A2(KEYINPUT20), .A3(new_n490), .A4(new_n493), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n496), .A2(new_n497), .B1(G116), .B2(new_n289), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n287), .A2(new_n489), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n488), .A2(G179), .A3(new_n311), .A4(new_n500), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n498), .A2(new_n499), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n309), .A2(G270), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n311), .B(new_n503), .C1(new_n486), .C2(new_n308), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(G200), .ZN(new_n505));
  OAI211_X1 g0305(.A(new_n502), .B(new_n505), .C1(new_n369), .C2(new_n504), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n388), .B1(new_n498), .B2(new_n499), .ZN(new_n507));
  INV_X1    g0307(.A(KEYINPUT21), .ZN(new_n508));
  AND3_X1   g0308(.A1(new_n507), .A2(new_n508), .A3(new_n504), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n507), .B2(new_n504), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n501), .B(new_n506), .C1(new_n509), .C2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n289), .A2(new_n407), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n293), .A2(new_n271), .A3(G68), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT19), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n420), .A2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(G87), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n516), .A2(new_n492), .A3(new_n217), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n421), .B2(new_n423), .ZN(new_n518));
  OAI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G20), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n513), .A2(new_n515), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n520), .A2(new_n253), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n371), .A2(new_n407), .ZN(new_n522));
  INV_X1    g0322(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(KEYINPUT86), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT86), .ZN(new_n525));
  AOI211_X1 g0325(.A(new_n525), .B(new_n522), .C1(new_n520), .C2(new_n253), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n512), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n301), .B1(new_n250), .B2(new_n489), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G244), .A2(G1698), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n362), .B2(new_n400), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n528), .B1(new_n530), .B2(new_n293), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n353), .A2(G45), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(G250), .ZN(new_n534));
  AOI21_X1  g0334(.A(G274), .B1(KEYINPUT84), .B2(G250), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n308), .B(new_n534), .C1(new_n532), .C2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(G179), .B1(new_n531), .B2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT85), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n297), .A2(G238), .ZN(new_n540));
  AOI22_X1  g0340(.A1(new_n540), .A2(new_n529), .B1(new_n261), .B2(new_n259), .ZN(new_n541));
  OAI211_X1 g0341(.A(G169), .B(new_n536), .C1(new_n541), .C2(new_n528), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n538), .A2(new_n539), .A3(new_n542), .ZN(new_n543));
  AOI21_X1  g0343(.A(new_n539), .B1(new_n538), .B2(new_n542), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n527), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n536), .B1(new_n541), .B2(new_n528), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(G190), .ZN(new_n548));
  OAI211_X1 g0348(.A(G200), .B(new_n536), .C1(new_n541), .C2(new_n528), .ZN(new_n549));
  AND2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g0350(.A1(new_n290), .A2(new_n516), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n550), .B(new_n552), .C1(new_n524), .C2(new_n526), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n546), .A2(new_n553), .ZN(new_n554));
  NOR2_X1   g0354(.A1(new_n511), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n325), .A2(G77), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n217), .A2(KEYINPUT6), .A3(G97), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n492), .A2(new_n217), .ZN(new_n558));
  NOR2_X1   g0358(.A1(G97), .A2(G107), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n560), .B2(KEYINPUT6), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n561), .A2(G20), .ZN(new_n562));
  OAI211_X1 g0362(.A(new_n556), .B(new_n562), .C1(new_n340), .C2(new_n217), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n563), .A2(new_n253), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n371), .A2(G97), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n289), .B2(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(new_n214), .B1(new_n295), .B2(new_n296), .ZN(new_n568));
  AND2_X1   g0368(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n569));
  NOR2_X1   g0369(.A1(KEYINPUT76), .A2(KEYINPUT3), .ZN(new_n570));
  NOR3_X1   g0370(.A1(new_n569), .A2(new_n570), .A3(new_n250), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n568), .B1(new_n571), .B2(new_n260), .ZN(new_n572));
  XOR2_X1   g0372(.A(KEYINPUT82), .B(KEYINPUT4), .Z(new_n573));
  OAI211_X1 g0373(.A(KEYINPUT4), .B(G244), .C1(new_n360), .C2(new_n361), .ZN(new_n574));
  NAND2_X1  g0374(.A1(G250), .A2(G1698), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  AOI22_X1  g0376(.A1(new_n572), .A2(new_n573), .B1(new_n576), .B2(new_n399), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n308), .B1(new_n577), .B2(new_n491), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n306), .A2(new_n308), .A3(G257), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n311), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT83), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT83), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n582), .A3(new_n311), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(G169), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n576), .A2(new_n399), .ZN(new_n586));
  OAI21_X1  g0386(.A(G244), .B1(new_n360), .B2(new_n361), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n261), .B2(new_n259), .ZN(new_n588));
  INV_X1    g0388(.A(new_n573), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n586), .B(new_n491), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n301), .ZN(new_n591));
  INV_X1    g0391(.A(new_n583), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n582), .B1(new_n579), .B2(new_n311), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n591), .A2(new_n594), .A3(G179), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n585), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n567), .A2(new_n596), .ZN(new_n597));
  INV_X1    g0397(.A(new_n566), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n598), .B1(new_n563), .B2(new_n253), .ZN(new_n599));
  OAI21_X1  g0399(.A(G200), .B1(new_n578), .B2(new_n584), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n591), .A2(new_n594), .A3(G190), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n312), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(G190), .ZN(new_n605));
  INV_X1    g0405(.A(G200), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n606), .B1(new_n310), .B2(new_n311), .ZN(new_n607));
  NOR4_X1   g0407(.A1(new_n281), .A2(new_n286), .A3(new_n291), .A4(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n603), .B1(new_n605), .B2(new_n608), .ZN(new_n609));
  AND4_X1   g0409(.A1(new_n319), .A2(new_n483), .A3(new_n555), .A4(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n472), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n382), .A2(new_n391), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT18), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n392), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n379), .A2(new_n381), .ZN(new_n616));
  INV_X1    g0416(.A(new_n477), .ZN(new_n617));
  INV_X1    g0417(.A(new_n479), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n447), .A2(new_n476), .A3(G169), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n473), .A2(new_n474), .ZN(new_n621));
  INV_X1    g0421(.A(new_n452), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(new_n449), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n615), .B1(new_n616), .B2(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n611), .B1(new_n624), .B2(new_n469), .ZN(new_n625));
  INV_X1    g0425(.A(new_n483), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n521), .A2(new_n523), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n525), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n521), .A2(KEYINPUT86), .A3(new_n523), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n551), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n548), .A2(KEYINPUT89), .A3(new_n549), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n631), .B1(KEYINPUT89), .B2(new_n549), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n538), .A2(new_n542), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n630), .A2(new_n632), .B1(new_n527), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n501), .B1(new_n509), .B2(new_n510), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n281), .A2(new_n286), .A3(new_n291), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n636), .A2(new_n315), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n609), .B(new_n634), .C1(new_n635), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n527), .A2(new_n633), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  AOI22_X1  g0440(.A1(new_n564), .A2(new_n566), .B1(new_n585), .B2(new_n595), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n546), .A2(new_n641), .A3(new_n553), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n640), .B1(new_n642), .B2(KEYINPUT26), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n585), .A2(new_n595), .ZN(new_n644));
  OAI21_X1  g0444(.A(KEYINPUT90), .B1(new_n644), .B2(new_n599), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT26), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT90), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n567), .A2(new_n596), .A3(new_n647), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n634), .A2(new_n645), .A3(new_n646), .A4(new_n648), .ZN(new_n649));
  AND3_X1   g0449(.A1(new_n643), .A2(KEYINPUT91), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(KEYINPUT91), .B1(new_n643), .B2(new_n649), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n638), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n625), .B1(new_n626), .B2(new_n653), .ZN(G369));
  NOR2_X1   g0454(.A1(new_n282), .A2(G20), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n353), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n659), .A2(G343), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT93), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n637), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n660), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n292), .A2(KEYINPUT92), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n608), .A2(new_n605), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT92), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n667), .B1(new_n636), .B2(new_n660), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n665), .A2(new_n319), .A3(new_n666), .A4(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n635), .A2(new_n660), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n663), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT94), .ZN(new_n672));
  INV_X1    g0472(.A(KEYINPUT94), .ZN(new_n673));
  OAI211_X1 g0473(.A(new_n673), .B(new_n663), .C1(new_n669), .C2(new_n670), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n319), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(new_n664), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n669), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n502), .A2(new_n660), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n635), .A2(new_n679), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n511), .B2(new_n679), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n681), .A2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n675), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g0485(.A(new_n685), .B(KEYINPUT95), .Z(G399));
  INV_X1    g0486(.A(new_n224), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n687), .A2(G41), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n517), .A2(G116), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G1), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n230), .B2(new_n689), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT96), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n609), .A2(new_n319), .A3(new_n555), .A4(new_n662), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n578), .A2(new_n584), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n488), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n310), .A2(G179), .A3(new_n311), .A4(new_n547), .ZN(new_n699));
  NOR3_X1   g0499(.A1(new_n698), .A2(KEYINPUT30), .A3(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT30), .B1(new_n698), .B2(new_n699), .ZN(new_n702));
  INV_X1    g0502(.A(new_n547), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n504), .A2(new_n703), .A3(new_n385), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT97), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n697), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n604), .B1(new_n705), .B2(new_n704), .ZN(new_n708));
  AOI22_X1  g0508(.A1(new_n701), .A2(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n696), .B1(new_n709), .B2(new_n660), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n708), .ZN(new_n711));
  INV_X1    g0511(.A(new_n702), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n700), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n661), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n695), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G330), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(KEYINPUT98), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT98), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n715), .A2(new_n718), .A3(G330), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT29), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n634), .A2(new_n645), .A3(new_n648), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(KEYINPUT26), .ZN(new_n723));
  OR2_X1    g0523(.A1(new_n642), .A2(KEYINPUT26), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(new_n639), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(KEYINPUT99), .ZN(new_n726));
  OAI211_X1 g0526(.A(new_n609), .B(new_n634), .C1(new_n676), .C2(new_n635), .ZN(new_n727));
  INV_X1    g0527(.A(KEYINPUT99), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n723), .A2(new_n724), .A3(new_n728), .A4(new_n639), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n726), .A2(new_n727), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g0530(.A(new_n721), .B1(new_n730), .B2(new_n660), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n652), .A2(new_n662), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  NOR3_X1   g0533(.A1(new_n720), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n694), .B1(new_n734), .B2(G1), .ZN(G364));
  NOR2_X1   g0535(.A1(new_n687), .A2(new_n293), .ZN(new_n736));
  XOR2_X1   g0536(.A(new_n736), .B(KEYINPUT101), .Z(new_n737));
  NAND3_X1  g0537(.A1(new_n202), .A2(new_n302), .A3(G50), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n737), .B(new_n738), .C1(new_n302), .C2(new_n247), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n224), .A2(G355), .A3(new_n399), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n739), .B(new_n740), .C1(G116), .C2(new_n224), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G13), .A2(G33), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT102), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(G20), .ZN(new_n745));
  AND2_X1   g0545(.A1(KEYINPUT103), .A2(G169), .ZN(new_n746));
  NOR2_X1   g0546(.A1(KEYINPUT103), .A2(G169), .ZN(new_n747));
  NOR3_X1   g0547(.A1(new_n746), .A2(new_n747), .A3(new_n271), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n227), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n745), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n741), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n655), .A2(G45), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT100), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n753), .A2(G1), .A3(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n688), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n271), .A2(new_n369), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n606), .A2(G179), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G303), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n398), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND3_X1  g0562(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(G317), .ZN(new_n765));
  OR2_X1    g0565(.A1(new_n765), .A2(KEYINPUT33), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(KEYINPUT33), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n764), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n763), .A2(new_n369), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G326), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n271), .B1(new_n771), .B2(G190), .ZN(new_n772));
  OAI211_X1 g0572(.A(new_n768), .B(new_n770), .C1(new_n299), .C2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n385), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n758), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n762), .B(new_n773), .C1(G322), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n271), .A2(G190), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n778), .A2(new_n759), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n778), .A2(new_n771), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G283), .A2(new_n780), .B1(new_n782), .B2(G329), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n783), .B(KEYINPUT105), .ZN(new_n784));
  INV_X1    g0584(.A(G311), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n778), .A2(new_n774), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n777), .B(new_n784), .C1(new_n785), .C2(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n782), .A2(G159), .ZN(new_n788));
  XNOR2_X1  g0588(.A(new_n788), .B(KEYINPUT104), .ZN(new_n789));
  XOR2_X1   g0589(.A(new_n789), .B(KEYINPUT32), .Z(new_n790));
  INV_X1    g0590(.A(new_n769), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n791), .A2(new_n436), .B1(new_n772), .B2(new_n492), .ZN(new_n792));
  INV_X1    g0592(.A(new_n764), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n399), .B1(new_n793), .B2(new_n341), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n760), .A2(new_n516), .ZN(new_n795));
  NOR3_X1   g0595(.A1(new_n792), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  AOI22_X1  g0596(.A1(G58), .A2(new_n776), .B1(new_n780), .B2(G107), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n796), .B(new_n797), .C1(new_n213), .C2(new_n786), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n787), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n757), .B1(new_n799), .B2(new_n749), .ZN(new_n800));
  INV_X1    g0600(.A(new_n745), .ZN(new_n801));
  OAI211_X1 g0601(.A(new_n751), .B(new_n800), .C1(new_n681), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n682), .A2(new_n757), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n681), .A2(G330), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n802), .B1(new_n803), .B2(new_n804), .ZN(G396));
  NAND2_X1  g0605(.A1(new_n413), .A2(new_n664), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n417), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(new_n452), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n622), .A2(new_n660), .ZN(new_n809));
  AND2_X1   g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n720), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n810), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(new_n717), .B2(new_n719), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  XNOR2_X1  g0614(.A(new_n814), .B(new_n732), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n757), .ZN(new_n816));
  AOI22_X1  g0616(.A1(new_n776), .A2(G143), .B1(G150), .B2(new_n764), .ZN(new_n817));
  INV_X1    g0617(.A(G137), .ZN(new_n818));
  INV_X1    g0618(.A(G159), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n791), .C1(new_n819), .C2(new_n786), .ZN(new_n820));
  INV_X1    g0620(.A(KEYINPUT34), .ZN(new_n821));
  OR2_X1    g0621(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n780), .A2(G68), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n820), .A2(new_n821), .ZN(new_n824));
  INV_X1    g0624(.A(G132), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n760), .A2(new_n436), .B1(new_n781), .B2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n772), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n294), .B(new_n826), .C1(G58), .C2(new_n827), .ZN(new_n828));
  NAND4_X1  g0628(.A1(new_n822), .A2(new_n823), .A3(new_n824), .A4(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(G283), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n793), .A2(new_n830), .B1(new_n791), .B2(new_n761), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G97), .B2(new_n827), .ZN(new_n832));
  INV_X1    g0632(.A(new_n786), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(G116), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n775), .A2(new_n299), .B1(new_n779), .B2(new_n516), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n835), .B1(G311), .B2(new_n782), .ZN(new_n836));
  INV_X1    g0636(.A(new_n760), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n399), .B1(new_n837), .B2(G107), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n832), .A2(new_n834), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n227), .B(new_n748), .C1(new_n829), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(G77), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n749), .A2(new_n742), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n757), .B(new_n840), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n843), .B(KEYINPUT106), .ZN(new_n844));
  OAI21_X1  g0644(.A(new_n844), .B1(new_n744), .B2(new_n810), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n816), .A2(new_n845), .ZN(G384));
  NAND2_X1  g0646(.A1(new_n348), .A2(new_n343), .ZN(new_n847));
  NAND4_X1  g0647(.A1(new_n349), .A2(new_n847), .A3(new_n253), .A4(new_n351), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n848), .A2(new_n375), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(new_n659), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n395), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n659), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n390), .A2(new_n853), .B1(new_n352), .B2(new_n375), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n378), .A2(new_n854), .ZN(new_n855));
  XNOR2_X1  g0655(.A(KEYINPUT109), .B(KEYINPUT37), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n391), .A2(new_n849), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n859), .A2(new_n850), .A3(new_n377), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(KEYINPUT37), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n377), .B(KEYINPUT17), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n850), .B1(new_n865), .B2(new_n615), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n855), .A2(new_n857), .B1(new_n860), .B2(KEYINPUT37), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n863), .A2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n449), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n660), .B1(new_n473), .B2(new_n474), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NOR3_X1   g0672(.A1(new_n480), .A2(new_n475), .A3(KEYINPUT108), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT108), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n874), .B1(new_n620), .B2(new_n621), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n872), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n871), .B1(new_n870), .B2(new_n620), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n652), .A2(new_n662), .A3(new_n808), .ZN(new_n879));
  INV_X1    g0679(.A(KEYINPUT107), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n879), .A2(new_n880), .A3(new_n809), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n879), .B2(new_n809), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n869), .B(new_n878), .C1(new_n881), .C2(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n853), .B1(new_n352), .B2(new_n375), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n395), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT111), .B1(new_n378), .B2(new_n854), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n382), .B1(new_n391), .B2(new_n659), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT111), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(new_n888), .A3(new_n377), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n856), .B1(new_n854), .B2(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n886), .A3(new_n889), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n885), .A2(new_n892), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n864), .ZN(new_n896));
  XOR2_X1   g0696(.A(KEYINPUT112), .B(KEYINPUT39), .Z(new_n897));
  NAND3_X1  g0697(.A1(new_n896), .A2(new_n863), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n869), .A2(KEYINPUT39), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n873), .A2(new_n875), .A3(new_n664), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n614), .A2(new_n392), .A3(new_n853), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n883), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n483), .B1(new_n731), .B2(new_n733), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(new_n625), .ZN(new_n906));
  XOR2_X1   g0706(.A(new_n904), .B(new_n906), .Z(new_n907));
  NAND3_X1  g0707(.A1(new_n713), .A2(KEYINPUT31), .A3(new_n664), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n695), .A2(new_n710), .A3(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n449), .B1(new_n475), .B2(new_n660), .ZN(new_n911));
  OAI21_X1  g0711(.A(KEYINPUT108), .B1(new_n480), .B2(new_n475), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n620), .A2(new_n621), .A3(new_n874), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g0714(.A(new_n877), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n810), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT113), .B1(new_n910), .B2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT113), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n878), .A2(new_n909), .A3(new_n918), .A4(new_n810), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n917), .A2(new_n869), .A3(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT40), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n910), .A2(new_n916), .ZN(new_n923));
  INV_X1    g0723(.A(new_n896), .ZN(new_n924));
  INV_X1    g0724(.A(new_n863), .ZN(new_n925));
  OAI211_X1 g0725(.A(KEYINPUT40), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n483), .A2(new_n909), .ZN(new_n928));
  XOR2_X1   g0728(.A(new_n927), .B(new_n928), .Z(new_n929));
  NAND2_X1  g0729(.A1(new_n929), .A2(G330), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n907), .B(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n353), .B2(new_n655), .ZN(new_n932));
  OAI211_X1 g0732(.A(G20), .B(new_n228), .C1(new_n561), .C2(KEYINPUT35), .ZN(new_n933));
  AOI211_X1 g0733(.A(new_n489), .B(new_n933), .C1(KEYINPUT35), .C2(new_n561), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT36), .Z(new_n935));
  NAND2_X1  g0735(.A1(new_n212), .A2(new_n320), .ZN(new_n936));
  OAI22_X1  g0736(.A1(new_n936), .A2(new_n230), .B1(G50), .B2(new_n341), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n937), .A2(G1), .A3(new_n282), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n932), .A2(new_n935), .A3(new_n938), .ZN(G367));
  NOR2_X1   g0739(.A1(new_n630), .A2(new_n660), .ZN(new_n940));
  MUX2_X1   g0740(.A(new_n634), .B(new_n640), .S(new_n940), .Z(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  OR2_X1    g0742(.A1(new_n669), .A2(new_n670), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n641), .A2(new_n661), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT114), .ZN(new_n945));
  OAI211_X1 g0745(.A(new_n597), .B(new_n602), .C1(new_n599), .C2(new_n662), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n949), .B(KEYINPUT42), .Z(new_n950));
  AOI21_X1  g0750(.A(new_n641), .B1(new_n947), .B2(new_n676), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT115), .ZN(new_n952));
  AND2_X1   g0752(.A1(new_n952), .A2(new_n662), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n942), .B1(new_n950), .B2(new_n953), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n684), .A2(new_n948), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  OAI221_X1 g0756(.A(new_n942), .B1(new_n684), .B2(new_n948), .C1(new_n950), .C2(new_n953), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n958));
  AND3_X1   g0758(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n958), .B1(new_n956), .B2(new_n957), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n688), .B(KEYINPUT41), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n684), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n948), .B1(new_n672), .B2(new_n674), .ZN(new_n965));
  OR2_X1    g0765(.A1(new_n965), .A2(KEYINPUT45), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n675), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n672), .A2(new_n674), .A3(new_n948), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n969), .A2(KEYINPUT44), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(KEYINPUT44), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n964), .B1(new_n968), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n966), .A2(new_n967), .ZN(new_n974));
  NAND4_X1  g0774(.A1(new_n974), .A2(new_n684), .A3(new_n971), .A4(new_n970), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n677), .A2(new_n669), .A3(new_n670), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n943), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(new_n683), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n734), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n973), .A2(new_n975), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n963), .B1(new_n981), .B2(new_n734), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n961), .B1(new_n982), .B2(new_n755), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n827), .A2(G68), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n398), .B1(new_n764), .B2(G159), .ZN(new_n985));
  INV_X1    g0785(.A(G143), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n984), .B(new_n985), .C1(new_n986), .C2(new_n791), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G50), .A2(new_n833), .B1(new_n780), .B2(new_n212), .ZN(new_n988));
  OAI221_X1 g0788(.A(new_n988), .B1(new_n205), .B2(new_n760), .C1(new_n818), .C2(new_n781), .ZN(new_n989));
  AOI211_X1 g0789(.A(new_n987), .B(new_n989), .C1(G150), .C2(new_n776), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n779), .A2(new_n492), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n760), .A2(new_n489), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n993), .A2(KEYINPUT46), .B1(G107), .B2(new_n827), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n994), .B1(new_n299), .B2(new_n793), .C1(new_n785), .C2(new_n791), .ZN(new_n995));
  AOI22_X1  g0795(.A1(G303), .A2(new_n776), .B1(new_n833), .B2(G283), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n765), .B2(new_n781), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n294), .B1(new_n993), .B2(KEYINPUT46), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n995), .A2(new_n997), .A3(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(new_n990), .B1(new_n992), .B2(new_n999), .ZN(new_n1000));
  XOR2_X1   g0800(.A(new_n1000), .B(KEYINPUT47), .Z(new_n1001));
  AOI21_X1  g0801(.A(new_n757), .B1(new_n1001), .B2(new_n749), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n407), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n737), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n750), .B1(new_n224), .B2(new_n1003), .C1(new_n1004), .C2(new_n239), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1002), .B(new_n1005), .C1(new_n941), .C2(new_n801), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n983), .A2(new_n1006), .ZN(G387));
  OR2_X1    g0807(.A1(new_n734), .A2(new_n978), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1008), .A2(new_n688), .A3(new_n979), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n978), .A2(new_n755), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n776), .A2(G317), .B1(G311), .B2(new_n764), .ZN(new_n1011));
  INV_X1    g0811(.A(G322), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1011), .B1(new_n761), .B2(new_n786), .C1(new_n1012), .C2(new_n791), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT48), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n830), .B2(new_n772), .C1(new_n299), .C2(new_n760), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n782), .A2(G326), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n293), .B1(G116), .B2(new_n780), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n1018), .A3(new_n1019), .A4(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(G150), .ZN(new_n1022));
  OAI22_X1  g0822(.A1(new_n775), .A2(new_n436), .B1(new_n781), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n213), .A2(new_n760), .ZN(new_n1024));
  AOI211_X1 g0824(.A(new_n1023), .B(new_n1024), .C1(G68), .C2(new_n833), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n819), .A2(new_n791), .B1(new_n793), .B2(new_n372), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n1003), .A2(new_n772), .ZN(new_n1027));
  NOR3_X1   g0827(.A1(new_n1026), .A2(new_n1027), .A3(new_n991), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1025), .A2(new_n293), .A3(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1021), .A2(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n757), .B1(new_n1030), .B2(new_n749), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n690), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n372), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1033), .A2(new_n436), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1032), .B1(new_n1034), .B2(KEYINPUT50), .ZN(new_n1035));
  OAI211_X1 g0835(.A(new_n1035), .B(new_n302), .C1(KEYINPUT50), .C2(new_n1034), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G68), .B2(G77), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n737), .B1(new_n302), .B2(new_n236), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n224), .A2(new_n399), .A3(new_n1032), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n224), .A2(G107), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n750), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1031), .B(new_n1042), .C1(new_n678), .C2(new_n801), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1009), .A2(new_n1010), .A3(new_n1043), .ZN(G393));
  OAI221_X1 g0844(.A(new_n750), .B1(new_n492), .B2(new_n224), .C1(new_n1004), .C2(new_n244), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n1033), .A2(new_n833), .B1(new_n780), .B2(G87), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n341), .B2(new_n760), .C1(new_n986), .C2(new_n781), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(G50), .B2(new_n764), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n772), .A2(new_n841), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n791), .A2(new_n1022), .B1(new_n775), .B2(new_n819), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1048), .A2(new_n293), .A3(new_n1050), .A4(new_n1052), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n791), .A2(new_n765), .B1(new_n775), .B2(new_n785), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n793), .A2(new_n761), .B1(new_n779), .B2(new_n217), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n760), .A2(new_n830), .B1(new_n786), .B2(new_n299), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n398), .B1(new_n772), .B2(new_n489), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1055), .B(new_n1059), .C1(new_n1012), .C2(new_n781), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1053), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n757), .B1(new_n1061), .B2(new_n749), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n1045), .B(new_n1062), .C1(new_n947), .C2(new_n801), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n973), .A2(new_n975), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n755), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n689), .B1(new_n1064), .B2(new_n979), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1066), .B1(new_n981), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  NAND3_X1  g0869(.A1(new_n483), .A2(G330), .A3(new_n909), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n905), .A2(new_n1070), .A3(new_n625), .ZN(new_n1071));
  INV_X1    g0871(.A(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n730), .A2(new_n660), .A3(new_n808), .ZN(new_n1073));
  AND2_X1   g0873(.A1(new_n1073), .A2(new_n809), .ZN(new_n1074));
  INV_X1    g0874(.A(KEYINPUT116), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n876), .A2(new_n1075), .A3(new_n877), .ZN(new_n1076));
  OAI21_X1  g0876(.A(KEYINPUT116), .B1(new_n914), .B2(new_n915), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n909), .A2(G330), .A3(new_n810), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n719), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n718), .B1(new_n715), .B2(G330), .ZN(new_n1083));
  OAI211_X1 g0883(.A(new_n810), .B(new_n878), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1084));
  NAND3_X1  g0884(.A1(new_n1074), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n878), .ZN(new_n1086));
  NOR2_X1   g0886(.A1(new_n1079), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n810), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n1086), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n881), .A2(new_n882), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1085), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(KEYINPUT117), .B1(new_n1072), .B2(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n901), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n900), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1094), .B1(new_n924), .B2(new_n925), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n1074), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1078), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1084), .ZN(new_n1100));
  NOR3_X1   g0900(.A1(new_n1095), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1087), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n900), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n879), .A2(new_n809), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT107), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n879), .A2(new_n880), .A3(new_n809), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1086), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g0907(.A(new_n1103), .B1(new_n1107), .B2(new_n901), .ZN(new_n1108));
  OAI221_X1 g0908(.A(new_n1094), .B1(new_n925), .B2(new_n924), .C1(new_n1074), .C2(new_n1078), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1102), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1092), .B1(new_n1101), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(KEYINPUT117), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1080), .B1(new_n813), .B2(new_n878), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1102), .B1(new_n813), .B2(new_n878), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n1074), .A2(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1116), .B2(new_n1071), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1108), .A2(new_n1109), .A3(new_n1084), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1087), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1111), .A2(new_n688), .A3(new_n1120), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1119), .A2(new_n1118), .A3(new_n755), .ZN(new_n1122));
  AOI22_X1  g0922(.A1(new_n827), .A2(G159), .B1(G137), .B2(new_n764), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(KEYINPUT54), .B(G143), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1123), .B1(new_n786), .B2(new_n1124), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT118), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n398), .B1(new_n780), .B2(G50), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n782), .A2(G125), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n825), .C2(new_n775), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1129), .B1(G128), .B2(new_n769), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n760), .A2(new_n1022), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT53), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1126), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n833), .A2(G97), .B1(G107), .B2(new_n764), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT119), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n823), .B1(new_n489), .B2(new_n775), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(G294), .B2(new_n782), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n399), .B(new_n795), .C1(G283), .C2(new_n769), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1137), .A3(new_n1050), .A4(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n757), .B1(new_n1140), .B2(new_n749), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n842), .ZN(new_n1142));
  OAI221_X1 g0942(.A(new_n1141), .B1(new_n1033), .B2(new_n1142), .C1(new_n900), .C2(new_n744), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1121), .A2(new_n1122), .A3(new_n1143), .ZN(G378));
  NAND2_X1  g0944(.A1(new_n469), .A2(new_n472), .ZN(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT55), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n458), .A2(new_n659), .ZN(new_n1147));
  XOR2_X1   g0947(.A(new_n1147), .B(KEYINPUT56), .Z(new_n1148));
  XNOR2_X1  g0948(.A(new_n1146), .B(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(new_n743), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n842), .A2(new_n436), .ZN(new_n1151));
  INV_X1    g0951(.A(G128), .ZN(new_n1152));
  OAI22_X1  g0952(.A1(new_n1152), .A2(new_n775), .B1(new_n760), .B2(new_n1124), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(G137), .B2(new_n833), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n827), .A2(G150), .B1(G125), .B2(new_n769), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n825), .C2(new_n793), .ZN(new_n1156));
  XOR2_X1   g0956(.A(new_n1156), .B(KEYINPUT120), .Z(new_n1157));
  INV_X1    g0957(.A(KEYINPUT59), .ZN(new_n1158));
  OR2_X1    g0958(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1158), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G33), .B1(new_n782), .B2(G124), .ZN(new_n1161));
  AOI21_X1  g0961(.A(G41), .B1(new_n780), .B2(G159), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n436), .B1(new_n571), .B2(G41), .ZN(new_n1164));
  OAI22_X1  g0964(.A1(new_n1003), .A2(new_n786), .B1(new_n217), .B2(new_n775), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n781), .A2(new_n830), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n779), .A2(new_n205), .ZN(new_n1167));
  OR4_X1    g0967(.A1(new_n1024), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n984), .B1(new_n791), .B2(new_n489), .C1(new_n492), .C2(new_n793), .ZN(new_n1169));
  NOR4_X1   g0969(.A1(new_n1168), .A2(new_n1169), .A3(G41), .A4(new_n293), .ZN(new_n1170));
  XOR2_X1   g0970(.A(new_n1170), .B(KEYINPUT58), .Z(new_n1171));
  NAND3_X1  g0971(.A1(new_n1163), .A2(new_n1164), .A3(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n757), .B1(new_n1172), .B2(new_n749), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1150), .A2(new_n1151), .A3(new_n1173), .ZN(new_n1174));
  AND3_X1   g0974(.A1(new_n922), .A2(new_n926), .A3(G330), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n904), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n922), .A2(new_n926), .A3(G330), .ZN(new_n1177));
  NAND4_X1  g0977(.A1(new_n1177), .A2(new_n903), .A3(new_n883), .A4(new_n902), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1176), .A2(new_n1149), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1149), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1174), .B1(new_n1181), .B2(new_n1065), .ZN(new_n1182));
  INV_X1    g0982(.A(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1149), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1184), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1176), .A2(new_n1149), .A3(new_n1178), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1119), .A2(new_n1118), .A3(new_n1091), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(new_n1072), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1190), .A3(KEYINPUT57), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1191), .A2(new_n688), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT57), .B1(new_n1188), .B2(new_n1190), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1183), .B1(new_n1192), .B2(new_n1193), .ZN(G375));
  NAND2_X1  g0994(.A1(new_n1078), .A2(new_n742), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n793), .A2(new_n489), .B1(new_n791), .B2(new_n299), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n398), .B1(new_n779), .B2(new_n841), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1196), .A2(new_n1027), .A3(new_n1197), .ZN(new_n1198));
  OAI22_X1  g0998(.A1(new_n775), .A2(new_n830), .B1(new_n786), .B2(new_n217), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1199), .B1(G97), .B2(new_n837), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n1198), .B(new_n1200), .C1(new_n761), .C2(new_n781), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT121), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n825), .A2(new_n791), .B1(new_n793), .B2(new_n1124), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G50), .B2(new_n827), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1204), .B1(new_n205), .B2(new_n779), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G137), .A2(new_n776), .B1(new_n833), .B2(G150), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n1206), .B1(new_n1152), .B2(new_n781), .C1(new_n819), .C2(new_n760), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n1205), .A2(new_n1207), .A3(new_n294), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n749), .B1(new_n1202), .B2(new_n1208), .ZN(new_n1209));
  NAND3_X1  g1009(.A1(new_n1195), .A2(new_n756), .A3(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1210), .B1(new_n341), .B2(new_n842), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1091), .B2(new_n755), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1072), .A2(new_n1091), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n962), .B1(new_n1072), .B2(new_n1091), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1212), .B1(new_n1214), .B2(new_n1215), .ZN(G381));
  AND3_X1   g1016(.A1(new_n1121), .A2(new_n1122), .A3(new_n1143), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n1217), .B(new_n1183), .C1(new_n1192), .C2(new_n1193), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(G384), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n983), .A2(new_n1068), .A3(new_n1006), .ZN(new_n1221));
  NOR4_X1   g1021(.A1(new_n1221), .A2(G396), .A3(G393), .A4(G381), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1222), .ZN(G407));
  INV_X1    g1023(.A(G213), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(G343), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT122), .Z(new_n1226));
  OAI211_X1 g1026(.A(G407), .B(G213), .C1(new_n1218), .C2(new_n1226), .ZN(G409));
  AND3_X1   g1027(.A1(new_n983), .A2(new_n1068), .A3(new_n1006), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n1068), .B1(new_n1006), .B2(new_n983), .ZN(new_n1229));
  OAI21_X1  g1029(.A(KEYINPUT125), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(G387), .A2(G390), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT125), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(new_n1232), .A3(new_n1221), .ZN(new_n1233));
  XOR2_X1   g1033(.A(G393), .B(G396), .Z(new_n1234));
  AND3_X1   g1034(.A1(new_n1230), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1234), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(G378), .A2(new_n1182), .ZN(new_n1238));
  AOI22_X1  g1038(.A1(new_n1187), .A2(new_n1186), .B1(new_n1189), .B2(new_n1072), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n962), .ZN(new_n1240));
  AOI22_X1  g1040(.A1(G375), .A2(G378), .B1(new_n1238), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT123), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1242), .B1(new_n1072), .B2(new_n1091), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1243), .A2(KEYINPUT60), .ZN(new_n1244));
  INV_X1    g1044(.A(KEYINPUT60), .ZN(new_n1245));
  OAI211_X1 g1045(.A(new_n1242), .B(new_n1245), .C1(new_n1072), .C2(new_n1091), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1244), .A2(new_n688), .A3(new_n1213), .A4(new_n1246), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1212), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1248), .A2(new_n1220), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1247), .A2(G384), .A3(new_n1212), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1241), .A2(KEYINPUT63), .A3(new_n1226), .A4(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1237), .A2(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT61), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT63), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1225), .A2(G2897), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1249), .A2(new_n1250), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT124), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(KEYINPUT124), .A3(new_n1256), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1251), .A2(new_n1226), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1259), .A2(new_n1260), .B1(new_n1261), .B2(G2897), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1225), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1241), .A2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1255), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1241), .A2(new_n1263), .A3(new_n1251), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1254), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1260), .A2(new_n1259), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1261), .A2(G2897), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT62), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1271), .A2(new_n1272), .B1(new_n1226), .B2(new_n1241), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1251), .ZN(new_n1274));
  AOI21_X1  g1074(.A(KEYINPUT61), .B1(new_n1274), .B2(KEYINPUT62), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n1266), .B2(KEYINPUT62), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1273), .A2(new_n1276), .ZN(new_n1277));
  OAI22_X1  g1077(.A1(new_n1253), .A2(new_n1268), .B1(new_n1277), .B2(new_n1237), .ZN(G405));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT57), .ZN(new_n1280));
  AND2_X1   g1080(.A1(new_n1189), .A2(new_n1072), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1280), .B1(new_n1281), .B2(new_n1181), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1282), .A2(new_n688), .A3(new_n1191), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1217), .B1(new_n1283), .B2(new_n1183), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1274), .B1(new_n1219), .B2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n689), .B1(new_n1239), .B2(KEYINPUT57), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1182), .B1(new_n1286), .B2(new_n1282), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1218), .B(new_n1251), .C1(new_n1287), .C2(new_n1217), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1279), .B1(new_n1289), .B2(KEYINPUT126), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT126), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1291), .B(KEYINPUT127), .C1(new_n1285), .C2(new_n1288), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1285), .A2(new_n1291), .A3(new_n1288), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(new_n1237), .ZN(new_n1294));
  NOR3_X1   g1094(.A1(new_n1290), .A2(new_n1292), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1288), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G375), .A2(G378), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1251), .B1(new_n1297), .B2(new_n1218), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT126), .B1(new_n1296), .B2(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1289), .A2(KEYINPUT126), .A3(new_n1279), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1300), .A2(new_n1301), .B1(new_n1237), .B2(new_n1293), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1295), .A2(new_n1302), .ZN(G402));
endmodule


