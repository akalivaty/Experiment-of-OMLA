//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n560, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n612, new_n613, new_n616, new_n617, new_n618,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT64), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT66), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT67), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n468), .B1(new_n465), .B2(KEYINPUT67), .ZN(new_n469));
  OAI21_X1  g044(.A(G2105), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  OR2_X1    g045(.A1(new_n461), .A2(new_n462), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n471), .A2(G137), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n473), .A2(KEYINPUT68), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n463), .A2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n475), .A2(new_n476), .A3(G137), .ZN(new_n477));
  AND2_X1   g052(.A1(new_n472), .A2(G2104), .ZN(new_n478));
  AOI22_X1  g053(.A1(new_n474), .A2(new_n477), .B1(G101), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n470), .A2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  NAND2_X1  g056(.A1(new_n475), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n463), .A2(new_n472), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n486));
  NAND3_X1  g061(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(G162));
  NOR2_X1   g063(.A1(new_n472), .A2(G114), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  NOR2_X1   g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n491), .B1(new_n483), .B2(G126), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n471), .A2(new_n472), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(KEYINPUT4), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n475), .A2(new_n497), .A3(G138), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n493), .B1(new_n496), .B2(new_n498), .ZN(G164));
  NAND2_X1  g074(.A1(G75), .A2(G543), .ZN(new_n500));
  XNOR2_X1  g075(.A(new_n500), .B(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G62), .ZN(new_n502));
  AND2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  NOR2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  NOR2_X1   g079(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n501), .B1(new_n502), .B2(new_n505), .ZN(new_n506));
  AND2_X1   g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(KEYINPUT6), .A2(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G543), .ZN(new_n510));
  NOR2_X1   g085(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  AOI22_X1  g086(.A1(new_n506), .A2(G651), .B1(G50), .B2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n508), .A2(new_n507), .B1(new_n503), .B2(new_n504), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT69), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g091(.A(KEYINPUT6), .B(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT69), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n516), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n512), .B1(new_n513), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT71), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT71), .ZN(new_n523));
  OAI211_X1 g098(.A(new_n512), .B(new_n523), .C1(new_n513), .C2(new_n520), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n522), .A2(new_n524), .ZN(G166));
  NAND3_X1  g100(.A1(new_n518), .A2(G63), .A3(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g103(.A1(new_n517), .A2(G51), .A3(G543), .ZN(new_n529));
  AND3_X1   g104(.A1(new_n526), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n516), .A2(G89), .A3(new_n519), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n530), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n505), .B2(new_n535), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n536), .A2(G651), .B1(new_n511), .B2(G52), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT72), .B(G90), .Z(new_n538));
  NAND3_X1  g113(.A1(new_n516), .A2(new_n519), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g115(.A(new_n540), .ZN(G171));
  AOI22_X1  g116(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(G651), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g119(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n516), .A2(G81), .A3(new_n519), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT73), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n511), .A2(G43), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n547), .B1(new_n546), .B2(new_n548), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n545), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT74), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g128(.A(KEYINPUT74), .B(new_n545), .C1(new_n549), .C2(new_n550), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  NAND4_X1  g132(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT76), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND4_X1  g137(.A1(G319), .A2(G483), .A3(G661), .A4(new_n562), .ZN(G188));
  NAND2_X1  g138(.A1(new_n511), .A2(G53), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT9), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n516), .A2(new_n519), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G91), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n518), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n543), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n565), .A2(new_n567), .A3(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n540), .A2(KEYINPUT77), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n537), .A2(new_n572), .A3(new_n539), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G301));
  INV_X1    g150(.A(G166), .ZN(G303));
  NAND3_X1  g151(.A1(new_n566), .A2(KEYINPUT78), .A3(G87), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n578));
  INV_X1    g153(.A(G87), .ZN(new_n579));
  OAI21_X1  g154(.A(new_n578), .B1(new_n520), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n518), .A2(G74), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n582), .A2(G651), .B1(new_n511), .B2(G49), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n581), .A2(new_n583), .ZN(G288));
  NAND2_X1  g159(.A1(G73), .A2(G543), .ZN(new_n585));
  INV_X1    g160(.A(G61), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n505), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n587), .A2(G651), .B1(new_n511), .B2(G48), .ZN(new_n588));
  INV_X1    g163(.A(G86), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n589), .B2(new_n520), .ZN(G305));
  NAND2_X1  g165(.A1(new_n566), .A2(G85), .ZN(new_n591));
  NAND2_X1  g166(.A1(G72), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G60), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n505), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n594), .A2(G651), .B1(new_n511), .B2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(G290));
  NAND3_X1  g171(.A1(new_n566), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n520), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(G54), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n517), .A2(G543), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT79), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n604), .B2(new_n603), .ZN(new_n606));
  AOI22_X1  g181(.A1(new_n518), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n607));
  OR2_X1    g182(.A1(new_n607), .A2(new_n543), .ZN(new_n608));
  NAND3_X1  g183(.A1(new_n601), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  MUX2_X1   g184(.A(new_n609), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g185(.A(new_n609), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g186(.A1(G286), .A2(G868), .ZN(new_n612));
  INV_X1    g187(.A(G299), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(G868), .ZN(G297));
  XOR2_X1   g189(.A(G297), .B(KEYINPUT80), .Z(G280));
  NAND2_X1  g190(.A1(new_n606), .A2(new_n608), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(new_n597), .B2(new_n600), .ZN(new_n617));
  INV_X1    g192(.A(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(G860), .ZN(G148));
  NAND2_X1  g194(.A1(new_n617), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n556), .B2(G868), .ZN(G323));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(KEYINPUT11), .ZN(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n471), .A2(new_n478), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  INV_X1    g202(.A(G2100), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n627), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n475), .A2(G135), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n483), .A2(G123), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(G2096), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND3_X1  g212(.A1(new_n629), .A2(new_n630), .A3(new_n637), .ZN(G156));
  INV_X1    g213(.A(KEYINPUT14), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2427), .B(G2438), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(G2430), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT15), .B(G2435), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n639), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n643), .B1(new_n642), .B2(new_n641), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  XNOR2_X1  g221(.A(G1341), .B(G1348), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n644), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n649), .A2(new_n650), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n651), .A2(G14), .A3(new_n652), .ZN(G401));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  XOR2_X1   g229(.A(G2084), .B(G2090), .Z(new_n655));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(KEYINPUT17), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n654), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n628), .ZN(new_n661));
  XOR2_X1   g236(.A(G2072), .B(G2078), .Z(new_n662));
  AOI21_X1  g237(.A(new_n662), .B1(new_n657), .B2(KEYINPUT18), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(new_n636), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n661), .B(new_n664), .ZN(G227));
  XOR2_X1   g240(.A(G1956), .B(G2474), .Z(new_n666));
  XOR2_X1   g241(.A(G1961), .B(G1966), .Z(new_n667));
  NAND2_X1  g242(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n668), .A2(KEYINPUT82), .ZN(new_n669));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n668), .A2(KEYINPUT82), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n669), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT20), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n666), .A2(new_n667), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n671), .B2(new_n668), .ZN(new_n676));
  NOR2_X1   g251(.A1(new_n671), .A2(KEYINPUT83), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(G1991), .B(G1996), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n681), .A2(new_n683), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n684), .A2(new_n687), .A3(new_n685), .ZN(new_n690));
  AND2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(G229));
  INV_X1    g266(.A(G29), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G26), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT28), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n475), .A2(G140), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT90), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n483), .A2(G128), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n472), .A2(G116), .ZN(new_n698));
  OAI21_X1  g273(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n699));
  OAI211_X1 g274(.A(new_n696), .B(new_n697), .C1(new_n698), .C2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT91), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n694), .B1(new_n701), .B2(new_n692), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(G2067), .ZN(new_n703));
  NOR2_X1   g278(.A1(G4), .A2(G16), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(new_n617), .B2(G16), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT89), .B(G1348), .Z(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n692), .A2(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G162), .B2(new_n692), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(KEYINPUT29), .Z(new_n711));
  INV_X1    g286(.A(G2090), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AND2_X1   g288(.A1(new_n692), .A2(G33), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n471), .A2(G127), .ZN(new_n715));
  AND2_X1   g290(.A1(G115), .A2(G2104), .ZN(new_n716));
  OAI21_X1  g291(.A(G2105), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT25), .ZN(new_n718));
  NAND2_X1  g293(.A1(G103), .A2(G2104), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n718), .B1(new_n719), .B2(G2105), .ZN(new_n720));
  NAND4_X1  g295(.A1(new_n472), .A2(KEYINPUT25), .A3(G103), .A4(G2104), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n475), .A2(G139), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n717), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n714), .B1(new_n723), .B2(G29), .ZN(new_n724));
  INV_X1    g299(.A(G2072), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  INV_X1    g302(.A(G34), .ZN(new_n728));
  AOI21_X1  g303(.A(G29), .B1(new_n728), .B2(KEYINPUT24), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(KEYINPUT24), .B2(new_n728), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(new_n480), .B2(new_n692), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2084), .ZN(new_n732));
  NAND3_X1  g307(.A1(new_n713), .A2(new_n727), .A3(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G16), .ZN(new_n734));
  NOR2_X1   g309(.A1(G171), .A2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n735), .B1(G5), .B2(new_n734), .ZN(new_n736));
  INV_X1    g311(.A(G1961), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n692), .A2(G27), .ZN(new_n740));
  OR2_X1    g315(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(KEYINPUT93), .ZN(new_n742));
  OAI211_X1 g317(.A(new_n741), .B(new_n742), .C1(G164), .C2(new_n692), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G2078), .ZN(new_n744));
  NOR2_X1   g319(.A1(G168), .A2(new_n734), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n734), .B2(G21), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g323(.A1(new_n738), .A2(new_n739), .A3(new_n744), .A4(new_n748), .ZN(new_n749));
  NAND3_X1  g324(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT26), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n751), .B1(G129), .B2(new_n483), .ZN(new_n752));
  AOI22_X1  g327(.A1(new_n475), .A2(G141), .B1(G105), .B2(new_n478), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  MUX2_X1   g329(.A(G32), .B(new_n754), .S(G29), .Z(new_n755));
  XNOR2_X1  g330(.A(KEYINPUT27), .B(G1996), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n724), .A2(new_n725), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n635), .A2(new_n692), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT30), .B(G28), .ZN(new_n760));
  OR2_X1    g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  NAND2_X1  g336(.A1(KEYINPUT31), .A2(G11), .ZN(new_n762));
  AOI22_X1  g337(.A1(new_n760), .A2(new_n692), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NAND4_X1  g338(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n763), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n746), .A2(new_n747), .B1(G2078), .B2(new_n743), .ZN(new_n765));
  NOR4_X1   g340(.A1(new_n733), .A2(new_n749), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(KEYINPUT85), .B(G16), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(G20), .ZN(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(KEYINPUT23), .Z(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G299), .B2(G16), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G1956), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(new_n711), .B2(new_n712), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(KEYINPUT94), .ZN(new_n773));
  NAND3_X1  g348(.A1(new_n708), .A2(new_n766), .A3(new_n773), .ZN(new_n774));
  INV_X1    g349(.A(new_n767), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(G19), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n556), .B2(new_n775), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(G1341), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n583), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n577), .B2(new_n580), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  INV_X1    g359(.A(new_n784), .ZN(new_n785));
  NOR2_X1   g360(.A1(new_n782), .A2(new_n783), .ZN(new_n786));
  OAI21_X1  g361(.A(G16), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n734), .A2(G23), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT88), .Z(new_n790));
  XOR2_X1   g365(.A(KEYINPUT33), .B(G1976), .Z(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n790), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n790), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n734), .A2(G6), .ZN(new_n795));
  INV_X1    g370(.A(G305), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n795), .B1(new_n796), .B2(new_n734), .ZN(new_n797));
  XOR2_X1   g372(.A(KEYINPUT32), .B(G1981), .Z(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n767), .A2(G22), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G166), .B2(new_n767), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n799), .B1(new_n801), .B2(G1971), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G1971), .B2(new_n801), .ZN(new_n803));
  NAND3_X1  g378(.A1(new_n793), .A2(new_n794), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n804), .A2(KEYINPUT34), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT34), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n793), .A2(new_n794), .A3(new_n806), .A4(new_n803), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n475), .A2(G131), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT84), .Z(new_n809));
  OAI21_X1  g384(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n810));
  INV_X1    g385(.A(G107), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(G2105), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n483), .B2(G119), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  MUX2_X1   g389(.A(G25), .B(new_n814), .S(G29), .Z(new_n815));
  XOR2_X1   g390(.A(KEYINPUT35), .B(G1991), .Z(new_n816));
  XOR2_X1   g391(.A(new_n815), .B(new_n816), .Z(new_n817));
  MUX2_X1   g392(.A(G24), .B(G290), .S(new_n775), .Z(new_n818));
  XNOR2_X1  g393(.A(KEYINPUT86), .B(G1986), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n805), .A2(new_n807), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT36), .ZN(new_n823));
  AND2_X1   g398(.A1(new_n807), .A2(new_n821), .ZN(new_n824));
  INV_X1    g399(.A(KEYINPUT36), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n824), .A2(new_n825), .A3(new_n805), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n780), .B1(new_n823), .B2(new_n826), .ZN(G311));
  NAND2_X1  g402(.A1(new_n823), .A2(new_n826), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(new_n779), .ZN(G150));
  NAND3_X1  g404(.A1(new_n516), .A2(G93), .A3(new_n519), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n511), .A2(G55), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n830), .A2(KEYINPUT97), .A3(new_n831), .ZN(new_n835));
  AND2_X1   g410(.A1(new_n518), .A2(G67), .ZN(new_n836));
  AND2_X1   g411(.A1(G80), .A2(G543), .ZN(new_n837));
  OAI211_X1 g412(.A(KEYINPUT96), .B(G651), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT96), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n837), .B1(new_n518), .B2(G67), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n839), .B1(new_n840), .B2(new_n543), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n834), .A2(new_n835), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(G860), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT99), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n845), .B(KEYINPUT37), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT98), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n546), .A2(new_n548), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT73), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n546), .A2(new_n547), .A3(new_n548), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n544), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n847), .B1(new_n851), .B2(new_n843), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n842), .A2(new_n835), .ZN(new_n853));
  AOI21_X1  g428(.A(KEYINPUT97), .B1(new_n830), .B2(new_n831), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(new_n551), .A3(KEYINPUT98), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n553), .A2(new_n554), .A3(new_n843), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n617), .A2(G559), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(KEYINPUT95), .B(KEYINPUT38), .Z(new_n862));
  XOR2_X1   g437(.A(new_n861), .B(new_n862), .Z(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  AND2_X1   g439(.A1(new_n864), .A2(KEYINPUT39), .ZN(new_n865));
  INV_X1    g440(.A(G860), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n866), .B1(new_n864), .B2(KEYINPUT39), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n846), .B1(new_n865), .B2(new_n867), .ZN(G145));
  XNOR2_X1  g443(.A(new_n814), .B(new_n626), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n723), .B(new_n754), .Z(new_n870));
  XNOR2_X1  g445(.A(new_n869), .B(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(KEYINPUT91), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n700), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n496), .A2(new_n498), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n875), .A2(new_n492), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n701), .A2(G164), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n483), .A2(G130), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n475), .A2(G142), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT101), .ZN(new_n881));
  OR3_X1    g456(.A1(new_n881), .A2(new_n472), .A3(G118), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n881), .B1(new_n472), .B2(G118), .ZN(new_n883));
  OR2_X1    g458(.A1(G106), .A2(G2105), .ZN(new_n884));
  NAND4_X1  g459(.A1(new_n882), .A2(G2104), .A3(new_n883), .A4(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n879), .A2(new_n880), .A3(new_n885), .ZN(new_n886));
  AND3_X1   g461(.A1(new_n877), .A2(new_n878), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n886), .B1(new_n877), .B2(new_n878), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n872), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n877), .A2(new_n878), .ZN(new_n890));
  INV_X1    g465(.A(new_n886), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n877), .A2(new_n878), .A3(new_n886), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(new_n893), .A3(new_n871), .ZN(new_n894));
  XOR2_X1   g469(.A(new_n487), .B(new_n635), .Z(new_n895));
  XNOR2_X1  g470(.A(new_n895), .B(KEYINPUT100), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(G160), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n889), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(G37), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g475(.A(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n897), .B1(new_n889), .B2(new_n894), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n906), .B1(new_n855), .B2(G868), .ZN(new_n907));
  XNOR2_X1  g482(.A(new_n859), .B(new_n620), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n613), .A2(new_n609), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n617), .A2(G299), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n908), .A2(KEYINPUT102), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(KEYINPUT102), .B1(new_n908), .B2(new_n912), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT103), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n613), .A2(new_n609), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(KEYINPUT103), .B1(new_n617), .B2(G299), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n917), .A3(new_n910), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT41), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT104), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n921), .B1(new_n911), .B2(new_n919), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n909), .A2(KEYINPUT104), .A3(KEYINPUT41), .A4(new_n910), .ZN(new_n923));
  AND3_X1   g498(.A1(new_n920), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n908), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n913), .A2(new_n914), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n796), .B1(new_n785), .B2(new_n786), .ZN(new_n928));
  INV_X1    g503(.A(new_n786), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n929), .A2(G305), .A3(new_n784), .ZN(new_n930));
  AND3_X1   g505(.A1(new_n522), .A2(new_n524), .A3(G290), .ZN(new_n931));
  AOI21_X1  g506(.A(G290), .B1(new_n522), .B2(new_n524), .ZN(new_n932));
  NOR2_X1   g507(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n928), .A2(new_n930), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n933), .B1(new_n928), .B2(new_n930), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n937), .B(KEYINPUT42), .ZN(new_n938));
  OR2_X1    g513(.A1(new_n927), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G868), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n927), .B2(new_n938), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n907), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n939), .A2(new_n941), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n942), .B1(KEYINPUT105), .B2(new_n943), .ZN(G295));
  AOI21_X1  g519(.A(new_n942), .B1(KEYINPUT105), .B2(new_n943), .ZN(G331));
  NAND3_X1  g520(.A1(new_n571), .A2(G168), .A3(new_n573), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT107), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(G168), .B2(new_n540), .ZN(new_n948));
  NAND3_X1  g523(.A1(G171), .A2(KEYINPUT107), .A3(G286), .ZN(new_n949));
  AND3_X1   g524(.A1(new_n946), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n950), .B1(new_n857), .B2(new_n858), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n851), .A2(new_n843), .A3(new_n847), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT98), .B1(new_n855), .B2(new_n551), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n858), .B(new_n950), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT108), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n857), .A2(KEYINPUT108), .A3(new_n858), .A4(new_n950), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n951), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OR2_X1    g533(.A1(new_n958), .A2(new_n924), .ZN(new_n959));
  NOR2_X1   g534(.A1(new_n951), .A2(new_n912), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n954), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n936), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n963), .A2(KEYINPUT109), .A3(new_n934), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n965), .B1(new_n935), .B2(new_n936), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n968), .ZN(new_n969));
  OAI211_X1 g544(.A(new_n937), .B(new_n961), .C1(new_n958), .C2(new_n924), .ZN(new_n970));
  AND2_X1   g545(.A1(new_n970), .A2(new_n899), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT43), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n969), .A2(new_n971), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(KEYINPUT112), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n956), .A2(new_n957), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT110), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n975), .A2(new_n976), .A3(new_n960), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n976), .B1(new_n975), .B2(new_n960), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n918), .A2(KEYINPUT41), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(KEYINPUT41), .B2(new_n911), .ZN(new_n980));
  INV_X1    g555(.A(new_n951), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(new_n954), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n977), .A2(new_n978), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n971), .B1(new_n983), .B2(new_n967), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n986));
  NAND4_X1  g561(.A1(new_n969), .A2(new_n971), .A3(new_n986), .A4(new_n972), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n974), .A2(KEYINPUT44), .A3(new_n985), .A4(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n971), .B(new_n972), .C1(new_n983), .C2(new_n967), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n967), .B1(new_n959), .B2(new_n961), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n970), .A2(new_n899), .ZN(new_n991));
  OAI21_X1  g566(.A(KEYINPUT43), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(KEYINPUT106), .B(KEYINPUT44), .ZN(new_n994));
  INV_X1    g569(.A(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(KEYINPUT111), .B1(new_n993), .B2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT111), .ZN(new_n997));
  AOI211_X1 g572(.A(new_n997), .B(new_n994), .C1(new_n989), .C2(new_n992), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n988), .B1(new_n996), .B2(new_n998), .ZN(G397));
  NAND2_X1  g574(.A1(new_n874), .A2(G2067), .ZN(new_n1000));
  INV_X1    g575(.A(G2067), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n701), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n754), .B(G1996), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n814), .B(new_n816), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n470), .A2(new_n479), .A3(G40), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT45), .B1(new_n876), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n470), .A2(new_n479), .A3(KEYINPUT113), .A4(G40), .ZN(new_n1013));
  AND3_X1   g588(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1007), .A2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(G290), .A2(G1986), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT114), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(new_n1014), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(G1986), .A3(G290), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  OR2_X1    g595(.A1(new_n1020), .A2(KEYINPUT115), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(KEYINPUT115), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1015), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n1023), .B(KEYINPUT116), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT57), .ZN(new_n1025));
  OAI21_X1  g600(.A(G299), .B1(KEYINPUT121), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(KEYINPUT121), .ZN(new_n1027));
  XNOR2_X1  g602(.A(new_n1026), .B(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n876), .A2(new_n1030), .A3(new_n1011), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1010), .A2(new_n1029), .A3(new_n1013), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(G1956), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n876), .A2(new_n1011), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT45), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1037), .A2(new_n1010), .A3(new_n1013), .A4(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1040));
  XNOR2_X1  g615(.A(new_n1040), .B(G2072), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1028), .B(new_n1034), .C1(new_n1039), .C2(new_n1042), .ZN(new_n1043));
  AND2_X1   g618(.A1(new_n1043), .A2(new_n617), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G164), .A2(G1384), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1010), .A2(new_n1045), .A3(new_n1013), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT123), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1010), .A2(KEYINPUT123), .A3(new_n1045), .A4(new_n1013), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1001), .ZN(new_n1051));
  INV_X1    g626(.A(G1348), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1032), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1051), .A2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1034), .B1(new_n1039), .B2(new_n1042), .ZN(new_n1055));
  INV_X1    g630(.A(new_n1028), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1044), .A2(new_n1054), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1056), .ZN(new_n1058));
  INV_X1    g633(.A(KEYINPUT61), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1058), .A2(new_n1043), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1059), .B1(new_n1058), .B2(new_n1043), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT59), .ZN(new_n1062));
  XOR2_X1   g637(.A(KEYINPUT58), .B(G1341), .Z(new_n1063));
  NAND3_X1  g638(.A1(new_n1048), .A2(new_n1049), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1039), .ZN(new_n1065));
  INV_X1    g640(.A(G1996), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1064), .A2(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1062), .B1(new_n1068), .B2(new_n556), .ZN(new_n1069));
  AOI211_X1 g644(.A(KEYINPUT59), .B(new_n555), .C1(new_n1064), .C2(new_n1067), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1060), .A2(new_n1061), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n617), .B1(new_n1054), .B2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1051), .A2(KEYINPUT60), .A3(new_n609), .A4(new_n1053), .ZN(new_n1074));
  AOI22_X1  g649(.A1(new_n1073), .A2(new_n1074), .B1(new_n1072), .B2(new_n1054), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1057), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(G305), .A2(G1981), .ZN(new_n1077));
  XNOR2_X1  g652(.A(KEYINPUT119), .B(G86), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n566), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1079), .A2(new_n588), .ZN(new_n1080));
  AOI21_X1  g655(.A(new_n1077), .B1(G1981), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT49), .ZN(new_n1082));
  XNOR2_X1  g657(.A(new_n1081), .B(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1046), .A2(G8), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G1976), .ZN(new_n1087));
  NOR3_X1   g662(.A1(new_n785), .A2(new_n1087), .A3(new_n786), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT52), .B1(new_n1088), .B2(new_n1084), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n1088), .A2(new_n1084), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT52), .B1(G288), .B2(new_n1087), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT118), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1091), .A2(new_n1095), .A3(new_n1092), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1090), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g672(.A1(new_n1065), .A2(G1971), .B1(G2090), .B2(new_n1032), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n1099));
  OAI211_X1 g674(.A(G303), .B(G8), .C1(new_n1099), .C2(KEYINPUT55), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G8), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1102), .B1(G166), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1104), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1098), .A2(G8), .A3(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1105), .B1(new_n1098), .B2(G8), .ZN(new_n1108));
  NOR2_X1   g683(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT53), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1110), .A2(G2078), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT125), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1008), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1112), .B1(new_n1037), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g689(.A1(new_n1012), .A2(KEYINPUT125), .A3(new_n1008), .ZN(new_n1115));
  OAI211_X1 g690(.A(new_n1038), .B(new_n1111), .C1(new_n1114), .C2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1110), .B1(new_n1039), .B2(G2078), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1032), .A2(new_n737), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(G171), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1037), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1121), .A2(KEYINPUT120), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1037), .A2(new_n1010), .A3(new_n1123), .A4(new_n1013), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1122), .A2(new_n1124), .A3(new_n1038), .A4(new_n1111), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1125), .A2(G301), .A3(new_n1117), .A4(new_n1118), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1120), .A2(new_n1126), .A3(KEYINPUT54), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1097), .A2(new_n1109), .A3(new_n1127), .ZN(new_n1128));
  OR2_X1    g703(.A1(new_n1119), .A2(new_n574), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1125), .A2(new_n1117), .A3(new_n1118), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(new_n574), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT54), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1128), .A2(new_n1132), .ZN(new_n1133));
  NOR2_X1   g708(.A1(new_n1032), .A2(G2084), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1122), .A2(new_n1124), .A3(new_n1038), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(new_n1135), .B2(new_n747), .ZN(new_n1136));
  NOR3_X1   g711(.A1(new_n1136), .A2(new_n1103), .A3(G168), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT51), .ZN(new_n1138));
  AOI211_X1 g713(.A(G286), .B(new_n1134), .C1(new_n1135), .C2(new_n747), .ZN(new_n1139));
  NOR2_X1   g714(.A1(new_n1103), .A2(KEYINPUT124), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1138), .B1(new_n1139), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1136), .A2(G168), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1143), .A2(KEYINPUT51), .A3(new_n1140), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1137), .B1(new_n1142), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1145), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1076), .A2(new_n1133), .A3(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1097), .A2(new_n1107), .ZN(new_n1148));
  AOI211_X1 g723(.A(G1976), .B(G288), .C1(new_n1083), .C2(new_n1085), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1085), .B1(new_n1149), .B2(new_n1077), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1148), .A2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n1136), .A2(new_n1103), .A3(G286), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1097), .A2(new_n1109), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT63), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1097), .A2(new_n1109), .A3(new_n1152), .A4(KEYINPUT63), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1151), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1147), .A2(new_n1157), .ZN(new_n1158));
  AND4_X1   g733(.A1(new_n574), .A2(new_n1097), .A3(new_n1109), .A4(new_n1130), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT62), .ZN(new_n1160));
  OAI21_X1  g735(.A(new_n1159), .B1(new_n1145), .B2(new_n1160), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1145), .A2(new_n1160), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1024), .B1(new_n1158), .B2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1014), .B1(new_n1003), .B2(new_n754), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1014), .A2(new_n1066), .ZN(new_n1166));
  AND2_X1   g741(.A1(new_n1166), .A2(KEYINPUT46), .ZN(new_n1167));
  NOR2_X1   g742(.A1(new_n1166), .A2(KEYINPUT46), .ZN(new_n1168));
  OAI21_X1  g743(.A(new_n1165), .B1(new_n1167), .B2(new_n1168), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n1169), .B(KEYINPUT126), .Z(new_n1170));
  NAND2_X1  g745(.A1(new_n1170), .A2(KEYINPUT47), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1017), .A2(KEYINPUT48), .A3(new_n1014), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT48), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1007), .A2(new_n1014), .B1(new_n1173), .B2(new_n1018), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1005), .A2(new_n816), .A3(new_n809), .A4(new_n813), .ZN(new_n1175));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1002), .ZN(new_n1176));
  AOI22_X1  g751(.A1(new_n1172), .A2(new_n1174), .B1(new_n1176), .B2(new_n1014), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1171), .A2(new_n1177), .ZN(new_n1178));
  NOR2_X1   g753(.A1(new_n1170), .A2(KEYINPUT47), .ZN(new_n1179));
  NOR2_X1   g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1164), .A2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g756(.A1(G401), .A2(new_n459), .A3(G227), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n1183), .B1(new_n689), .B2(new_n690), .ZN(new_n1184));
  OAI21_X1  g758(.A(new_n1184), .B1(new_n900), .B2(new_n902), .ZN(new_n1185));
  AOI21_X1  g759(.A(new_n1185), .B1(new_n989), .B2(new_n992), .ZN(new_n1186));
  XNOR2_X1  g760(.A(new_n1186), .B(KEYINPUT127), .ZN(G308));
  INV_X1    g761(.A(new_n1186), .ZN(G225));
endmodule


