//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 1 1 1 0 1 0 0 1 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:01 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n753, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n773, new_n774, new_n775, new_n776,
    new_n778, new_n779, new_n780, new_n781, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n791, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n876, new_n877, new_n878,
    new_n879, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n944,
    new_n945, new_n946, new_n947, new_n949, new_n950, new_n951, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  INV_X1    g002(.A(G29gat), .ZN(new_n204));
  INV_X1    g003(.A(G36gat), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT88), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n208), .B(new_n209), .ZN(new_n210));
  XOR2_X1   g009(.A(G43gat), .B(G50gat), .Z(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT85), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT85), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT87), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n210), .A2(new_n216), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n207), .A2(KEYINPUT86), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n206), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n207), .A2(KEYINPUT86), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n218), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n224), .A2(KEYINPUT15), .A3(new_n212), .A4(new_n215), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n220), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT17), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT89), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(new_n226), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n232));
  XNOR2_X1  g031(.A(G15gat), .B(G22gat), .ZN(new_n233));
  INV_X1    g032(.A(G1gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT16), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G1gat), .B2(new_n233), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(G8gat), .Z(new_n238));
  AND2_X1   g037(.A1(new_n232), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n230), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(G229gat), .A2(G233gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n238), .B(KEYINPUT90), .ZN(new_n242));
  OR2_X1    g041(.A1(new_n242), .A2(new_n231), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n240), .A2(new_n243), .A3(KEYINPUT18), .A4(new_n241), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n242), .B(new_n231), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT91), .B(KEYINPUT13), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(new_n241), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n246), .A2(new_n247), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G141gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G197gat), .ZN(new_n255));
  XOR2_X1   g054(.A(KEYINPUT11), .B(G169gat), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(new_n257), .B(KEYINPUT12), .Z(new_n258));
  NOR2_X1   g057(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(new_n258), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n244), .A2(new_n245), .B1(new_n248), .B2(new_n251), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n260), .B1(new_n261), .B2(new_n247), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n202), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n253), .A2(new_n258), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n261), .A2(new_n260), .A3(new_n247), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n264), .A2(KEYINPUT92), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n263), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  XOR2_X1   g067(.A(G8gat), .B(G36gat), .Z(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT77), .ZN(new_n270));
  XNOR2_X1  g069(.A(G64gat), .B(G92gat), .ZN(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  XNOR2_X1  g071(.A(G197gat), .B(G204gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT22), .ZN(new_n274));
  INV_X1    g073(.A(G211gat), .ZN(new_n275));
  INV_X1    g074(.A(G218gat), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n274), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n273), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(G211gat), .B(G218gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n279), .A2(new_n273), .A3(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(G190gat), .ZN(new_n284));
  INV_X1    g083(.A(G183gat), .ZN(new_n285));
  OAI211_X1 g084(.A(KEYINPUT67), .B(new_n284), .C1(new_n285), .C2(KEYINPUT27), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT28), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n285), .B2(KEYINPUT27), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT27), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(G183gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n286), .B(new_n287), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(G190gat), .B1(new_n289), .B2(G183gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n285), .A2(KEYINPUT27), .ZN(new_n293));
  OAI211_X1 g092(.A(new_n292), .B(new_n293), .C1(KEYINPUT67), .C2(KEYINPUT28), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT68), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT68), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n298), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G169gat), .A2(G176gat), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT64), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT64), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n305), .B1(G169gat), .B2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT26), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n304), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n300), .A2(new_n301), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(G183gat), .A2(G190gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NAND4_X1  g112(.A1(new_n295), .A2(new_n309), .A3(KEYINPUT69), .A4(new_n310), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT25), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT23), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n303), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n316), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n304), .A2(new_n306), .A3(KEYINPUT23), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT65), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n310), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT24), .ZN(new_n324));
  NAND3_X1  g123(.A1(KEYINPUT65), .A2(G183gat), .A3(G190gat), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n323), .A2(new_n324), .A3(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n327));
  OAI21_X1  g126(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n328));
  INV_X1    g127(.A(new_n328), .ZN(new_n329));
  NOR3_X1   g128(.A1(KEYINPUT66), .A2(G183gat), .A3(G190gat), .ZN(new_n330));
  OAI211_X1 g129(.A(new_n326), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n310), .A2(new_n324), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n285), .A2(new_n284), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n332), .A2(new_n327), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n318), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n302), .A2(new_n303), .A3(KEYINPUT23), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI22_X1  g136(.A1(new_n321), .A2(new_n331), .B1(new_n337), .B2(new_n316), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n315), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(KEYINPUT74), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT74), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n315), .A2(new_n342), .A3(new_n339), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT75), .B(KEYINPUT29), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G226gat), .A2(G233gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n347), .ZN(new_n349));
  INV_X1    g148(.A(new_n311), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n349), .B1(new_n350), .B2(new_n338), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT76), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n283), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n283), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n342), .B1(new_n315), .B2(new_n339), .ZN(new_n356));
  AOI211_X1 g155(.A(KEYINPUT74), .B(new_n338), .C1(new_n313), .C2(new_n314), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n349), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI211_X1 g157(.A(KEYINPUT29), .B(new_n349), .C1(new_n339), .C2(new_n311), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n355), .B1(new_n358), .B2(new_n360), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n272), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n360), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n283), .ZN(new_n364));
  INV_X1    g163(.A(new_n272), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n352), .B1(new_n346), .B2(new_n347), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n364), .B(new_n365), .C1(new_n366), .C2(new_n283), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n362), .A2(KEYINPUT30), .A3(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n356), .A2(new_n357), .A3(new_n344), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n353), .B1(new_n369), .B2(new_n349), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n361), .B1(new_n370), .B2(new_n355), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT30), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n371), .A2(new_n372), .A3(new_n365), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n376));
  NAND2_X1  g175(.A1(G155gat), .A2(G162gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(KEYINPUT2), .ZN(new_n378));
  INV_X1    g177(.A(G141gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n379), .A2(G148gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n381), .A2(G141gat), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n376), .B(new_n378), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  XNOR2_X1  g182(.A(G155gat), .B(G162gat), .ZN(new_n384));
  INV_X1    g183(.A(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(G141gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n379), .A2(G148gat), .ZN(new_n389));
  AOI21_X1  g188(.A(KEYINPUT78), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n390), .A2(new_n384), .A3(new_n378), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n386), .A2(new_n387), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n345), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(new_n355), .ZN(new_n394));
  NAND2_X1  g193(.A1(G228gat), .A2(G233gat), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n383), .A2(new_n385), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n384), .B1(new_n390), .B2(new_n378), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT29), .ZN(new_n400));
  AOI21_X1  g199(.A(KEYINPUT3), .B1(new_n283), .B2(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n394), .B(new_n396), .C1(new_n399), .C2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT79), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n397), .B2(new_n398), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n386), .A2(KEYINPUT79), .A3(new_n391), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n344), .B1(new_n281), .B2(new_n282), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n405), .C1(KEYINPUT3), .C2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n394), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT82), .B1(new_n408), .B2(new_n395), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n410));
  AOI211_X1 g209(.A(new_n410), .B(new_n396), .C1(new_n407), .C2(new_n394), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n402), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(KEYINPUT31), .B(G50gat), .Z(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G78gat), .B(G106gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(G22gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n413), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n417), .B(new_n402), .C1(new_n409), .C2(new_n411), .ZN(new_n418));
  AND3_X1   g217(.A1(new_n414), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n416), .B1(new_n414), .B2(new_n418), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT32), .ZN(new_n422));
  INV_X1    g221(.A(G113gat), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(G120gat), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(G120gat), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G113gat), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n423), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n426), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT1), .ZN(new_n431));
  XNOR2_X1  g230(.A(G127gat), .B(G134gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NOR2_X1   g232(.A1(new_n423), .A2(G120gat), .ZN(new_n434));
  NOR2_X1   g233(.A1(new_n427), .A2(G113gat), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n431), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  XOR2_X1   g235(.A(G127gat), .B(G134gat), .Z(new_n437));
  AOI21_X1  g236(.A(KEYINPUT70), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(KEYINPUT1), .B1(new_n428), .B2(new_n424), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n439), .A2(new_n440), .A3(new_n432), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n433), .B1(new_n438), .B2(new_n441), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n315), .B2(new_n339), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n436), .A2(KEYINPUT70), .A3(new_n437), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n440), .B1(new_n439), .B2(new_n432), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n437), .A2(KEYINPUT1), .ZN(new_n446));
  AOI22_X1  g245(.A1(new_n444), .A2(new_n445), .B1(new_n446), .B2(new_n430), .ZN(new_n447));
  AOI211_X1 g246(.A(new_n447), .B(new_n338), .C1(new_n313), .C2(new_n314), .ZN(new_n448));
  NOR2_X1   g247(.A1(new_n443), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(G227gat), .A2(G233gat), .ZN(new_n450));
  INV_X1    g249(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n422), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT34), .B1(new_n451), .B2(KEYINPUT73), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n340), .A2(new_n447), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n315), .A2(new_n442), .A3(new_n339), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n453), .B1(new_n456), .B2(new_n450), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n450), .B(new_n453), .C1(new_n443), .C2(new_n448), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n452), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n453), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n461), .B1(new_n449), .B2(new_n451), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n454), .A2(new_n451), .A3(new_n455), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(KEYINPUT32), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(new_n464), .A3(new_n458), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT72), .B(KEYINPUT33), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  XOR2_X1   g267(.A(G15gat), .B(G43gat), .Z(new_n469));
  XNOR2_X1  g268(.A(G71gat), .B(G99gat), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n469), .B(new_n470), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n466), .A2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(KEYINPUT35), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n460), .A2(new_n472), .A3(new_n465), .ZN(new_n476));
  NAND4_X1  g275(.A1(new_n421), .A2(new_n474), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n375), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT83), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT6), .ZN(new_n480));
  OAI21_X1  g279(.A(KEYINPUT3), .B1(new_n397), .B2(new_n398), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n442), .A2(new_n481), .A3(new_n392), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT5), .ZN(new_n483));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n386), .A2(new_n391), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n487), .B1(new_n442), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n447), .A2(new_n399), .A3(KEYINPUT80), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n486), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n405), .ZN(new_n492));
  AOI21_X1  g291(.A(KEYINPUT79), .B1(new_n386), .B2(new_n391), .ZN(new_n493));
  OAI211_X1 g292(.A(new_n486), .B(new_n447), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n485), .B1(new_n491), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT81), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT81), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n485), .B(new_n498), .C1(new_n491), .C2(new_n495), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n442), .A2(new_n487), .A3(new_n488), .ZN(new_n500));
  AOI21_X1  g299(.A(KEYINPUT80), .B1(new_n447), .B2(new_n399), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n486), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(KEYINPUT4), .B(new_n447), .C1(new_n492), .C2(new_n493), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n502), .A2(new_n503), .A3(new_n484), .A4(new_n482), .ZN(new_n504));
  OAI22_X1  g303(.A1(new_n500), .A2(new_n501), .B1(new_n399), .B2(new_n447), .ZN(new_n505));
  INV_X1    g304(.A(new_n484), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n483), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  AOI22_X1  g306(.A1(new_n497), .A2(new_n499), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g307(.A(G1gat), .B(G29gat), .ZN(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT0), .ZN(new_n510));
  XNOR2_X1  g309(.A(G57gat), .B(G85gat), .ZN(new_n511));
  XOR2_X1   g310(.A(new_n510), .B(new_n511), .Z(new_n512));
  OAI21_X1  g311(.A(new_n480), .B1(new_n508), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n499), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n507), .A2(new_n504), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n514), .A2(new_n512), .A3(new_n515), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n479), .B1(new_n513), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(KEYINPUT4), .B1(new_n500), .B2(new_n501), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n494), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n498), .B1(new_n519), .B2(new_n485), .ZN(new_n520));
  INV_X1    g319(.A(new_n499), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n515), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n512), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT6), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n522), .A2(new_n523), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n514), .A2(new_n512), .A3(new_n515), .ZN(new_n526));
  NAND4_X1  g325(.A1(new_n525), .A2(KEYINPUT83), .A3(new_n480), .A4(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n517), .A2(new_n524), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n478), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n525), .A2(new_n480), .A3(new_n526), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n524), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n374), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n421), .A2(new_n474), .A3(new_n476), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT84), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AND3_X1   g334(.A1(new_n460), .A2(new_n472), .A3(new_n465), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n472), .B1(new_n460), .B2(new_n465), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n538), .A2(KEYINPUT84), .A3(new_n421), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n532), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n529), .B1(new_n540), .B2(new_n475), .ZN(new_n541));
  INV_X1    g340(.A(new_n421), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n532), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT36), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n544), .B1(new_n536), .B2(new_n537), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n474), .A2(KEYINPUT36), .A3(new_n476), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT38), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT37), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n365), .B1(new_n371), .B2(new_n549), .ZN(new_n550));
  OAI21_X1  g349(.A(KEYINPUT37), .B1(new_n354), .B2(new_n361), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n364), .B(new_n549), .C1(new_n366), .C2(new_n283), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(new_n272), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n341), .A2(new_n343), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n359), .B1(new_n555), .B2(new_n349), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT37), .B1(new_n556), .B2(new_n283), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n355), .B1(new_n348), .B2(new_n353), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n548), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n367), .B1(new_n554), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n528), .A2(new_n552), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT39), .ZN(new_n562));
  AOI22_X1  g361(.A1(new_n489), .A2(new_n490), .B1(new_n488), .B2(new_n442), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n563), .B2(new_n484), .ZN(new_n564));
  INV_X1    g363(.A(new_n482), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n565), .B1(new_n518), .B2(new_n494), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n564), .B1(new_n566), .B2(new_n484), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n482), .B1(new_n491), .B2(new_n495), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n562), .A3(new_n506), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n567), .A2(new_n512), .A3(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT40), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n567), .A2(KEYINPUT40), .A3(new_n512), .A4(new_n569), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n572), .A2(new_n525), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n574), .A2(new_n368), .A3(new_n373), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n575), .A2(new_n421), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n543), .B(new_n547), .C1(new_n561), .C2(new_n576), .ZN(new_n577));
  AOI21_X1  g376(.A(new_n268), .B1(new_n541), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n579));
  NAND2_X1  g378(.A1(G85gat), .A2(G92gat), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT7), .ZN(new_n581));
  NAND2_X1  g380(.A1(G99gat), .A2(G106gat), .ZN(new_n582));
  INV_X1    g381(.A(G85gat), .ZN(new_n583));
  INV_X1    g382(.A(G92gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(KEYINPUT8), .A2(new_n582), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  AND2_X1   g385(.A1(G99gat), .A2(G106gat), .ZN(new_n587));
  NOR2_X1   g386(.A1(G99gat), .A2(G106gat), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n579), .B1(new_n586), .B2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n589), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n581), .A2(new_n591), .A3(KEYINPUT97), .A4(new_n585), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n586), .A2(new_n589), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n230), .A2(new_n232), .A3(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n226), .ZN(new_n599));
  AND3_X1   g398(.A1(new_n596), .A2(new_n284), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n284), .B1(new_n596), .B2(new_n599), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n276), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n599), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n603), .A2(G190gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n596), .A2(new_n284), .A3(new_n599), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(G218gat), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT96), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G134gat), .B(G162gat), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(G64gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n614), .A2(G57gat), .ZN(new_n615));
  INV_X1    g414(.A(G57gat), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(G64gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n618), .B1(KEYINPUT93), .B2(KEYINPUT9), .ZN(new_n619));
  INV_X1    g418(.A(G71gat), .ZN(new_n620));
  INV_X1    g419(.A(G78gat), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  OR3_X1    g421(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT93), .ZN(new_n623));
  OAI21_X1  g422(.A(KEYINPUT93), .B1(new_n620), .B2(new_n621), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n619), .A2(new_n622), .A3(new_n623), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT9), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n626), .B1(new_n620), .B2(new_n621), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n615), .A2(KEYINPUT94), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n628), .A2(new_n617), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n615), .A2(KEYINPUT94), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n627), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  AOI21_X1  g430(.A(KEYINPUT21), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(G231gat), .A2(G233gat), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G127gat), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n625), .A2(new_n631), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT95), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n242), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n635), .B(new_n639), .Z(new_n640));
  XNOR2_X1  g439(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G155gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(G183gat), .B(G211gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n640), .B(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n602), .A2(new_n606), .A3(new_n607), .A4(new_n611), .ZN(new_n646));
  INV_X1    g445(.A(new_n594), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n636), .B1(new_n647), .B2(KEYINPUT98), .ZN(new_n648));
  OR2_X1    g447(.A1(new_n647), .A2(KEYINPUT98), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n648), .A2(new_n593), .A3(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(KEYINPUT99), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n595), .A2(new_n636), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT99), .ZN(new_n654));
  NAND4_X1  g453(.A1(new_n648), .A2(new_n649), .A3(new_n654), .A4(new_n593), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n651), .A2(new_n652), .A3(new_n653), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n637), .A2(new_n598), .A3(KEYINPUT10), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(G230gat), .A2(G233gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n651), .A2(new_n653), .A3(new_n655), .ZN(new_n661));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n663), .A2(KEYINPUT100), .ZN(new_n664));
  XOR2_X1   g463(.A(G120gat), .B(G148gat), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT101), .ZN(new_n666));
  XNOR2_X1  g465(.A(G176gat), .B(G204gat), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n666), .B(new_n667), .Z(new_n668));
  INV_X1    g467(.A(KEYINPUT100), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n661), .A2(new_n669), .A3(new_n662), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n660), .A2(new_n664), .A3(new_n668), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n668), .ZN(new_n673));
  INV_X1    g472(.A(new_n663), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n662), .B1(new_n656), .B2(new_n657), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT102), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT102), .B(new_n673), .C1(new_n674), .C2(new_n675), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n672), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n613), .A2(new_n645), .A3(new_n646), .A4(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT103), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n613), .A2(new_n646), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND4_X1  g484(.A1(new_n685), .A2(KEYINPUT103), .A3(new_n645), .A4(new_n680), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n578), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  NOR2_X1   g486(.A1(new_n687), .A2(new_n531), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(new_n234), .ZN(G1324gat));
  INV_X1    g488(.A(new_n687), .ZN(new_n690));
  XOR2_X1   g489(.A(KEYINPUT16), .B(G8gat), .Z(new_n691));
  NAND3_X1  g490(.A1(new_n690), .A2(new_n375), .A3(new_n691), .ZN(new_n692));
  OAI21_X1  g491(.A(G8gat), .B1(new_n687), .B2(new_n374), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g493(.A(new_n692), .B(new_n694), .S(KEYINPUT42), .Z(G1325gat));
  INV_X1    g494(.A(new_n538), .ZN(new_n696));
  OR3_X1    g495(.A1(new_n687), .A2(G15gat), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(G15gat), .B1(new_n687), .B2(new_n547), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(G1326gat));
  NOR2_X1   g498(.A1(new_n687), .A2(new_n421), .ZN(new_n700));
  XOR2_X1   g499(.A(KEYINPUT43), .B(G22gat), .Z(new_n701));
  XNOR2_X1  g500(.A(new_n700), .B(new_n701), .ZN(G1327gat));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n703));
  AOI211_X1 g502(.A(new_n703), .B(new_n685), .C1(new_n541), .C2(new_n577), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n535), .A2(new_n539), .ZN(new_n705));
  AOI22_X1  g504(.A1(new_n368), .A2(new_n373), .B1(new_n530), .B2(new_n524), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n475), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n477), .ZN(new_n708));
  AND3_X1   g507(.A1(new_n708), .A2(new_n528), .A3(new_n374), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n577), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  AOI21_X1  g509(.A(KEYINPUT44), .B1(new_n710), .B2(new_n684), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  INV_X1    g512(.A(new_n531), .ZN(new_n714));
  INV_X1    g513(.A(new_n680), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n715), .A2(new_n645), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n264), .A2(new_n265), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n712), .A2(new_n713), .A3(new_n714), .A4(new_n719), .ZN(new_n720));
  AOI21_X1  g519(.A(KEYINPUT84), .B1(new_n538), .B2(new_n421), .ZN(new_n721));
  AND4_X1   g520(.A1(KEYINPUT84), .A2(new_n421), .A3(new_n476), .A4(new_n474), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n706), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n723), .A2(KEYINPUT35), .B1(new_n528), .B2(new_n478), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n547), .B1(new_n706), .B2(new_n421), .ZN(new_n725));
  OR3_X1    g524(.A1(new_n528), .A2(new_n552), .A3(new_n560), .ZN(new_n726));
  INV_X1    g525(.A(new_n576), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n684), .B1(new_n724), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n703), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n710), .A2(KEYINPUT44), .A3(new_n684), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n730), .A2(new_n714), .A3(new_n731), .A4(new_n719), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT105), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n720), .A2(new_n733), .A3(G29gat), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n716), .A2(new_n684), .ZN(new_n735));
  OAI211_X1 g534(.A(new_n267), .B(new_n735), .C1(new_n724), .C2(new_n728), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n714), .A2(new_n204), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT104), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT104), .ZN(new_n739));
  INV_X1    g538(.A(new_n737), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n578), .A2(new_n739), .A3(new_n735), .A4(new_n740), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n738), .A2(KEYINPUT45), .A3(new_n741), .ZN(new_n742));
  AOI21_X1  g541(.A(KEYINPUT45), .B1(new_n738), .B2(new_n741), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n734), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT106), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n734), .A2(new_n744), .A3(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n746), .A2(new_n748), .ZN(G1328gat));
  NOR3_X1   g548(.A1(new_n736), .A2(G36gat), .A3(new_n374), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT46), .ZN(new_n751));
  INV_X1    g550(.A(new_n712), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n374), .A3(new_n718), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(new_n205), .ZN(G1329gat));
  OR2_X1    g553(.A1(new_n696), .A2(G43gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n736), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT107), .ZN(new_n757));
  INV_X1    g556(.A(new_n547), .ZN(new_n758));
  NAND4_X1  g557(.A1(new_n730), .A2(new_n758), .A3(new_n731), .A4(new_n719), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G43gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n761), .B(new_n762), .ZN(G1330gat));
  OR3_X1    g562(.A1(new_n736), .A2(G50gat), .A3(new_n421), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n730), .A2(new_n542), .A3(new_n731), .A4(new_n719), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(G50gat), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(KEYINPUT108), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT48), .B(new_n764), .C1(new_n767), .C2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n765), .A2(G50gat), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n764), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(KEYINPUT48), .B2(new_n771), .ZN(G1331gat));
  INV_X1    g571(.A(new_n645), .ZN(new_n773));
  NOR4_X1   g572(.A1(new_n684), .A2(new_n773), .A3(new_n717), .A4(new_n680), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n710), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n775), .A2(new_n531), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(new_n616), .ZN(G1332gat));
  XNOR2_X1  g576(.A(new_n775), .B(KEYINPUT109), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n375), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n780));
  XOR2_X1   g579(.A(KEYINPUT49), .B(G64gat), .Z(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(G1333gat));
  AOI21_X1  g581(.A(new_n620), .B1(new_n778), .B2(new_n758), .ZN(new_n783));
  XNOR2_X1  g582(.A(new_n538), .B(KEYINPUT110), .ZN(new_n784));
  NOR3_X1   g583(.A1(new_n775), .A2(G71gat), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g584(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  OR3_X1    g586(.A1(new_n783), .A2(new_n785), .A3(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n787), .B1(new_n783), .B2(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(G1334gat));
  NAND2_X1  g589(.A1(new_n778), .A2(new_n542), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g591(.A1(new_n645), .A2(new_n717), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n710), .A2(new_n684), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT51), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n795), .A2(new_n680), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n796), .A2(new_n583), .A3(new_n714), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n793), .A2(new_n715), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n752), .A2(new_n531), .A3(new_n798), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n797), .B1(new_n583), .B2(new_n799), .ZN(G1336gat));
  INV_X1    g599(.A(new_n798), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n712), .A2(new_n375), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n715), .A2(new_n584), .A3(new_n375), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n803), .B1(new_n795), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(KEYINPUT52), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n803), .B(new_n807), .C1(new_n795), .C2(new_n804), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(G1337gat));
  INV_X1    g608(.A(G99gat), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n796), .A2(new_n810), .A3(new_n538), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n712), .A2(new_n758), .A3(new_n801), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(G99gat), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n812), .A2(new_n813), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n811), .B1(new_n815), .B2(new_n816), .ZN(G1338gat));
  NAND3_X1  g616(.A1(new_n712), .A2(new_n542), .A3(new_n801), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(G106gat), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT53), .ZN(new_n820));
  NOR3_X1   g619(.A1(new_n680), .A2(G106gat), .A3(new_n421), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n819), .B(new_n820), .C1(new_n795), .C2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(new_n795), .ZN(new_n824));
  XOR2_X1   g623(.A(new_n821), .B(KEYINPUT113), .Z(new_n825));
  AOI22_X1  g624(.A1(new_n824), .A2(new_n825), .B1(new_n818), .B2(G106gat), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n823), .B1(new_n826), .B2(new_n820), .ZN(G1339gat));
  NOR2_X1   g626(.A1(new_n681), .A2(new_n717), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n656), .A2(new_n662), .A3(new_n657), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n660), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n668), .B1(new_n675), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n830), .B2(new_n832), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n833), .A2(new_n672), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n259), .A2(new_n262), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n241), .B1(new_n240), .B2(new_n243), .ZN(new_n838));
  OAI22_X1  g637(.A1(new_n838), .A2(KEYINPUT114), .B1(new_n248), .B2(new_n251), .ZN(new_n839));
  AND2_X1   g638(.A1(new_n838), .A2(KEYINPUT114), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n257), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n265), .ZN(new_n842));
  OAI22_X1  g641(.A1(new_n836), .A2(new_n837), .B1(new_n842), .B2(new_n680), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n685), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n842), .B1(new_n613), .B2(new_n646), .ZN(new_n845));
  INV_X1    g644(.A(new_n835), .ZN(new_n846));
  NOR3_X1   g645(.A1(new_n846), .A2(new_n833), .A3(new_n672), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n828), .B1(new_n849), .B2(new_n773), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n850), .A2(new_n531), .ZN(new_n851));
  INV_X1    g650(.A(new_n705), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n375), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n423), .A3(new_n717), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n850), .A2(new_n542), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n714), .A2(new_n374), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n858), .A2(new_n696), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(G113gat), .B1(new_n860), .B2(new_n268), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT115), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n856), .B1(new_n863), .B2(new_n864), .ZN(G1340gat));
  NOR3_X1   g664(.A1(new_n860), .A2(new_n427), .A3(new_n680), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n855), .A2(new_n715), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n866), .B1(new_n427), .B2(new_n867), .ZN(G1341gat));
  NAND4_X1  g667(.A1(new_n857), .A2(G127gat), .A3(new_n645), .A4(new_n859), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n869), .B(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(KEYINPUT117), .B1(new_n854), .B2(new_n773), .ZN(new_n872));
  NOR3_X1   g671(.A1(new_n854), .A2(KEYINPUT117), .A3(new_n773), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(G127gat), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(G1342gat));
  OR4_X1    g674(.A1(KEYINPUT56), .A2(new_n854), .A3(G134gat), .A4(new_n685), .ZN(new_n876));
  OAI21_X1  g675(.A(G134gat), .B1(new_n860), .B2(new_n685), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n685), .A2(G134gat), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT56), .B1(new_n854), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n876), .A2(new_n877), .A3(new_n879), .ZN(G1343gat));
  NOR2_X1   g679(.A1(new_n758), .A2(new_n858), .ZN(new_n881));
  INV_X1    g680(.A(new_n828), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n843), .A2(new_n685), .B1(new_n845), .B2(new_n847), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n882), .B1(new_n883), .B2(new_n645), .ZN(new_n884));
  AOI21_X1  g683(.A(KEYINPUT57), .B1(new_n884), .B2(new_n542), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n542), .A2(KEYINPUT57), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n259), .A2(new_n262), .A3(new_n202), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT92), .B1(new_n264), .B2(new_n265), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n847), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n841), .A2(new_n265), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(new_n715), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n684), .B1(new_n889), .B2(new_n891), .ZN(new_n892));
  AND3_X1   g691(.A1(new_n684), .A2(new_n890), .A3(new_n847), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n773), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n886), .B1(new_n894), .B2(new_n882), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n267), .B(new_n881), .C1(new_n885), .C2(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(KEYINPUT118), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n847), .A2(new_n717), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n684), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n773), .B1(new_n899), .B2(new_n893), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n421), .B1(new_n900), .B2(new_n882), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n842), .A2(new_n680), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n902), .B1(new_n267), .B2(new_n847), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n848), .B1(new_n903), .B2(new_n684), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n828), .B1(new_n904), .B2(new_n773), .ZN(new_n905));
  OAI22_X1  g704(.A1(new_n901), .A2(KEYINPUT57), .B1(new_n905), .B2(new_n886), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT118), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n906), .A2(new_n907), .A3(new_n267), .A4(new_n881), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n897), .A2(new_n908), .A3(G141gat), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n758), .A2(new_n421), .ZN(new_n910));
  INV_X1    g709(.A(new_n910), .ZN(new_n911));
  NOR4_X1   g710(.A1(new_n850), .A2(new_n531), .A3(new_n375), .A4(new_n911), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n268), .A2(G141gat), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n914), .A2(KEYINPUT58), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n909), .A2(new_n915), .ZN(new_n916));
  INV_X1    g715(.A(new_n881), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n884), .A2(new_n542), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n894), .A2(new_n882), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n421), .A2(new_n919), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n917), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n379), .B1(new_n924), .B2(new_n717), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT58), .B1(new_n925), .B2(new_n914), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n916), .A2(new_n926), .ZN(G1344gat));
  XOR2_X1   g726(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n928));
  NAND2_X1  g727(.A1(new_n918), .A2(KEYINPUT57), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n686), .A2(new_n268), .A3(new_n683), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n894), .A2(new_n930), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n421), .A2(KEYINPUT57), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n680), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n929), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n928), .B1(new_n935), .B2(new_n381), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n715), .B(new_n881), .C1(new_n885), .C2(new_n895), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n381), .A2(KEYINPUT59), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(KEYINPUT119), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT119), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n936), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n912), .A2(new_n381), .A3(new_n715), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1345gat));
  INV_X1    g742(.A(new_n924), .ZN(new_n944));
  OAI21_X1  g743(.A(G155gat), .B1(new_n944), .B2(new_n773), .ZN(new_n945));
  INV_X1    g744(.A(G155gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n912), .A2(new_n946), .A3(new_n645), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n947), .ZN(G1346gat));
  OAI21_X1  g747(.A(G162gat), .B1(new_n944), .B2(new_n685), .ZN(new_n949));
  INV_X1    g748(.A(G162gat), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n912), .A2(new_n950), .A3(new_n684), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n949), .A2(new_n951), .ZN(G1347gat));
  NAND2_X1  g751(.A1(new_n375), .A2(new_n531), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n784), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n857), .A2(new_n954), .ZN(new_n955));
  NOR3_X1   g754(.A1(new_n955), .A2(new_n302), .A3(new_n268), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n852), .A2(new_n374), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n884), .A2(new_n531), .A3(new_n957), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT121), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n717), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n956), .B1(new_n960), .B2(new_n302), .ZN(G1348gat));
  NAND3_X1  g760(.A1(new_n959), .A2(new_n303), .A3(new_n715), .ZN(new_n962));
  OAI21_X1  g761(.A(G176gat), .B1(new_n955), .B2(new_n680), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(G1349gat));
  OAI21_X1  g763(.A(G183gat), .B1(new_n955), .B2(new_n773), .ZN(new_n965));
  INV_X1    g764(.A(new_n958), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n289), .A2(G183gat), .ZN(new_n967));
  NAND4_X1  g766(.A1(new_n966), .A2(new_n967), .A3(new_n293), .A4(new_n645), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT60), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n970), .A2(KEYINPUT122), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n969), .B(new_n971), .ZN(G1350gat));
  NAND3_X1  g771(.A1(new_n959), .A2(new_n284), .A3(new_n684), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n857), .A2(new_n684), .A3(new_n954), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT61), .ZN(new_n975));
  AND3_X1   g774(.A1(new_n974), .A2(new_n975), .A3(G190gat), .ZN(new_n976));
  AOI21_X1  g775(.A(new_n975), .B1(new_n974), .B2(G190gat), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n973), .B1(new_n976), .B2(new_n977), .ZN(G1351gat));
  NOR2_X1   g777(.A1(new_n953), .A2(new_n758), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT124), .Z(new_n980));
  NAND3_X1  g779(.A1(new_n929), .A2(new_n933), .A3(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n268), .ZN(new_n982));
  NOR3_X1   g781(.A1(new_n850), .A2(new_n714), .A3(new_n911), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(new_n375), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n837), .A2(G197gat), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AND2_X1   g785(.A1(new_n986), .A2(KEYINPUT123), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n986), .A2(KEYINPUT123), .ZN(new_n988));
  OAI21_X1  g787(.A(new_n982), .B1(new_n987), .B2(new_n988), .ZN(G1352gat));
  NAND4_X1  g788(.A1(new_n929), .A2(new_n933), .A3(new_n715), .A4(new_n980), .ZN(new_n990));
  NAND2_X1  g789(.A1(new_n990), .A2(G204gat), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n715), .A2(new_n375), .ZN(new_n992));
  AOI211_X1 g791(.A(G204gat), .B(new_n992), .C1(KEYINPUT125), .C2(KEYINPUT62), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n884), .A2(new_n531), .A3(new_n910), .A4(new_n993), .ZN(new_n994));
  NOR2_X1   g793(.A1(KEYINPUT125), .A2(KEYINPUT62), .ZN(new_n995));
  XNOR2_X1  g794(.A(new_n994), .B(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n991), .A2(new_n996), .ZN(new_n997));
  INV_X1    g796(.A(KEYINPUT126), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n991), .A2(KEYINPUT126), .A3(new_n996), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n999), .A2(new_n1000), .ZN(G1353gat));
  NOR2_X1   g800(.A1(new_n773), .A2(G211gat), .ZN(new_n1002));
  NAND3_X1  g801(.A1(new_n983), .A2(new_n375), .A3(new_n1002), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1004));
  XNOR2_X1  g803(.A(new_n1003), .B(new_n1004), .ZN(new_n1005));
  NAND4_X1  g804(.A1(new_n929), .A2(new_n933), .A3(new_n645), .A4(new_n980), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n1006), .A2(G211gat), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1007), .A2(KEYINPUT63), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT63), .ZN(new_n1009));
  NAND3_X1  g808(.A1(new_n1006), .A2(new_n1009), .A3(G211gat), .ZN(new_n1010));
  NAND3_X1  g809(.A1(new_n1005), .A2(new_n1008), .A3(new_n1010), .ZN(G1354gat));
  OAI21_X1  g810(.A(G218gat), .B1(new_n981), .B2(new_n685), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n684), .A2(new_n276), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1012), .B1(new_n984), .B2(new_n1013), .ZN(G1355gat));
endmodule


