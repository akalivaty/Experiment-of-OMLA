//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 1 1 1 0 0 1 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:35 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1291, new_n1292, new_n1294, new_n1295, new_n1296, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1362, new_n1363, new_n1364;
  NOR2_X1   g0000(.A1(G50), .A2(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  INV_X1    g0002(.A(G77), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT64), .ZN(G353));
  NOR2_X1   g0005(.A1(G97), .A2(G107), .ZN(new_n206));
  INV_X1    g0006(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  OAI21_X1  g0008(.A(G50), .B1(G58), .B2(G68), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G1), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n212), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n221));
  INV_X1    g0021(.A(G87), .ZN(new_n222));
  INV_X1    g0022(.A(G250), .ZN(new_n223));
  INV_X1    g0023(.A(G97), .ZN(new_n224));
  INV_X1    g0024(.A(G257), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT67), .Z(new_n227));
  AOI22_X1  g0027(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n228));
  INV_X1    g0028(.A(G238), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n228), .B1(new_n202), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT65), .B(G77), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n230), .B1(G244), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n227), .A2(new_n233), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n217), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI211_X1 g0036(.A(new_n214), .B(new_n220), .C1(new_n236), .C2(KEYINPUT1), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n237), .B1(KEYINPUT1), .B2(new_n236), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G250), .B(G257), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G264), .B(G270), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n243), .B(new_n246), .Z(G358));
  XNOR2_X1  g0047(.A(G68), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT68), .ZN(new_n249));
  XOR2_X1   g0049(.A(G50), .B(G58), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(G107), .B(G116), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n251), .B(new_n254), .ZN(G351));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n211), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n215), .B2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n231), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n215), .A2(G13), .A3(G20), .ZN(new_n260));
  INV_X1    g0060(.A(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n258), .A2(G77), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n231), .A2(G20), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n212), .A2(G33), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT15), .B(G87), .ZN(new_n268));
  OAI221_X1 g0068(.A(new_n263), .B1(new_n265), .B2(new_n266), .C1(new_n267), .C2(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n269), .A2(KEYINPUT73), .A3(new_n257), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(KEYINPUT73), .B1(new_n269), .B2(new_n257), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n262), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G169), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n215), .B1(G41), .B2(G45), .ZN(new_n279));
  INV_X1    g0079(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n211), .B1(G33), .B2(G41), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(new_n280), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n282), .B1(G244), .B2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n287));
  AND2_X1   g0087(.A1(KEYINPUT3), .A2(G33), .ZN(new_n288));
  NOR2_X1   g0088(.A1(KEYINPUT3), .A2(G33), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G1698), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n292), .A2(G238), .B1(G107), .B2(new_n290), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT72), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n291), .A2(G232), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n294), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT3), .ZN(new_n297));
  INV_X1    g0097(.A(G33), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g0099(.A1(KEYINPUT3), .A2(G33), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND4_X1  g0101(.A1(new_n301), .A2(KEYINPUT72), .A3(G232), .A4(new_n291), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n296), .A2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n287), .B1(new_n293), .B2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n274), .B1(new_n286), .B2(new_n304), .ZN(new_n305));
  AND2_X1   g0105(.A1(new_n273), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(G179), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n293), .A2(new_n303), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n307), .B(new_n285), .C1(new_n308), .C2(new_n287), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n272), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(new_n270), .ZN(new_n312));
  OAI211_X1 g0112(.A(G190), .B(new_n285), .C1(new_n308), .C2(new_n287), .ZN(new_n313));
  OAI21_X1  g0113(.A(G200), .B1(new_n286), .B2(new_n304), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n262), .ZN(new_n315));
  AND2_X1   g0115(.A1(new_n310), .A2(new_n315), .ZN(new_n316));
  OR2_X1    g0116(.A1(new_n316), .A2(KEYINPUT74), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n310), .A2(KEYINPUT74), .A3(new_n315), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n301), .A2(G222), .A3(new_n291), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n319), .B(KEYINPUT69), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n292), .A2(G223), .ZN(new_n321));
  OAI21_X1  g0121(.A(new_n321), .B1(new_n259), .B2(new_n301), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n283), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n282), .B1(G226), .B2(new_n284), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n274), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n212), .B1(new_n201), .B2(new_n202), .ZN(new_n327));
  INV_X1    g0127(.A(G150), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n266), .A2(new_n267), .B1(new_n328), .B2(new_n265), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n327), .B1(new_n329), .B2(KEYINPUT70), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(KEYINPUT70), .B2(new_n329), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n257), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n260), .A2(G50), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n258), .B2(G50), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n326), .B(new_n335), .C1(G179), .C2(new_n325), .ZN(new_n336));
  XNOR2_X1  g0136(.A(new_n336), .B(KEYINPUT71), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n317), .A2(new_n318), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT10), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n325), .A2(G200), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(KEYINPUT75), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(new_n335), .B(KEYINPUT9), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n323), .A2(G190), .A3(new_n324), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n342), .A2(new_n340), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  XOR2_X1   g0145(.A(new_n335), .B(KEYINPUT9), .Z(new_n346));
  NAND2_X1  g0146(.A1(new_n340), .A2(new_n344), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n341), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n345), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g0149(.A(KEYINPUT76), .B1(new_n260), .B2(G68), .ZN(new_n350));
  XOR2_X1   g0150(.A(new_n350), .B(KEYINPUT12), .Z(new_n351));
  NAND2_X1  g0151(.A1(new_n202), .A2(G20), .ZN(new_n352));
  INV_X1    g0152(.A(G50), .ZN(new_n353));
  OAI221_X1 g0153(.A(new_n352), .B1(new_n267), .B2(new_n203), .C1(new_n265), .C2(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(new_n257), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT11), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n258), .A2(G68), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n354), .A2(KEYINPUT11), .A3(new_n257), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n351), .A2(new_n357), .A3(new_n358), .A4(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT14), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT13), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n287), .A2(G238), .A3(new_n279), .ZN(new_n363));
  AND2_X1   g0163(.A1(new_n281), .A2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G226), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n291), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n240), .A2(G1698), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n366), .B(new_n367), .C1(new_n288), .C2(new_n289), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n283), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n362), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n281), .A2(new_n363), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n287), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  NOR3_X1   g0174(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT13), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n361), .B(G169), .C1(new_n372), .C2(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n364), .A2(new_n371), .A3(new_n362), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT13), .B1(new_n373), .B2(new_n374), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(G179), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n377), .A2(new_n378), .ZN(new_n381));
  AOI21_X1  g0181(.A(new_n361), .B1(new_n381), .B2(G169), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n360), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G190), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G200), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n386), .B1(new_n377), .B2(new_n378), .ZN(new_n387));
  OR3_X1    g0187(.A1(new_n385), .A2(new_n360), .A3(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n349), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n266), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n392), .A2(new_n260), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n393), .B1(new_n392), .B2(new_n258), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n257), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n299), .A2(new_n212), .A3(new_n300), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n299), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n300), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n202), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G58), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n402), .A2(new_n202), .ZN(new_n403));
  NOR2_X1   g0203(.A1(G58), .A2(G68), .ZN(new_n404));
  OAI21_X1  g0204(.A(G20), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n264), .A2(G159), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n401), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n396), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT16), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(new_n401), .B2(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n395), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n287), .A2(G232), .A3(new_n279), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n281), .A2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(new_n414), .ZN(new_n415));
  OR2_X1    g0215(.A1(G223), .A2(G1698), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n365), .A2(G1698), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n416), .B(new_n417), .C1(new_n288), .C2(new_n289), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G33), .A2(G87), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n283), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n274), .B1(new_n415), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n287), .B1(new_n418), .B2(new_n419), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n414), .A2(new_n423), .A3(new_n307), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(KEYINPUT18), .B1(new_n412), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(KEYINPUT7), .B1(new_n290), .B2(new_n212), .ZN(new_n427));
  INV_X1    g0227(.A(new_n400), .ZN(new_n428));
  OAI21_X1  g0228(.A(G68), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n407), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n429), .A2(KEYINPUT16), .A3(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n411), .A2(new_n431), .A3(new_n257), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n415), .A2(new_n421), .A3(new_n384), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n386), .B1(new_n414), .B2(new_n423), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(new_n394), .A3(new_n435), .ZN(new_n436));
  NOR2_X1   g0236(.A1(KEYINPUT77), .A2(KEYINPUT17), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n432), .A2(new_n394), .ZN(new_n439));
  INV_X1    g0239(.A(new_n425), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n439), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  XOR2_X1   g0242(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n443));
  NAND4_X1  g0243(.A1(new_n432), .A2(new_n394), .A3(new_n435), .A4(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n426), .A2(new_n438), .A3(new_n442), .A4(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n338), .A2(new_n391), .A3(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(G107), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n448), .A2(KEYINPUT6), .A3(G97), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n224), .A2(new_n448), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n450), .A2(new_n206), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n449), .B1(new_n451), .B2(KEYINPUT6), .ZN(new_n452));
  AOI22_X1  g0252(.A1(new_n452), .A2(G20), .B1(G77), .B2(new_n264), .ZN(new_n453));
  OAI21_X1  g0253(.A(G107), .B1(new_n427), .B2(new_n428), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n396), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT78), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n456), .B1(new_n298), .B2(G1), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n215), .A2(KEYINPUT78), .A3(G33), .ZN(new_n458));
  AND3_X1   g0258(.A1(new_n457), .A2(new_n458), .A3(new_n260), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT79), .B1(new_n459), .B2(new_n396), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n457), .A2(new_n458), .A3(new_n260), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT79), .ZN(new_n462));
  NOR3_X1   g0262(.A1(new_n461), .A2(new_n462), .A3(new_n257), .ZN(new_n463));
  OAI21_X1  g0263(.A(G97), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT80), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n260), .A2(new_n224), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n458), .A2(new_n260), .ZN(new_n468));
  NAND4_X1  g0268(.A1(new_n468), .A2(KEYINPUT79), .A3(new_n396), .A4(new_n457), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n462), .B1(new_n461), .B2(new_n257), .ZN(new_n470));
  AOI21_X1  g0270(.A(new_n224), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n466), .ZN(new_n472));
  OAI21_X1  g0272(.A(KEYINPUT80), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n455), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(G244), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(G1698), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n476), .B1(new_n288), .B2(new_n289), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  OAI211_X1 g0280(.A(G250), .B(G1698), .C1(new_n288), .C2(new_n289), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n476), .B(KEYINPUT4), .C1(new_n289), .C2(new_n288), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n483), .A2(new_n283), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n215), .A2(G45), .ZN(new_n485));
  OR2_X1    g0285(.A1(KEYINPUT5), .A2(G41), .ZN(new_n486));
  NAND2_X1  g0286(.A1(KEYINPUT5), .A2(G41), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n278), .ZN(new_n489));
  NOR3_X1   g0289(.A1(new_n488), .A2(new_n225), .A3(new_n283), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n484), .A2(new_n384), .A3(new_n489), .A4(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(new_n278), .ZN(new_n493));
  INV_X1    g0293(.A(G45), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G1), .ZN(new_n495));
  INV_X1    g0295(.A(new_n487), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT5), .A2(G41), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  AOI211_X1 g0299(.A(new_n499), .B(new_n490), .C1(new_n483), .C2(new_n283), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n492), .B1(new_n500), .B2(G200), .ZN(new_n501));
  AND2_X1   g0301(.A1(new_n474), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n484), .A2(new_n307), .A3(new_n489), .A4(new_n491), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n503), .B1(new_n500), .B2(G169), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n474), .A2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n225), .A2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(G250), .B2(G1698), .ZN(new_n508));
  INV_X1    g0308(.A(G294), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n508), .A2(new_n290), .B1(new_n298), .B2(new_n509), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT5), .B(G41), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n495), .B1(new_n276), .B2(new_n277), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n510), .A2(new_n283), .B1(new_n512), .B2(G264), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(G179), .A3(new_n489), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n498), .A2(G264), .A3(new_n287), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n298), .A2(new_n509), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G250), .A2(G1698), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n225), .B2(G1698), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n516), .B1(new_n518), .B2(new_n301), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n489), .B(new_n515), .C1(new_n519), .C2(new_n287), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT85), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(G169), .ZN(new_n522));
  AND2_X1   g0322(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n521), .B1(new_n520), .B2(G169), .ZN(new_n524));
  INV_X1    g0324(.A(new_n524), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n212), .B(G87), .C1(new_n288), .C2(new_n289), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT22), .ZN(new_n527));
  OR2_X1    g0327(.A1(new_n527), .A2(KEYINPUT83), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n301), .A2(new_n212), .A3(G87), .A4(new_n528), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT24), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT23), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n212), .B2(G107), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n448), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(G33), .A2(G116), .ZN(new_n538));
  INV_X1    g0338(.A(new_n538), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(KEYINPUT84), .A3(new_n212), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT84), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n538), .B2(G20), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  AND3_X1   g0343(.A1(new_n532), .A2(new_n533), .A3(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n533), .B1(new_n532), .B2(new_n543), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n257), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n469), .A2(new_n470), .A3(G107), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n260), .A2(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(new_n548), .B(KEYINPUT25), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n523), .A2(new_n525), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n520), .A2(new_n386), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n510), .A2(new_n283), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(new_n384), .A3(new_n515), .A4(new_n489), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  AND3_X1   g0356(.A1(new_n546), .A2(new_n551), .A3(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT86), .B1(new_n552), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n532), .A2(new_n543), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n532), .A2(new_n533), .A3(new_n543), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n396), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n514), .A2(new_n522), .ZN(new_n563));
  OAI22_X1  g0363(.A1(new_n562), .A2(new_n550), .B1(new_n563), .B2(new_n524), .ZN(new_n564));
  INV_X1    g0364(.A(KEYINPUT86), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n546), .A2(new_n551), .A3(new_n556), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n468), .A2(G116), .A3(new_n396), .A4(new_n457), .ZN(new_n568));
  INV_X1    g0368(.A(G116), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n261), .A2(new_n569), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n256), .A2(new_n211), .B1(G20), .B2(new_n569), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n480), .B(new_n212), .C1(G33), .C2(new_n224), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n571), .A2(KEYINPUT20), .A3(new_n572), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT20), .B1(new_n571), .B2(new_n572), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n568), .B(new_n570), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(G303), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n299), .A2(new_n576), .A3(new_n300), .ZN(new_n577));
  MUX2_X1   g0377(.A(G257), .B(G264), .S(G1698), .Z(new_n578));
  OAI211_X1 g0378(.A(new_n283), .B(new_n577), .C1(new_n578), .C2(new_n290), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n498), .A2(G270), .A3(new_n287), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n579), .A2(new_n489), .A3(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n575), .A2(G169), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT21), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AND4_X1   g0384(.A1(G179), .A2(new_n579), .A3(new_n489), .A4(new_n580), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n575), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n581), .A2(G200), .ZN(new_n587));
  OR2_X1    g0387(.A1(new_n573), .A2(new_n574), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n568), .A2(new_n570), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n579), .A2(new_n489), .A3(G190), .A4(new_n580), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n587), .A2(new_n588), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n575), .A2(KEYINPUT21), .A3(G169), .A4(new_n581), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n584), .A2(new_n586), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n223), .B1(new_n215), .B2(G45), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n278), .A2(new_n495), .B1(new_n287), .B2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(G238), .A2(G1698), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n596), .B1(new_n475), .B2(G1698), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n539), .B1(new_n597), .B2(new_n301), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n595), .B1(new_n598), .B2(new_n287), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G200), .ZN(new_n600));
  INV_X1    g0400(.A(new_n268), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n260), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT19), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n212), .B1(new_n369), .B2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n604), .B1(G87), .B2(new_n207), .ZN(new_n605));
  OAI211_X1 g0405(.A(new_n212), .B(G68), .C1(new_n288), .C2(new_n289), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n212), .A2(G33), .A3(G97), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT82), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n607), .A2(new_n608), .A3(new_n603), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n608), .B1(new_n607), .B2(new_n603), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n605), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n602), .B1(new_n611), .B2(new_n257), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n469), .A2(new_n470), .A3(G87), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n229), .A2(new_n291), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n475), .A2(G1698), .ZN(new_n615));
  OAI211_X1 g0415(.A(new_n614), .B(new_n615), .C1(new_n288), .C2(new_n289), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n538), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(new_n283), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n618), .A2(G190), .A3(new_n595), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n600), .A2(new_n612), .A3(new_n613), .A4(new_n619), .ZN(new_n620));
  AOI21_X1  g0420(.A(new_n287), .B1(new_n616), .B2(new_n538), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n287), .A2(G274), .A3(new_n495), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n594), .A2(new_n287), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g0424(.A1(new_n621), .A2(new_n624), .A3(G179), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT81), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n595), .B(new_n307), .C1(new_n598), .C2(new_n287), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT81), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n599), .A2(new_n274), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n469), .A2(new_n470), .A3(new_n601), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n612), .A2(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n620), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n593), .A2(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n506), .A2(new_n558), .A3(new_n567), .A4(new_n635), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n447), .A2(new_n636), .ZN(G372));
  AND3_X1   g0437(.A1(new_n439), .A2(new_n441), .A3(new_n440), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n441), .B1(new_n439), .B2(new_n440), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g0440(.A(new_n383), .ZN(new_n641));
  INV_X1    g0441(.A(new_n310), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n641), .B1(new_n642), .B2(new_n388), .ZN(new_n643));
  INV_X1    g0443(.A(new_n437), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n644), .B1(new_n412), .B2(new_n435), .ZN(new_n645));
  INV_X1    g0445(.A(new_n444), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n640), .B1(new_n643), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(new_n349), .ZN(new_n650));
  AND2_X1   g0450(.A1(new_n650), .A2(new_n337), .ZN(new_n651));
  INV_X1    g0451(.A(new_n504), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n467), .A2(new_n473), .ZN(new_n653));
  INV_X1    g0453(.A(new_n455), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n652), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(KEYINPUT26), .B1(new_n656), .B2(new_n634), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n625), .B1(new_n612), .B2(new_n632), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT87), .ZN(new_n659));
  AND3_X1   g0459(.A1(new_n622), .A2(new_n623), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n622), .B2(new_n623), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n618), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(new_n274), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n658), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  AND3_X1   g0465(.A1(new_n612), .A2(new_n613), .A3(new_n619), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n662), .A2(G200), .ZN(new_n667));
  AOI22_X1  g0467(.A1(new_n666), .A2(new_n667), .B1(new_n658), .B2(new_n663), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n505), .A2(new_n665), .A3(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n657), .A2(new_n664), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n592), .A2(new_n586), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n580), .A2(new_n489), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n274), .B1(new_n672), .B2(new_n579), .ZN(new_n673));
  AOI21_X1  g0473(.A(KEYINPUT21), .B1(new_n673), .B2(new_n575), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n564), .A2(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n666), .A2(new_n667), .ZN(new_n678));
  AND3_X1   g0478(.A1(new_n566), .A2(new_n678), .A3(new_n664), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n474), .A2(new_n501), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(new_n656), .A3(new_n680), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT88), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n677), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n679), .A2(KEYINPUT88), .A3(new_n656), .A4(new_n680), .ZN(new_n684));
  AOI21_X1  g0484(.A(new_n670), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n651), .B1(new_n447), .B2(new_n685), .ZN(G369));
  INV_X1    g0486(.A(new_n593), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n215), .A2(new_n212), .A3(G13), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT89), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n692), .A2(new_n694), .A3(G213), .ZN(new_n695));
  INV_X1    g0495(.A(G343), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n575), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n687), .A2(new_n698), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n699), .B1(new_n675), .B2(new_n698), .ZN(new_n700));
  XOR2_X1   g0500(.A(new_n700), .B(KEYINPUT90), .Z(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(G330), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  AND2_X1   g0503(.A1(new_n558), .A2(new_n567), .ZN(new_n704));
  OAI21_X1  g0504(.A(new_n697), .B1(new_n562), .B2(new_n550), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n552), .A2(new_n697), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(new_n697), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n552), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n675), .A2(new_n697), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n704), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n709), .A2(new_n711), .A3(new_n713), .ZN(G399));
  INV_X1    g0514(.A(new_n218), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(G41), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR3_X1   g0517(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n717), .A2(G1), .A3(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n719), .B1(new_n209), .B2(new_n717), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n721), .B(KEYINPUT28), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n668), .A2(new_n652), .A3(new_n655), .A4(KEYINPUT26), .ZN(new_n723));
  NOR3_X1   g0523(.A1(new_n634), .A2(new_n474), .A3(new_n504), .ZN(new_n724));
  OAI21_X1  g0524(.A(new_n723), .B1(new_n724), .B2(KEYINPUT26), .ZN(new_n725));
  NAND4_X1  g0525(.A1(new_n679), .A2(new_n676), .A3(new_n656), .A4(new_n680), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n725), .A2(new_n726), .A3(new_n664), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n727), .A2(new_n710), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n727), .A2(KEYINPUT94), .A3(new_n710), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT29), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n685), .B2(new_n697), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n520), .A2(new_n581), .A3(new_n307), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n490), .B1(new_n483), .B2(new_n283), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n489), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT93), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n662), .A2(new_n741), .ZN(new_n742));
  OAI211_X1 g0542(.A(new_n618), .B(KEYINPUT93), .C1(new_n660), .C2(new_n661), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n738), .A2(new_n740), .A3(new_n742), .A4(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n739), .A2(new_n585), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT92), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n621), .A2(new_n624), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n746), .B1(new_n513), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n513), .A2(new_n747), .A3(new_n746), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n745), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n744), .B1(new_n751), .B2(KEYINPUT30), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n513), .A2(new_n746), .A3(new_n747), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n739), .B(new_n585), .C1(new_n753), .C2(new_n748), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT30), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n697), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n754), .A2(new_n755), .ZN(new_n760));
  INV_X1    g0560(.A(new_n745), .ZN(new_n761));
  OAI211_X1 g0561(.A(new_n761), .B(KEYINPUT30), .C1(new_n753), .C2(new_n748), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n760), .A2(new_n762), .A3(new_n744), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n697), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n759), .B(new_n764), .C1(new_n636), .C2(new_n697), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G330), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n736), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  OAI21_X1  g0568(.A(new_n722), .B1(new_n768), .B2(G1), .ZN(G364));
  INV_X1    g0569(.A(G13), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n215), .B1(new_n771), .B2(G45), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n716), .A2(new_n773), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n703), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n701), .A2(G330), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  OR2_X1    g0581(.A1(new_n700), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n218), .A2(new_n301), .ZN(new_n783));
  INV_X1    g0583(.A(G355), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n783), .A2(new_n784), .B1(G116), .B2(new_n218), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT95), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n251), .A2(G45), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n715), .A2(new_n301), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n789), .B1(new_n494), .B2(new_n210), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n786), .B1(new_n787), .B2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n211), .B1(G20), .B2(new_n274), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n781), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n774), .B1(new_n791), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n212), .A2(new_n384), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n386), .A2(G179), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n290), .B1(new_n798), .B2(new_n576), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n212), .B1(new_n800), .B2(G190), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  AOI21_X1  g0602(.A(new_n799), .B1(G294), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n796), .A2(G179), .A3(new_n386), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n212), .A2(G190), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(new_n800), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n805), .A2(G322), .B1(new_n808), .B2(G329), .ZN(new_n809));
  NAND3_X1  g0609(.A1(new_n806), .A2(G179), .A3(new_n386), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n806), .A2(new_n797), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n811), .B1(new_n813), .B2(G283), .ZN(new_n814));
  NAND3_X1  g0614(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n815), .A2(G190), .ZN(new_n816));
  XNOR2_X1  g0616(.A(KEYINPUT33), .B(G317), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n815), .A2(new_n384), .ZN(new_n818));
  AOI22_X1  g0618(.A1(new_n816), .A2(new_n817), .B1(new_n818), .B2(G326), .ZN(new_n819));
  NAND4_X1  g0619(.A1(new_n803), .A2(new_n809), .A3(new_n814), .A4(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n811), .A2(KEYINPUT96), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n811), .A2(KEYINPUT96), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n824), .A2(new_n259), .B1(new_n402), .B2(new_n804), .ZN(new_n825));
  XNOR2_X1  g0625(.A(new_n825), .B(KEYINPUT97), .ZN(new_n826));
  INV_X1    g0626(.A(G159), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n807), .A2(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(KEYINPUT32), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n816), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n224), .B2(new_n801), .C1(new_n831), .C2(new_n202), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n301), .B1(new_n812), .B2(new_n448), .C1(new_n222), .C2(new_n798), .ZN(new_n833));
  INV_X1    g0633(.A(new_n818), .ZN(new_n834));
  OAI22_X1  g0634(.A1(new_n828), .A2(new_n829), .B1(new_n353), .B2(new_n834), .ZN(new_n835));
  OR3_X1    g0635(.A1(new_n832), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n820), .B1(new_n826), .B2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(KEYINPUT98), .ZN(new_n838));
  OR2_X1    g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n793), .B1(new_n837), .B2(new_n838), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n795), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI22_X1  g0641(.A1(new_n775), .A2(new_n777), .B1(new_n782), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(G396));
  NOR2_X1   g0643(.A1(new_n685), .A2(new_n697), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n273), .A2(new_n697), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n315), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n310), .A2(new_n846), .ZN(new_n847));
  AND4_X1   g0647(.A1(new_n309), .A2(new_n273), .A3(new_n305), .A4(new_n710), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(KEYINPUT99), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n316), .A2(new_n710), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n844), .A2(new_n851), .B1(new_n685), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n774), .B1(new_n853), .B2(new_n766), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(new_n766), .B2(new_n853), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n805), .A2(G143), .B1(G137), .B2(new_n818), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n856), .B1(new_n328), .B2(new_n831), .C1(new_n824), .C2(new_n827), .ZN(new_n857));
  XOR2_X1   g0657(.A(new_n857), .B(KEYINPUT34), .Z(new_n858));
  NOR2_X1   g0658(.A1(new_n801), .A2(new_n402), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n301), .B1(new_n798), .B2(new_n353), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n813), .A2(G68), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n862), .B2(new_n807), .ZN(new_n863));
  NOR4_X1   g0663(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(new_n798), .ZN(new_n865));
  AOI22_X1  g0665(.A1(new_n805), .A2(G294), .B1(new_n865), .B2(G107), .ZN(new_n866));
  OAI221_X1 g0666(.A(new_n866), .B1(new_n222), .B2(new_n812), .C1(new_n824), .C2(new_n569), .ZN(new_n867));
  INV_X1    g0667(.A(G311), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n290), .B1(new_n801), .B2(new_n224), .C1(new_n868), .C2(new_n807), .ZN(new_n869));
  INV_X1    g0669(.A(G283), .ZN(new_n870));
  OAI22_X1  g0670(.A1(new_n831), .A2(new_n870), .B1(new_n834), .B2(new_n576), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n867), .A2(new_n869), .A3(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n792), .B1(new_n864), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n774), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n792), .A2(new_n778), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n874), .B1(new_n203), .B2(new_n875), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n848), .B1(new_n310), .B2(new_n846), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n873), .B(new_n876), .C1(new_n779), .C2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n855), .A2(new_n878), .ZN(G384));
  NOR2_X1   g0679(.A1(new_n771), .A2(new_n215), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n733), .A2(new_n446), .A3(new_n735), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n651), .ZN(new_n882));
  XNOR2_X1  g0682(.A(new_n882), .B(KEYINPUT105), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT106), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n695), .B1(new_n638), .B2(new_n639), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n697), .A2(new_n360), .ZN(new_n886));
  AND3_X1   g0686(.A1(new_n383), .A2(new_n388), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n886), .B1(new_n383), .B2(new_n388), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n680), .B1(new_n474), .B2(new_n504), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n668), .A2(new_n566), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n682), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n893), .A2(new_n684), .A3(new_n676), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n657), .A2(new_n664), .A3(new_n669), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n852), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n890), .B1(new_n896), .B2(new_n848), .ZN(new_n897));
  OAI21_X1  g0697(.A(KEYINPUT100), .B1(new_n401), .B2(new_n407), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT100), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n429), .A2(new_n899), .A3(new_n430), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n900), .A3(new_n410), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n395), .B1(new_n901), .B2(new_n409), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n436), .B1(new_n902), .B2(new_n425), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n902), .A2(new_n695), .ZN(new_n904));
  OAI21_X1  g0704(.A(KEYINPUT37), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n425), .B1(new_n432), .B2(new_n394), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n695), .B1(new_n432), .B2(new_n394), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(KEYINPUT101), .B(KEYINPUT37), .Z(new_n910));
  NAND4_X1  g0710(.A1(new_n907), .A2(new_n909), .A3(new_n436), .A4(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n905), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n445), .A2(new_n904), .ZN(new_n913));
  AND3_X1   g0713(.A1(new_n912), .A2(KEYINPUT38), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(KEYINPUT38), .B1(new_n912), .B2(new_n913), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI211_X1 g0716(.A(KEYINPUT102), .B(new_n885), .C1(new_n897), .C2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n912), .A2(new_n913), .A3(KEYINPUT38), .ZN(new_n918));
  OAI21_X1  g0718(.A(KEYINPUT104), .B1(new_n645), .B2(new_n646), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n438), .A2(new_n920), .A3(new_n444), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n919), .A2(new_n640), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n907), .A2(new_n909), .A3(new_n436), .ZN(new_n923));
  INV_X1    g0723(.A(new_n910), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n922), .A2(new_n908), .B1(new_n911), .B2(new_n925), .ZN(new_n926));
  XOR2_X1   g0726(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n918), .B1(new_n926), .B2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT39), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n916), .A2(KEYINPUT39), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n641), .A2(new_n710), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n917), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n849), .B1(new_n685), .B2(new_n852), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT38), .ZN(new_n938));
  INV_X1    g0738(.A(new_n695), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n431), .A2(new_n257), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n429), .A2(new_n430), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT16), .B1(new_n941), .B2(KEYINPUT100), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n942), .B2(new_n900), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n939), .B1(new_n943), .B2(new_n395), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n440), .B1(new_n943), .B2(new_n395), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n944), .A2(new_n945), .A3(new_n436), .ZN(new_n946));
  INV_X1    g0746(.A(new_n436), .ZN(new_n947));
  NOR3_X1   g0747(.A1(new_n947), .A2(new_n906), .A3(new_n908), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n946), .A2(KEYINPUT37), .B1(new_n948), .B2(new_n910), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n944), .B1(new_n640), .B2(new_n647), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n938), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n918), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n937), .A2(new_n952), .A3(new_n890), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT102), .B1(new_n953), .B2(new_n885), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n936), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g0755(.A(new_n884), .B(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n877), .B1(new_n887), .B2(new_n888), .ZN(new_n957));
  INV_X1    g0757(.A(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n765), .B(new_n958), .C1(new_n914), .C2(new_n915), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT40), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT107), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n959), .A2(KEYINPUT107), .A3(new_n960), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AND3_X1   g0765(.A1(new_n765), .A2(KEYINPUT40), .A3(new_n958), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n929), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n446), .A2(new_n765), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n969), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n970), .A2(G330), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT108), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n880), .B1(new_n956), .B2(new_n973), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n974), .B1(new_n973), .B2(new_n956), .ZN(new_n975));
  OR2_X1    g0775(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n452), .A2(KEYINPUT35), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n976), .A2(G116), .A3(new_n213), .A4(new_n977), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT36), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n259), .A2(new_n209), .A3(new_n403), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n202), .A2(G50), .ZN(new_n981));
  OAI211_X1 g0781(.A(G1), .B(new_n770), .C1(new_n980), .C2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n975), .A2(new_n979), .A3(new_n982), .ZN(G367));
  OAI21_X1  g0783(.A(new_n506), .B1(new_n474), .B2(new_n710), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n505), .A2(new_n697), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n987), .A2(new_n713), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT42), .Z(new_n989));
  XNOR2_X1  g0789(.A(new_n986), .B(KEYINPUT110), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n990), .A2(new_n552), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n697), .B1(new_n991), .B2(new_n656), .ZN(new_n992));
  NOR2_X1   g0792(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n612), .A2(new_n613), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n697), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n668), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n664), .B2(new_n995), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  XNOR2_X1  g0798(.A(KEYINPUT109), .B(KEYINPUT43), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT43), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n998), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n993), .A2(new_n1002), .ZN(new_n1003));
  NOR3_X1   g0803(.A1(new_n989), .A2(new_n992), .A3(new_n1000), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n990), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n1003), .A2(new_n1004), .B1(new_n709), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n709), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n1008), .A3(new_n990), .ZN(new_n1009));
  XOR2_X1   g0809(.A(new_n716), .B(KEYINPUT41), .Z(new_n1010));
  OAI21_X1  g0810(.A(new_n713), .B1(new_n708), .B2(new_n712), .ZN(new_n1011));
  XNOR2_X1  g0811(.A(new_n702), .B(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n767), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT111), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n713), .A2(new_n986), .A3(new_n711), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT45), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1018));
  AND2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT44), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n713), .A2(new_n711), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1020), .B1(new_n1022), .B2(new_n986), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n1021), .A2(KEYINPUT44), .A3(new_n987), .ZN(new_n1024));
  AND2_X1   g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  OAI211_X1 g0825(.A(new_n1008), .B(new_n1014), .C1(new_n1019), .C2(new_n1025), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1023), .A2(new_n1024), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT111), .B1(new_n1027), .B2(new_n709), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1027), .A2(new_n709), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1013), .A2(new_n1026), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1010), .B1(new_n1030), .B2(new_n768), .ZN(new_n1031));
  OAI211_X1 g0831(.A(new_n1006), .B(new_n1009), .C1(new_n1031), .C2(new_n773), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n788), .A2(new_n246), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n794), .B1(new_n715), .B2(new_n601), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n874), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n824), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n1036), .A2(G50), .B1(G159), .B2(new_n816), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT113), .ZN(new_n1038));
  OR2_X1    g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n301), .B1(new_n798), .B2(new_n402), .ZN(new_n1040));
  INV_X1    g0840(.A(G137), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n259), .A2(new_n812), .B1(new_n807), .B2(new_n1041), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1040), .B(new_n1042), .C1(G143), .C2(new_n818), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n801), .A2(new_n202), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(G150), .B2(new_n805), .ZN(new_n1046));
  XNOR2_X1  g0846(.A(new_n1046), .B(KEYINPUT112), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1039), .A2(new_n1043), .A3(new_n1044), .A4(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1036), .A2(G283), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n798), .A2(new_n569), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n1050), .A2(KEYINPUT46), .B1(new_n868), .B2(new_n834), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT46), .B2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n812), .A2(new_n224), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n290), .B1(new_n804), .B2(new_n576), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1053), .B(new_n1054), .C1(G317), .C2(new_n808), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n802), .A2(G107), .B1(G294), .B2(new_n816), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1049), .A2(new_n1052), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1048), .A2(new_n1057), .ZN(new_n1058));
  XOR2_X1   g0858(.A(new_n1058), .B(KEYINPUT47), .Z(new_n1059));
  OAI221_X1 g0859(.A(new_n1035), .B1(new_n781), .B2(new_n997), .C1(new_n1059), .C2(new_n793), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1032), .A2(new_n1060), .ZN(G387));
  INV_X1    g0861(.A(new_n1012), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n706), .A2(new_n707), .A3(new_n780), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n783), .A2(new_n718), .B1(G107), .B2(new_n218), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n243), .A2(new_n494), .ZN(new_n1065));
  XOR2_X1   g0865(.A(new_n1065), .B(KEYINPUT114), .Z(new_n1066));
  INV_X1    g0866(.A(new_n718), .ZN(new_n1067));
  AOI211_X1 g0867(.A(G45), .B(new_n1067), .C1(G68), .C2(G77), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n266), .A2(G50), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT50), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n789), .B1(new_n1068), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1064), .B1(new_n1066), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n774), .B1(new_n1072), .B2(new_n794), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n805), .A2(G317), .B1(G311), .B2(new_n816), .ZN(new_n1074));
  INV_X1    g0874(.A(G322), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n834), .C1(new_n824), .C2(new_n576), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT48), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(new_n865), .A2(G294), .B1(new_n802), .B2(G283), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1078), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT49), .ZN(new_n1082));
  OR2_X1    g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n812), .A2(new_n569), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n301), .B(new_n1085), .C1(G326), .C2(new_n808), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  AOI211_X1 g0887(.A(new_n290), .B(new_n1053), .C1(G159), .C2(new_n818), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n259), .A2(new_n798), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G50), .B2(new_n805), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT115), .B(G150), .Z(new_n1091));
  AOI22_X1  g0891(.A1(new_n811), .A2(G68), .B1(new_n808), .B2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n801), .A2(new_n268), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(new_n816), .B2(new_n392), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1073), .B1(new_n1096), .B2(new_n792), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n1062), .A2(new_n773), .B1(new_n1063), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n768), .A2(new_n1062), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n716), .B1(new_n767), .B2(new_n1012), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(G393));
  INV_X1    g0901(.A(KEYINPUT117), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1027), .B(new_n1008), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1030), .B(new_n716), .C1(new_n1013), .C2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n788), .A2(new_n254), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n794), .B1(G97), .B2(new_n715), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n874), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n805), .A2(G311), .B1(G317), .B2(new_n818), .ZN(new_n1108));
  XOR2_X1   g0908(.A(new_n1108), .B(KEYINPUT52), .Z(new_n1109));
  OAI221_X1 g0909(.A(new_n290), .B1(new_n812), .B2(new_n448), .C1(new_n831), .C2(new_n576), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n1110), .B1(G116), .B2(new_n802), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n810), .A2(new_n509), .B1(new_n807), .B2(new_n1075), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1112), .B1(G283), .B2(new_n865), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1109), .A2(new_n1111), .A3(new_n1113), .ZN(new_n1114));
  AOI22_X1  g0914(.A1(new_n805), .A2(G159), .B1(G150), .B2(new_n818), .ZN(new_n1115));
  XNOR2_X1  g0915(.A(new_n1115), .B(KEYINPUT51), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n798), .A2(new_n202), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n301), .B1(new_n812), .B2(new_n222), .ZN(new_n1118));
  AOI211_X1 g0918(.A(new_n1117), .B(new_n1118), .C1(G143), .C2(new_n808), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n802), .A2(G77), .B1(G50), .B2(new_n816), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1119), .B(new_n1120), .C1(new_n266), .C2(new_n824), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1114), .B1(new_n1116), .B2(new_n1121), .ZN(new_n1122));
  XOR2_X1   g0922(.A(new_n1122), .B(KEYINPUT116), .Z(new_n1123));
  OAI21_X1  g0923(.A(new_n1107), .B1(new_n1123), .B2(new_n793), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1124), .B1(new_n1005), .B2(new_n780), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1103), .B2(new_n773), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1102), .B1(new_n1104), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1104), .A2(new_n1102), .A3(new_n1126), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(G390));
  NAND2_X1  g0930(.A1(new_n931), .A2(new_n932), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n778), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n805), .A2(G132), .B1(new_n808), .B2(G125), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n290), .B1(new_n813), .B2(G50), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n802), .A2(G159), .B1(G137), .B2(new_n816), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1133), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n865), .A2(new_n1091), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n1137), .A2(KEYINPUT53), .B1(new_n818), .B2(G128), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(KEYINPUT53), .B2(new_n1137), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI211_X1 g0941(.A(new_n1136), .B(new_n1139), .C1(new_n1036), .C2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n824), .A2(new_n224), .ZN(new_n1143));
  AOI22_X1  g0943(.A1(new_n802), .A2(G77), .B1(G283), .B2(new_n818), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n448), .B2(new_n831), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n290), .B1(new_n798), .B2(new_n222), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1146), .B(KEYINPUT118), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n861), .B1(new_n569), .B2(new_n804), .C1(new_n509), .C2(new_n807), .ZN(new_n1148));
  NOR4_X1   g0948(.A1(new_n1143), .A2(new_n1145), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n792), .B1(new_n1142), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n874), .B1(new_n266), .B2(new_n875), .ZN(new_n1151));
  NAND3_X1  g0951(.A1(new_n1132), .A2(new_n1150), .A3(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n730), .A2(new_n731), .A3(new_n849), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n847), .A3(new_n890), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n929), .A2(new_n933), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n897), .A2(new_n933), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1131), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NOR3_X1   g0959(.A1(new_n766), .A2(new_n850), .A3(new_n889), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1160), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1156), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1161), .A2(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1152), .B1(new_n1164), .B2(new_n772), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1153), .A2(new_n847), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n766), .ZN(new_n1167));
  AND2_X1   g0967(.A1(new_n1167), .A2(new_n851), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1162), .B(new_n1166), .C1(new_n1168), .C2(new_n890), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n890), .B1(new_n1167), .B2(new_n877), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n937), .B1(new_n1170), .B2(new_n1160), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n446), .A2(new_n1167), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n881), .A2(new_n651), .A3(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1172), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n717), .B1(new_n1164), .B2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1161), .A2(new_n1172), .A3(new_n1163), .A4(new_n1174), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1165), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(G378));
  INV_X1    g0979(.A(KEYINPUT57), .ZN(new_n1180));
  INV_X1    g0980(.A(G330), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n1181), .B1(new_n966), .B2(new_n929), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n742), .A2(new_n743), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n500), .A2(new_n737), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n754), .A2(new_n755), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n758), .B(new_n710), .C1(new_n1185), .C2(new_n762), .ZN(new_n1186));
  AOI21_X1  g0986(.A(KEYINPUT31), .B1(new_n763), .B2(new_n697), .ZN(new_n1187));
  NOR2_X1   g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n634), .ZN(new_n1189));
  AND4_X1   g0989(.A1(new_n656), .A2(new_n687), .A3(new_n1189), .A4(new_n680), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1190), .A2(new_n558), .A3(new_n567), .A4(new_n710), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n957), .B1(new_n1188), .B2(new_n1191), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n962), .B(KEYINPUT40), .C1(new_n952), .C2(new_n1192), .ZN(new_n1193));
  AOI21_X1  g0993(.A(KEYINPUT107), .B1(new_n959), .B2(new_n960), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1182), .B1(new_n1193), .B2(new_n1194), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n335), .A2(new_n939), .ZN(new_n1198));
  AND3_X1   g0998(.A1(new_n349), .A2(new_n336), .A3(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1198), .B1(new_n349), .B2(new_n336), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1197), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n349), .A2(new_n336), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1198), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n349), .A2(new_n336), .A3(new_n1198), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1204), .A2(new_n1205), .A3(new_n1196), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1201), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1195), .A2(new_n1208), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1207), .B(new_n1182), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1210));
  AND3_X1   g1010(.A1(new_n955), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n954), .ZN(new_n1212));
  AND2_X1   g1012(.A1(new_n917), .A2(new_n935), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1209), .A2(new_n1210), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n881), .A2(new_n651), .A3(new_n1173), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1156), .A2(new_n1158), .A3(new_n1162), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1162), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1216), .B1(new_n1219), .B2(new_n1172), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1180), .B1(new_n1215), .B2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1213), .A2(new_n1212), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1207), .B1(new_n965), .B2(new_n1182), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1210), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n1222), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n955), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1180), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1177), .A2(new_n1174), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n717), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1221), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT121), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n772), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1208), .A2(new_n778), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n875), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n774), .B1(G50), .B2(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(G33), .A2(G41), .ZN(new_n1236));
  INV_X1    g1036(.A(G41), .ZN(new_n1237));
  AOI211_X1 g1037(.A(G50), .B(new_n1236), .C1(new_n290), .C2(new_n1237), .ZN(new_n1238));
  NOR4_X1   g1038(.A1(new_n1089), .A2(new_n1045), .A3(G41), .A4(new_n301), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n812), .A2(new_n402), .ZN(new_n1240));
  XNOR2_X1  g1040(.A(new_n1240), .B(KEYINPUT119), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n804), .A2(new_n448), .B1(new_n807), .B2(new_n870), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(new_n601), .B2(new_n811), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(G97), .A2(new_n816), .B1(new_n818), .B2(G116), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1239), .A2(new_n1241), .A3(new_n1243), .A4(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT58), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1238), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  OAI22_X1  g1047(.A1(new_n831), .A2(new_n862), .B1(new_n801), .B2(new_n328), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(G125), .B2(new_n818), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n805), .A2(G128), .B1(new_n865), .B2(new_n1141), .ZN(new_n1250));
  OAI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(new_n1041), .C2(new_n810), .ZN(new_n1251));
  XOR2_X1   g1051(.A(new_n1251), .B(KEYINPUT120), .Z(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n808), .A2(G124), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n813), .A2(G159), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .A4(new_n1236), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1252), .A2(KEYINPUT59), .ZN(new_n1257));
  OAI221_X1 g1057(.A(new_n1247), .B1(new_n1246), .B2(new_n1245), .C1(new_n1256), .C2(new_n1257), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1235), .B1(new_n1258), .B2(new_n792), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1233), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1231), .B1(new_n1232), .B2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n773), .B1(new_n1211), .B2(new_n1214), .ZN(new_n1263));
  NAND3_X1  g1063(.A1(new_n1263), .A2(KEYINPUT121), .A3(new_n1260), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1262), .A2(new_n1264), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1230), .A2(new_n1265), .ZN(G375));
  INV_X1    g1066(.A(new_n1010), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1169), .A2(new_n1216), .A3(new_n1171), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1175), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n889), .A2(new_n778), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n774), .B1(G68), .B2(new_n1234), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G97), .A2(new_n865), .B1(new_n808), .B2(G303), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1272), .B1(new_n870), .B2(new_n804), .C1(new_n824), .C2(new_n448), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n290), .B1(new_n812), .B2(new_n203), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n831), .A2(new_n569), .B1(new_n834), .B2(new_n509), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1273), .A2(new_n1093), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  OR2_X1    g1077(.A1(new_n1277), .A2(KEYINPUT122), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(KEYINPUT122), .ZN(new_n1279));
  INV_X1    g1079(.A(G128), .ZN(new_n1280));
  OAI22_X1  g1080(.A1(new_n804), .A2(new_n1041), .B1(new_n807), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(G159), .B2(new_n865), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n301), .B1(new_n810), .B2(new_n328), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1283), .B1(G50), .B2(new_n802), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1141), .A2(new_n816), .B1(G132), .B2(new_n818), .ZN(new_n1285));
  NAND4_X1  g1085(.A1(new_n1241), .A2(new_n1282), .A3(new_n1284), .A4(new_n1285), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1278), .A2(new_n1279), .A3(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1271), .B1(new_n1287), .B2(new_n792), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(new_n1172), .A2(new_n773), .B1(new_n1270), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1269), .A2(new_n1289), .ZN(G381));
  OR4_X1    g1090(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1291));
  NOR3_X1   g1091(.A1(G390), .A2(new_n1291), .A3(G387), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1292), .A2(new_n1178), .A3(new_n1230), .A4(new_n1265), .ZN(G407));
  NAND2_X1  g1093(.A1(new_n696), .A2(G213), .ZN(new_n1294));
  XOR2_X1   g1094(.A(new_n1294), .B(KEYINPUT123), .Z(new_n1295));
  NAND2_X1  g1095(.A1(new_n1178), .A2(new_n1295), .ZN(new_n1296));
  OAI211_X1 g1096(.A(G407), .B(G213), .C1(G375), .C2(new_n1296), .ZN(G409));
  INV_X1    g1097(.A(KEYINPUT63), .ZN(new_n1298));
  INV_X1    g1098(.A(KEYINPUT124), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1230), .A2(new_n1265), .A3(G378), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1215), .A2(new_n1220), .A3(new_n1010), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1263), .A2(new_n1260), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1178), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1300), .A2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1175), .A2(KEYINPUT60), .ZN(new_n1305));
  AND2_X1   g1105(.A1(new_n1305), .A2(new_n1268), .ZN(new_n1306));
  NAND4_X1  g1106(.A1(new_n1216), .A2(KEYINPUT60), .A3(new_n1171), .A4(new_n1169), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1307), .A2(new_n716), .ZN(new_n1308));
  OAI211_X1 g1108(.A(G384), .B(new_n1289), .C1(new_n1306), .C2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(G384), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1308), .B1(new_n1305), .B2(new_n1268), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1289), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1310), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1309), .A2(new_n1313), .ZN(new_n1314));
  INV_X1    g1114(.A(new_n1314), .ZN(new_n1315));
  AND4_X1   g1115(.A1(new_n1299), .A2(new_n1304), .A3(new_n1294), .A4(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1294), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1317), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1299), .B1(new_n1318), .B2(new_n1315), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1298), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(G387), .A2(new_n1129), .A3(new_n1128), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1129), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1032), .B(new_n1060), .C1(new_n1322), .C2(new_n1127), .ZN(new_n1323));
  XNOR2_X1  g1123(.A(G393), .B(new_n842), .ZN(new_n1324));
  AND3_X1   g1124(.A1(new_n1321), .A2(new_n1323), .A3(new_n1324), .ZN(new_n1325));
  AOI21_X1  g1125(.A(new_n1324), .B1(new_n1321), .B2(new_n1323), .ZN(new_n1326));
  OR2_X1    g1126(.A1(new_n1325), .A2(new_n1326), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1309), .A2(new_n1313), .B1(G2897), .B2(new_n1295), .ZN(new_n1328));
  INV_X1    g1128(.A(G2897), .ZN(new_n1329));
  NOR2_X1   g1129(.A1(new_n1294), .A2(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1315), .B2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1331), .A2(new_n1318), .ZN(new_n1332));
  NOR3_X1   g1132(.A1(new_n1327), .A2(KEYINPUT61), .A3(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1295), .B1(new_n1300), .B2(new_n1303), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NOR3_X1   g1135(.A1(new_n1335), .A2(new_n1298), .A3(new_n1314), .ZN(new_n1336));
  AND2_X1   g1136(.A1(new_n1336), .A2(KEYINPUT125), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1336), .A2(KEYINPUT125), .ZN(new_n1338));
  OAI211_X1 g1138(.A(new_n1320), .B(new_n1333), .C1(new_n1337), .C2(new_n1338), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1331), .A2(new_n1334), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1340), .A2(KEYINPUT61), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1304), .A2(new_n1294), .A3(new_n1315), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(KEYINPUT124), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1318), .A2(new_n1299), .A3(new_n1315), .ZN(new_n1344));
  AOI21_X1  g1144(.A(KEYINPUT62), .B1(new_n1343), .B2(new_n1344), .ZN(new_n1345));
  INV_X1    g1145(.A(KEYINPUT62), .ZN(new_n1346));
  NOR2_X1   g1146(.A1(new_n1314), .A2(new_n1346), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1334), .A2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(KEYINPUT126), .ZN(new_n1349));
  INV_X1    g1149(.A(KEYINPUT126), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1334), .A2(new_n1350), .A3(new_n1347), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1349), .A2(new_n1351), .ZN(new_n1352));
  OAI211_X1 g1152(.A(KEYINPUT127), .B(new_n1341), .C1(new_n1345), .C2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1327), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1346), .B1(new_n1316), .B2(new_n1319), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1334), .A2(new_n1350), .A3(new_n1347), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1350), .B1(new_n1334), .B2(new_n1347), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1355), .A2(new_n1358), .ZN(new_n1359));
  AOI21_X1  g1159(.A(KEYINPUT127), .B1(new_n1359), .B2(new_n1341), .ZN(new_n1360));
  OAI21_X1  g1160(.A(new_n1339), .B1(new_n1354), .B2(new_n1360), .ZN(G405));
  NAND2_X1  g1161(.A1(G375), .A2(new_n1178), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n1300), .ZN(new_n1363));
  XNOR2_X1  g1163(.A(new_n1363), .B(new_n1315), .ZN(new_n1364));
  XNOR2_X1  g1164(.A(new_n1364), .B(new_n1327), .ZN(G402));
endmodule


