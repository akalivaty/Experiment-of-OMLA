//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 0 1 1 1 1 0 0 1 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 1 0 0 1 0 1 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:21:16 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n826, new_n827, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987;
  INV_X1    g000(.A(KEYINPUT35), .ZN(new_n202));
  XNOR2_X1  g001(.A(G197gat), .B(G204gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(KEYINPUT72), .B(G218gat), .ZN(new_n204));
  AND2_X1   g003(.A1(new_n204), .A2(G211gat), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n203), .B1(new_n205), .B2(KEYINPUT22), .ZN(new_n206));
  XNOR2_X1  g005(.A(G211gat), .B(G218gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G226gat), .A2(G233gat), .ZN(new_n210));
  XOR2_X1   g009(.A(new_n210), .B(KEYINPUT73), .Z(new_n211));
  XNOR2_X1  g010(.A(KEYINPUT27), .B(G183gat), .ZN(new_n212));
  INV_X1    g011(.A(G190gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OR2_X1    g013(.A1(new_n214), .A2(KEYINPUT28), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n214), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n216));
  INV_X1    g015(.A(G169gat), .ZN(new_n217));
  INV_X1    g016(.A(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OR3_X1    g018(.A1(new_n219), .A2(KEYINPUT67), .A3(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  OAI21_X1  g020(.A(KEYINPUT26), .B1(new_n219), .B2(KEYINPUT67), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  AND3_X1   g022(.A1(new_n215), .A2(new_n216), .A3(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT23), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n219), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT66), .ZN(new_n227));
  NOR2_X1   g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(KEYINPUT23), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n219), .A2(KEYINPUT66), .A3(new_n225), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n232));
  AOI21_X1  g031(.A(KEYINPUT25), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT24), .ZN(new_n234));
  INV_X1    g033(.A(G183gat), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n234), .A2(new_n235), .A3(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n235), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n213), .B1(KEYINPUT24), .B2(G183gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n231), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n233), .A2(new_n240), .ZN(new_n241));
  OAI211_X1 g040(.A(new_n231), .B(new_n239), .C1(new_n232), .C2(KEYINPUT25), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n224), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n211), .B1(new_n243), .B2(KEYINPUT29), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n241), .A2(new_n242), .ZN(new_n246));
  INV_X1    g045(.A(new_n224), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  XOR2_X1   g047(.A(new_n211), .B(KEYINPUT74), .Z(new_n249));
  AOI21_X1  g048(.A(new_n245), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n249), .ZN(new_n251));
  NOR3_X1   g050(.A1(new_n243), .A2(KEYINPUT76), .A3(new_n251), .ZN(new_n252));
  OAI211_X1 g051(.A(new_n209), .B(new_n244), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n248), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n243), .A2(new_n211), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n208), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(G8gat), .B(G36gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n258), .B(KEYINPUT77), .ZN(new_n259));
  XNOR2_X1  g058(.A(G64gat), .B(G92gat), .ZN(new_n260));
  XOR2_X1   g059(.A(new_n259), .B(new_n260), .Z(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AND3_X1   g061(.A1(new_n253), .A2(new_n257), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n262), .B1(new_n253), .B2(new_n257), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT30), .ZN(new_n265));
  NOR3_X1   g064(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n253), .A2(new_n257), .ZN(new_n267));
  NOR3_X1   g066(.A1(new_n267), .A2(KEYINPUT30), .A3(new_n261), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(G1gat), .B(G29gat), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n270), .B(KEYINPUT0), .ZN(new_n271));
  XNOR2_X1  g070(.A(G57gat), .B(G85gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT79), .B(G141gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(G148gat), .ZN(new_n277));
  OR2_X1    g076(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(KEYINPUT80), .A2(G148gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n278), .A2(G141gat), .A3(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT81), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT81), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n277), .A2(new_n283), .A3(new_n280), .ZN(new_n284));
  NAND2_X1  g083(.A1(G155gat), .A2(G162gat), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT2), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI22_X1  g088(.A1(new_n282), .A2(new_n284), .B1(new_n285), .B2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(G148gat), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n291), .A2(G141gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(G141gat), .ZN(new_n293));
  AOI21_X1  g092(.A(KEYINPUT2), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR3_X1   g093(.A1(KEYINPUT78), .A2(G155gat), .A3(G162gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT78), .B1(G155gat), .B2(G162gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n285), .ZN(new_n297));
  NOR3_X1   g096(.A1(new_n294), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n275), .B1(new_n290), .B2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n289), .A2(new_n285), .ZN(new_n300));
  INV_X1    g099(.A(new_n284), .ZN(new_n301));
  AOI21_X1  g100(.A(new_n283), .B1(new_n277), .B2(new_n280), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n298), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n303), .A2(KEYINPUT82), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(G127gat), .B(G134gat), .ZN(new_n306));
  INV_X1    g105(.A(G113gat), .ZN(new_n307));
  INV_X1    g106(.A(G120gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT1), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  AND2_X1   g108(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT68), .B(G120gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n311), .A2(G113gat), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(new_n307), .B2(new_n308), .ZN(new_n313));
  INV_X1    g112(.A(new_n306), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n310), .A2(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n299), .A2(new_n305), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT83), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n303), .A2(new_n304), .A3(new_n315), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT83), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n299), .A2(new_n305), .A3(new_n320), .A4(new_n316), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G225gat), .A2(G233gat), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n274), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n299), .A2(new_n305), .A3(KEYINPUT3), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n290), .A2(new_n298), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n326), .A2(new_n316), .A3(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n319), .B(KEYINPUT4), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n330), .A2(new_n323), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n325), .A2(new_n333), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n274), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n273), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT6), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n333), .A2(KEYINPUT5), .ZN(new_n338));
  INV_X1    g137(.A(new_n273), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n338), .B(new_n339), .C1(new_n333), .C2(new_n325), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n336), .A2(new_n337), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n322), .A2(new_n324), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(KEYINPUT5), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n335), .B1(new_n343), .B2(new_n332), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n344), .A2(KEYINPUT6), .A3(new_n339), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n269), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n248), .A2(new_n315), .ZN(new_n347));
  NAND2_X1  g146(.A1(G227gat), .A2(G233gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n348), .B(KEYINPUT64), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n243), .A2(new_n316), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT32), .ZN(new_n352));
  XNOR2_X1  g151(.A(G15gat), .B(G43gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(G71gat), .B(G99gat), .ZN(new_n354));
  XNOR2_X1  g153(.A(new_n353), .B(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n352), .B1(new_n356), .B2(KEYINPUT33), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n351), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n352), .A2(KEYINPUT33), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n351), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT69), .B1(new_n360), .B2(new_n356), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT69), .ZN(new_n362));
  AOI211_X1 g161(.A(new_n362), .B(new_n355), .C1(new_n351), .C2(new_n359), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n358), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n347), .A2(new_n350), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT34), .ZN(new_n366));
  INV_X1    g165(.A(new_n349), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n366), .B1(new_n365), .B2(new_n367), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n364), .A2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n209), .B1(new_n329), .B2(new_n254), .ZN(new_n374));
  NAND2_X1  g173(.A1(G228gat), .A2(G233gat), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n328), .B1(new_n208), .B2(KEYINPUT29), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n377), .A2(new_n299), .A3(new_n305), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n209), .A2(new_n254), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n327), .B1(new_n380), .B2(new_n328), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n375), .B1(new_n381), .B2(new_n374), .ZN(new_n382));
  XNOR2_X1  g181(.A(G78gat), .B(G106gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(KEYINPUT31), .B(G50gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT84), .ZN(new_n386));
  INV_X1    g185(.A(G22gat), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n385), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n388), .B1(new_n387), .B2(new_n385), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n379), .A2(new_n382), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n389), .B1(new_n379), .B2(new_n382), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n371), .B(new_n358), .C1(new_n361), .C2(new_n363), .ZN(new_n393));
  AND3_X1   g192(.A1(new_n373), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n202), .B1(new_n346), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n265), .B1(new_n267), .B2(new_n261), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n243), .A2(new_n211), .ZN(new_n398));
  INV_X1    g197(.A(new_n254), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n251), .B1(new_n243), .B2(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n209), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n248), .A2(new_n245), .A3(new_n249), .ZN(new_n402));
  OAI21_X1  g201(.A(KEYINPUT76), .B1(new_n243), .B2(new_n251), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT29), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n248), .A2(new_n404), .ZN(new_n405));
  AOI22_X1  g204(.A1(new_n402), .A2(new_n403), .B1(new_n405), .B2(new_n211), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n401), .B1(new_n406), .B2(new_n209), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(new_n262), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n397), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(new_n268), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n411), .A2(new_n202), .A3(new_n392), .ZN(new_n412));
  OAI21_X1  g211(.A(KEYINPUT87), .B1(new_n340), .B2(new_n337), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT87), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n344), .A2(new_n414), .A3(KEYINPUT6), .A4(new_n339), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n412), .B1(new_n341), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT71), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n373), .A2(new_n418), .A3(new_n393), .ZN(new_n419));
  OR2_X1    g218(.A1(new_n361), .A2(new_n363), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n420), .A2(KEYINPUT71), .A3(new_n371), .A4(new_n358), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(KEYINPUT88), .A3(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(KEYINPUT88), .B1(new_n419), .B2(new_n421), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n417), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n341), .A2(new_n345), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n411), .ZN(new_n427));
  INV_X1    g226(.A(new_n392), .ZN(new_n428));
  XNOR2_X1  g227(.A(KEYINPUT70), .B(KEYINPUT36), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n419), .A2(new_n429), .A3(new_n421), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n373), .A2(KEYINPUT36), .A3(new_n393), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n427), .A2(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT38), .Z(new_n433));
  INV_X1    g232(.A(KEYINPUT37), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n262), .B1(new_n407), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n267), .A2(KEYINPUT37), .ZN(new_n436));
  AOI21_X1  g235(.A(new_n433), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n253), .A2(new_n434), .A3(new_n257), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n208), .B(new_n244), .C1(new_n250), .C2(new_n252), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n209), .B1(new_n255), .B2(new_n256), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n439), .A2(KEYINPUT37), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n438), .A2(new_n441), .A3(new_n261), .A4(new_n433), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(new_n408), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n437), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n416), .A2(new_n444), .A3(new_n341), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n323), .B1(new_n330), .B2(new_n331), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT39), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n324), .B2(new_n322), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n446), .A2(new_n447), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n273), .ZN(new_n452));
  AOI211_X1 g251(.A(KEYINPUT85), .B(new_n339), .C1(new_n446), .C2(new_n447), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n449), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT40), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  OAI211_X1 g255(.A(KEYINPUT40), .B(new_n449), .C1(new_n452), .C2(new_n453), .ZN(new_n457));
  NAND4_X1  g256(.A1(new_n456), .A2(new_n340), .A3(new_n269), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n445), .A2(new_n392), .A3(new_n458), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n396), .A2(new_n425), .B1(new_n432), .B2(new_n459), .ZN(new_n460));
  XNOR2_X1  g259(.A(G15gat), .B(G22gat), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT16), .ZN(new_n462));
  AOI21_X1  g261(.A(G1gat), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n387), .A2(G15gat), .ZN(new_n464));
  INV_X1    g263(.A(G15gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(G22gat), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT89), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(G8gat), .ZN(new_n469));
  INV_X1    g268(.A(G8gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n467), .A3(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n463), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n463), .A2(new_n469), .A3(new_n471), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(G36gat), .ZN(new_n476));
  AND2_X1   g275(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n477));
  NOR2_X1   g276(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(G29gat), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n480), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(KEYINPUT15), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT15), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n479), .A2(new_n484), .A3(new_n481), .ZN(new_n485));
  XNOR2_X1  g284(.A(G43gat), .B(G50gat), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT17), .ZN(new_n488));
  INV_X1    g287(.A(new_n486), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n482), .A2(KEYINPUT15), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n487), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n488), .B1(new_n487), .B2(new_n490), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n475), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494));
  INV_X1    g293(.A(new_n474), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n495), .A2(new_n472), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n487), .A2(new_n490), .ZN(new_n497));
  AOI21_X1  g296(.A(KEYINPUT90), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND3_X1   g297(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT90), .ZN(new_n499));
  OAI211_X1 g298(.A(new_n493), .B(new_n494), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n500), .A2(KEYINPUT91), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT90), .ZN(new_n502));
  AOI211_X1 g301(.A(new_n484), .B(new_n486), .C1(new_n479), .C2(new_n481), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n489), .B1(new_n482), .B2(KEYINPUT15), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n503), .B1(new_n485), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n475), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT90), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT91), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n494), .A4(new_n493), .ZN(new_n510));
  XOR2_X1   g309(.A(KEYINPUT92), .B(KEYINPUT18), .Z(new_n511));
  NAND3_X1  g310(.A1(new_n501), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G113gat), .B(G141gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n513), .B(G197gat), .ZN(new_n514));
  XOR2_X1   g313(.A(KEYINPUT11), .B(G169gat), .Z(new_n515));
  XNOR2_X1  g314(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(new_n516), .B(KEYINPUT12), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n475), .A2(new_n505), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(new_n499), .B2(new_n498), .ZN(new_n519));
  XOR2_X1   g318(.A(new_n494), .B(KEYINPUT13), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n508), .A2(KEYINPUT18), .A3(new_n494), .A4(new_n493), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n512), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n517), .B1(new_n512), .B2(new_n523), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n460), .A2(new_n526), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n341), .A2(new_n345), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(new_n287), .ZN(new_n530));
  XNOR2_X1  g329(.A(G183gat), .B(G211gat), .ZN(new_n531));
  XOR2_X1   g330(.A(new_n530), .B(new_n531), .Z(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT21), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n535));
  NAND2_X1  g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT9), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(G57gat), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n539), .A2(G64gat), .ZN(new_n540));
  INV_X1    g339(.A(G64gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n541), .A2(G57gat), .ZN(new_n542));
  OAI211_X1 g341(.A(new_n535), .B(new_n538), .C1(new_n540), .C2(new_n542), .ZN(new_n543));
  XNOR2_X1  g342(.A(G71gat), .B(G78gat), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n541), .A2(G57gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n539), .A2(G64gat), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT93), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(new_n544), .A3(new_n538), .ZN(new_n550));
  AND3_X1   g349(.A1(new_n546), .A2(KEYINPUT94), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT94), .B1(new_n546), .B2(new_n550), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n534), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(G231gat), .A2(G233gat), .ZN(new_n554));
  OR2_X1    g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n553), .A2(new_n554), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(G127gat), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT95), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n559), .B1(new_n551), .B2(new_n552), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n546), .A2(new_n550), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT94), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n546), .A2(new_n550), .A3(KEYINPUT94), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(KEYINPUT95), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n560), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n496), .B1(new_n566), .B2(KEYINPUT21), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(G127gat), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n555), .A2(new_n569), .A3(new_n556), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n558), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n568), .B1(new_n558), .B2(new_n570), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n533), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n572), .A2(new_n573), .A3(new_n533), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(G99gat), .A2(G106gat), .ZN(new_n578));
  INV_X1    g377(.A(new_n578), .ZN(new_n579));
  NOR2_X1   g378(.A1(G99gat), .A2(G106gat), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(G85gat), .ZN(new_n582));
  INV_X1    g381(.A(G92gat), .ZN(new_n583));
  AOI22_X1  g382(.A1(KEYINPUT8), .A2(new_n578), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT7), .ZN(new_n586));
  OAI21_X1  g385(.A(KEYINPUT97), .B1(new_n586), .B2(KEYINPUT96), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT7), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G85gat), .A2(G92gat), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n592), .B1(new_n588), .B2(KEYINPUT7), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n587), .A3(new_n590), .ZN(new_n596));
  AOI211_X1 g395(.A(new_n581), .B(new_n585), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(new_n581), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n596), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n598), .B1(new_n599), .B2(new_n584), .ZN(new_n600));
  OAI22_X1  g399(.A1(new_n491), .A2(new_n492), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n600), .A2(new_n597), .ZN(new_n602));
  AND2_X1   g401(.A1(G232gat), .A2(G233gat), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n602), .A2(new_n497), .B1(KEYINPUT41), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G190gat), .B(G218gat), .Z(new_n606));
  OR2_X1    g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n606), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G134gat), .B(G162gat), .Z(new_n610));
  NOR2_X1   g409(.A1(new_n603), .A2(KEYINPUT41), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT98), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  NAND4_X1  g414(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n615), .A4(new_n608), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n577), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  OAI211_X1 g421(.A(new_n563), .B(new_n564), .C1(new_n600), .C2(new_n597), .ZN(new_n623));
  INV_X1    g422(.A(G230gat), .ZN(new_n624));
  INV_X1    g423(.A(G233gat), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  AND3_X1   g425(.A1(new_n593), .A2(new_n587), .A3(new_n590), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n593), .B1(new_n587), .B2(new_n590), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n584), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n629), .A2(new_n581), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n599), .A2(new_n598), .A3(new_n584), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n630), .A2(new_n561), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n623), .A2(new_n626), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n622), .B1(new_n634), .B2(KEYINPUT99), .ZN(new_n635));
  INV_X1    g434(.A(new_n626), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT10), .B1(new_n623), .B2(new_n632), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n630), .A2(KEYINPUT10), .A3(new_n631), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n638), .B1(new_n565), .B2(new_n560), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n636), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OAI211_X1 g439(.A(new_n635), .B(new_n640), .C1(KEYINPUT99), .C2(new_n634), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(new_n622), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n527), .A2(new_n528), .A3(new_n619), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(new_n646), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g446(.A1(new_n619), .A2(new_n645), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n460), .A2(new_n526), .A3(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(new_n649), .A2(new_n269), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT100), .B1(new_n650), .B2(new_n470), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n650), .A2(KEYINPUT100), .A3(new_n470), .ZN(new_n652));
  XOR2_X1   g451(.A(KEYINPUT16), .B(G8gat), .Z(new_n653));
  NAND2_X1  g452(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  AND2_X1   g453(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n656));
  OAI211_X1 g455(.A(new_n651), .B(new_n652), .C1(new_n655), .C2(new_n656), .ZN(G1325gat));
  NAND2_X1  g456(.A1(new_n419), .A2(new_n421), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT88), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(new_n422), .ZN(new_n661));
  AOI21_X1  g460(.A(G15gat), .B1(new_n649), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n430), .A2(new_n431), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n663), .A2(new_n465), .ZN(new_n664));
  XNOR2_X1  g463(.A(new_n664), .B(KEYINPUT101), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n662), .B1(new_n649), .B2(new_n665), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n649), .A2(new_n428), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  INV_X1    g468(.A(new_n577), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n670), .A2(new_n617), .A3(new_n644), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n527), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n673), .A2(new_n480), .A3(new_n528), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n674), .B(KEYINPUT45), .ZN(new_n675));
  XOR2_X1   g474(.A(new_n577), .B(KEYINPUT102), .Z(new_n676));
  INV_X1    g475(.A(new_n526), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(new_n677), .A3(new_n645), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n678), .B(KEYINPUT103), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT104), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n427), .A2(new_n428), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n459), .A2(new_n681), .A3(new_n663), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n395), .B1(new_n661), .B2(new_n417), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n680), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n425), .A2(new_n396), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n432), .A2(new_n459), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT104), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n617), .B(KEYINPUT105), .ZN(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n689), .A2(KEYINPUT44), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT44), .B1(new_n460), .B2(new_n617), .ZN(new_n692));
  AOI21_X1  g491(.A(new_n679), .B1(new_n691), .B2(new_n692), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n693), .A2(new_n528), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n675), .B1(new_n480), .B2(new_n694), .ZN(G1328gat));
  NOR3_X1   g494(.A1(new_n672), .A2(G36gat), .A3(new_n411), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT46), .ZN(new_n697));
  AND2_X1   g496(.A1(new_n693), .A2(new_n269), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n476), .B2(new_n698), .ZN(G1329gat));
  INV_X1    g498(.A(G43gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n663), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n700), .B1(new_n693), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT47), .ZN(new_n703));
  INV_X1    g502(.A(new_n661), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n672), .A2(G43gat), .A3(new_n704), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n702), .A2(new_n703), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n703), .B1(new_n702), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n706), .A2(new_n707), .ZN(G1330gat));
  INV_X1    g507(.A(G50gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n673), .A2(new_n709), .A3(new_n428), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n710), .A2(KEYINPUT48), .ZN(new_n711));
  AOI211_X1 g510(.A(new_n392), .B(new_n679), .C1(new_n691), .C2(new_n692), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT106), .ZN(new_n713));
  OAI21_X1  g512(.A(G50gat), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n693), .A2(new_n713), .A3(new_n428), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n711), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n710), .B1(new_n712), .B2(new_n709), .ZN(new_n717));
  INV_X1    g516(.A(KEYINPUT48), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n716), .A2(new_n719), .ZN(G1331gat));
  AND2_X1   g519(.A1(new_n684), .A2(new_n687), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n677), .A2(new_n645), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n619), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(new_n426), .ZN(new_n725));
  XNOR2_X1  g524(.A(new_n725), .B(new_n539), .ZN(G1332gat));
  NOR2_X1   g525(.A1(new_n724), .A2(new_n411), .ZN(new_n727));
  NOR2_X1   g526(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n728));
  AND2_X1   g527(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n729));
  OAI21_X1  g528(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n727), .B2(new_n728), .ZN(G1333gat));
  INV_X1    g530(.A(new_n724), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n732), .A2(G71gat), .A3(new_n701), .ZN(new_n733));
  INV_X1    g532(.A(G71gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n661), .B(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n734), .B1(new_n724), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(KEYINPUT50), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT50), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n733), .A2(new_n738), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(G1334gat));
  NAND2_X1  g542(.A1(new_n732), .A2(new_n428), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n744), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g544(.A1(new_n722), .A2(new_n577), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n746), .B1(new_n691), .B2(new_n692), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(new_n528), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n670), .A2(new_n677), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n617), .B1(new_n685), .B2(new_n686), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n750), .B2(KEYINPUT108), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n460), .A2(new_n752), .A3(new_n617), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT51), .B1(new_n751), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n750), .A2(KEYINPUT108), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n752), .B1(new_n460), .B2(new_n617), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND4_X1  g556(.A1(new_n755), .A2(new_n756), .A3(new_n757), .A4(new_n749), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n754), .A2(new_n644), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n528), .A2(new_n582), .ZN(new_n760));
  OAI22_X1  g559(.A1(new_n748), .A2(new_n582), .B1(new_n759), .B2(new_n760), .ZN(G1336gat));
  NOR2_X1   g560(.A1(new_n411), .A2(G92gat), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n754), .A2(new_n644), .A3(new_n758), .A4(new_n762), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n583), .B1(new_n747), .B2(new_n269), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT52), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT52), .ZN(new_n767));
  AND2_X1   g566(.A1(new_n747), .A2(new_n269), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n767), .B(new_n763), .C1(new_n768), .C2(new_n583), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n766), .A2(new_n769), .ZN(G1337gat));
  NAND2_X1  g569(.A1(new_n747), .A2(new_n701), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G99gat), .ZN(new_n772));
  OR2_X1    g571(.A1(new_n704), .A2(G99gat), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n759), .B2(new_n773), .ZN(G1338gat));
  NAND2_X1  g573(.A1(new_n691), .A2(new_n692), .ZN(new_n775));
  INV_X1    g574(.A(new_n746), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n428), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n777), .A2(G106gat), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n392), .A2(G106gat), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n754), .A2(new_n644), .A3(new_n758), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n781));
  AND3_X1   g580(.A1(new_n778), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g581(.A(new_n781), .B1(new_n778), .B2(new_n780), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n782), .A2(new_n783), .ZN(G1339gat));
  OR3_X1    g583(.A1(new_n637), .A2(new_n639), .A3(new_n636), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n785), .A2(KEYINPUT54), .A3(new_n640), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  OAI211_X1 g586(.A(new_n787), .B(new_n636), .C1(new_n637), .C2(new_n639), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT110), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n788), .A2(new_n789), .A3(new_n622), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n789), .B1(new_n788), .B2(new_n622), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n790), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT55), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n641), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  OAI211_X1 g595(.A(KEYINPUT111), .B(new_n641), .C1(new_n792), .C2(new_n793), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n792), .A2(new_n793), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n796), .A2(new_n677), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n512), .A2(new_n523), .A3(new_n517), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n519), .A2(new_n520), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n494), .B1(new_n508), .B2(new_n493), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n516), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n800), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n644), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n688), .B1(new_n799), .B2(new_n805), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n794), .A2(new_n795), .B1(new_n793), .B2(new_n792), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n688), .A3(new_n804), .A4(new_n797), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n676), .B1(new_n806), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n648), .A2(new_n677), .ZN(new_n811));
  INV_X1    g610(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n428), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n528), .A2(new_n411), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n704), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n816), .A2(new_n307), .A3(new_n526), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n810), .A2(new_n812), .ZN(new_n818));
  AND3_X1   g617(.A1(new_n818), .A2(new_n528), .A3(new_n394), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n819), .A2(new_n677), .A3(new_n411), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n817), .B1(new_n820), .B2(new_n307), .ZN(G1340gat));
  OAI21_X1  g620(.A(G120gat), .B1(new_n816), .B2(new_n645), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n411), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n645), .A2(new_n311), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(G1341gat));
  OAI21_X1  g624(.A(G127gat), .B1(new_n816), .B2(new_n676), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n670), .A2(new_n569), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n826), .B1(new_n823), .B2(new_n827), .ZN(G1342gat));
  NOR3_X1   g627(.A1(new_n269), .A2(G134gat), .A3(new_n617), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n819), .A2(new_n829), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n816), .B2(new_n617), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(KEYINPUT56), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n831), .A2(new_n832), .A3(new_n833), .ZN(G1343gat));
  INV_X1    g633(.A(KEYINPUT58), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n701), .A2(new_n814), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT113), .ZN(new_n837));
  AND2_X1   g636(.A1(new_n804), .A2(new_n644), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n793), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT112), .B1(new_n792), .B2(new_n793), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n794), .A2(new_n526), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n808), .B1(new_n843), .B2(new_n618), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n811), .B1(new_n844), .B2(new_n577), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n392), .A2(new_n846), .ZN(new_n847));
  INV_X1    g646(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n837), .B1(new_n845), .B2(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT112), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n798), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n792), .A2(KEYINPUT112), .A3(new_n793), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI221_X1 g652(.A(new_n641), .B1(new_n792), .B2(new_n793), .C1(new_n525), .C2(new_n524), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n805), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n617), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n670), .B1(new_n856), .B2(new_n808), .ZN(new_n857));
  OAI211_X1 g656(.A(KEYINPUT113), .B(new_n847), .C1(new_n857), .C2(new_n811), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n849), .A2(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT57), .B1(new_n818), .B2(new_n428), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n677), .B(new_n836), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(new_n276), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n663), .A2(new_n428), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT114), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n663), .A2(KEYINPUT114), .A3(new_n428), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n818), .A2(new_n528), .A3(new_n866), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT116), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n426), .B1(new_n810), .B2(new_n812), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n871), .A2(KEYINPUT116), .A3(new_n866), .A4(new_n867), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n526), .A2(G141gat), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n870), .A2(new_n411), .A3(new_n872), .A4(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT117), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n874), .A2(new_n875), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n835), .B(new_n863), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT115), .ZN(new_n879));
  INV_X1    g678(.A(new_n873), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n868), .A2(new_n269), .A3(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n863), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n879), .B1(new_n883), .B2(KEYINPUT58), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n881), .B1(new_n861), .B2(new_n862), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n885), .A2(KEYINPUT115), .A3(new_n835), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n878), .B1(new_n884), .B2(new_n886), .ZN(G1344gat));
  XOR2_X1   g686(.A(KEYINPUT118), .B(KEYINPUT59), .Z(new_n888));
  NOR2_X1   g687(.A1(new_n843), .A2(new_n618), .ZN(new_n889));
  AND4_X1   g688(.A1(new_n618), .A2(new_n807), .A3(new_n804), .A4(new_n797), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n577), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(new_n812), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n892), .A2(new_n428), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n893), .A2(new_n846), .B1(new_n818), .B2(new_n847), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n836), .A2(new_n644), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT119), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n291), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(KEYINPUT119), .B1(new_n894), .B2(new_n895), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n888), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n278), .A2(new_n279), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n836), .B1(new_n859), .B2(new_n860), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  AOI211_X1 g702(.A(KEYINPUT59), .B(new_n901), .C1(new_n903), .C2(new_n644), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n870), .A2(new_n872), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n411), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n644), .A2(new_n901), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n900), .A2(new_n904), .B1(new_n907), .B2(new_n908), .ZN(G1345gat));
  NAND3_X1  g708(.A1(new_n906), .A2(new_n411), .A3(new_n670), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n676), .A2(new_n287), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT120), .ZN(new_n912));
  AOI22_X1  g711(.A1(new_n910), .A2(new_n287), .B1(new_n903), .B2(new_n912), .ZN(G1346gat));
  OAI21_X1  g712(.A(G162gat), .B1(new_n902), .B2(new_n689), .ZN(new_n914));
  NAND3_X1  g713(.A1(new_n411), .A2(new_n288), .A3(new_n618), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n914), .B1(new_n905), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(KEYINPUT121), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT121), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n914), .B(new_n918), .C1(new_n905), .C2(new_n915), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n917), .A2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n528), .A2(new_n411), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n394), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n818), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(G169gat), .B1(new_n924), .B2(new_n677), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n736), .A2(new_n921), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(new_n813), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n526), .A2(new_n217), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n925), .B1(new_n928), .B2(new_n929), .ZN(G1348gat));
  OAI21_X1  g729(.A(G176gat), .B1(new_n927), .B2(new_n645), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n924), .A2(new_n218), .A3(new_n644), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(G1349gat));
  OAI21_X1  g732(.A(G183gat), .B1(new_n927), .B2(new_n676), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n924), .A2(new_n212), .A3(new_n670), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g735(.A(new_n936), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n924), .A2(new_n213), .A3(new_n688), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n928), .A2(new_n618), .ZN(new_n940));
  AOI21_X1  g739(.A(new_n939), .B1(new_n940), .B2(G190gat), .ZN(new_n941));
  AOI211_X1 g740(.A(KEYINPUT61), .B(new_n213), .C1(new_n928), .C2(new_n618), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1351gat));
  INV_X1    g742(.A(KEYINPUT125), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n921), .A2(new_n663), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT124), .ZN(new_n946));
  OR2_X1    g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n944), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  AND2_X1   g748(.A1(new_n945), .A2(new_n946), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n945), .A2(new_n946), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n950), .A2(new_n951), .A3(KEYINPUT125), .ZN(new_n952));
  NOR3_X1   g751(.A1(new_n894), .A2(new_n949), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n953), .A2(new_n677), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(G197gat), .ZN(new_n955));
  INV_X1    g754(.A(KEYINPUT123), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n392), .B1(new_n810), .B2(new_n812), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(new_n945), .ZN(new_n958));
  INV_X1    g757(.A(KEYINPUT122), .ZN(new_n959));
  XNOR2_X1  g758(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n526), .A2(G197gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n956), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n960), .A2(new_n956), .A3(new_n961), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n955), .B1(new_n962), .B2(new_n963), .ZN(G1352gat));
  INV_X1    g763(.A(G204gat), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n952), .A2(new_n949), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n893), .A2(new_n846), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n818), .A2(new_n847), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(new_n644), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n965), .B1(new_n970), .B2(KEYINPUT126), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n971), .B1(KEYINPUT126), .B2(new_n970), .ZN(new_n972));
  NOR3_X1   g771(.A1(new_n958), .A2(G204gat), .A3(new_n645), .ZN(new_n973));
  XNOR2_X1  g772(.A(new_n973), .B(KEYINPUT62), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n972), .A2(new_n974), .ZN(G1353gat));
  INV_X1    g774(.A(G211gat), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n976), .A3(new_n670), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n670), .B1(new_n950), .B2(new_n951), .ZN(new_n978));
  OAI21_X1  g777(.A(G211gat), .B1(new_n894), .B2(new_n978), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT63), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n979), .A2(new_n980), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n977), .B1(new_n981), .B2(new_n982), .ZN(G1354gat));
  AOI21_X1  g782(.A(G218gat), .B1(new_n960), .B2(new_n688), .ZN(new_n984));
  OR2_X1    g783(.A1(new_n953), .A2(KEYINPUT127), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n618), .A2(new_n204), .ZN(new_n986));
  AOI21_X1  g785(.A(new_n986), .B1(new_n953), .B2(KEYINPUT127), .ZN(new_n987));
  AOI21_X1  g786(.A(new_n984), .B1(new_n985), .B2(new_n987), .ZN(G1355gat));
endmodule


