

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728;

  XNOR2_X1 U366 ( .A(n509), .B(KEYINPUT104), .ZN(n728) );
  NOR2_X1 U367 ( .A1(n534), .A2(n366), .ZN(n359) );
  XNOR2_X1 U368 ( .A(n568), .B(KEYINPUT1), .ZN(n535) );
  NOR2_X1 U369 ( .A1(G953), .A2(G237), .ZN(n440) );
  NOR2_X2 U370 ( .A1(n628), .A2(n627), .ZN(n717) );
  XNOR2_X1 U371 ( .A(KEYINPUT38), .B(n621), .ZN(n577) );
  XNOR2_X1 U372 ( .A(n352), .B(n349), .ZN(n496) );
  XNOR2_X1 U373 ( .A(n357), .B(KEYINPUT41), .ZN(n565) );
  NOR2_X1 U374 ( .A1(n486), .A2(n494), .ZN(n357) );
  XNOR2_X1 U375 ( .A(n590), .B(n497), .ZN(n599) );
  INV_X1 U376 ( .A(n496), .ZN(n621) );
  OR2_X1 U377 ( .A1(n680), .A2(n643), .ZN(n352) );
  INV_X1 U378 ( .A(n380), .ZN(n424) );
  XOR2_X1 U379 ( .A(G122), .B(G107), .Z(n464) );
  INV_X1 U380 ( .A(KEYINPUT64), .ZN(n378) );
  XNOR2_X1 U381 ( .A(KEYINPUT65), .B(KEYINPUT4), .ZN(n395) );
  XNOR2_X1 U382 ( .A(G146), .B(G125), .ZN(n380) );
  XOR2_X1 U383 ( .A(G119), .B(G110), .Z(n432) );
  XNOR2_X1 U384 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U385 ( .A(G143), .B(G122), .ZN(n450) );
  NAND2_X1 U386 ( .A1(n684), .A2(G475), .ZN(n356) );
  INV_X1 U387 ( .A(KEYINPUT83), .ZN(n374) );
  OR2_X1 U388 ( .A1(n722), .A2(n546), .ZN(n543) );
  NAND2_X1 U389 ( .A1(n496), .A2(n616), .ZN(n590) );
  XNOR2_X1 U390 ( .A(n424), .B(n368), .ZN(n712) );
  XNOR2_X1 U391 ( .A(G140), .B(KEYINPUT10), .ZN(n368) );
  XNOR2_X1 U392 ( .A(G128), .B(KEYINPUT23), .ZN(n381) );
  INV_X1 U393 ( .A(KEYINPUT8), .ZN(n370) );
  XNOR2_X1 U394 ( .A(n461), .B(n347), .ZN(n365) );
  OR2_X1 U395 ( .A1(n480), .A2(n536), .ZN(n421) );
  AND2_X1 U396 ( .A1(n576), .A2(n575), .ZN(n595) );
  XNOR2_X1 U397 ( .A(n456), .B(n455), .ZN(n521) );
  XNOR2_X1 U398 ( .A(n454), .B(G475), .ZN(n455) );
  XNOR2_X1 U399 ( .A(n389), .B(n346), .ZN(n390) );
  NAND2_X1 U400 ( .A1(n373), .A2(n642), .ZN(n372) );
  NAND2_X1 U401 ( .A1(n684), .A2(G210), .ZN(n363) );
  NAND2_X1 U402 ( .A1(n595), .A2(n376), .ZN(n375) );
  NOR2_X1 U403 ( .A1(n348), .A2(n621), .ZN(n376) );
  XNOR2_X1 U404 ( .A(n375), .B(n374), .ZN(n597) );
  XNOR2_X1 U405 ( .A(n582), .B(KEYINPUT87), .ZN(n583) );
  XOR2_X1 U406 ( .A(G113), .B(G119), .Z(n410) );
  XOR2_X1 U407 ( .A(G113), .B(G104), .Z(n442) );
  XOR2_X1 U408 ( .A(KEYINPUT66), .B(G101), .Z(n413) );
  NAND2_X1 U409 ( .A1(G234), .A2(G237), .ZN(n469) );
  NOR2_X1 U410 ( .A1(G902), .A2(G237), .ZN(n438) );
  XNOR2_X1 U411 ( .A(n358), .B(KEYINPUT108), .ZN(n486) );
  NAND2_X1 U412 ( .A1(n577), .A2(n616), .ZN(n358) );
  INV_X1 U413 ( .A(KEYINPUT74), .ZN(n571) );
  NAND2_X1 U414 ( .A1(n717), .A2(n641), .ZN(n373) );
  XNOR2_X1 U415 ( .A(G110), .B(G104), .ZN(n401) );
  XNOR2_X1 U416 ( .A(n437), .B(n697), .ZN(n680) );
  INV_X1 U417 ( .A(KEYINPUT19), .ZN(n497) );
  NAND2_X1 U418 ( .A1(n366), .A2(n470), .ZN(n394) );
  XNOR2_X1 U419 ( .A(n386), .B(n367), .ZN(n694) );
  XNOR2_X1 U420 ( .A(n369), .B(n712), .ZN(n367) );
  XNOR2_X1 U421 ( .A(n364), .B(n458), .ZN(n646) );
  XNOR2_X1 U422 ( .A(n365), .B(n465), .ZN(n364) );
  NOR2_X1 U423 ( .A1(n565), .A2(n600), .ZN(n566) );
  XNOR2_X1 U424 ( .A(n592), .B(n591), .ZN(n593) );
  XNOR2_X1 U425 ( .A(KEYINPUT109), .B(KEYINPUT36), .ZN(n591) );
  OR2_X1 U426 ( .A1(n522), .A2(n348), .ZN(n524) );
  AND2_X1 U427 ( .A1(n359), .A2(n377), .ZN(n509) );
  INV_X1 U428 ( .A(KEYINPUT60), .ZN(n353) );
  XNOR2_X1 U429 ( .A(n356), .B(n351), .ZN(n355) );
  INV_X1 U430 ( .A(KEYINPUT56), .ZN(n360) );
  XNOR2_X1 U431 ( .A(n363), .B(n683), .ZN(n362) );
  INV_X1 U432 ( .A(n375), .ZN(n669) );
  XOR2_X1 U433 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n346) );
  XNOR2_X1 U434 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n347) );
  NAND2_X1 U435 ( .A1(n521), .A2(n520), .ZN(n348) );
  AND2_X1 U436 ( .A1(G210), .A2(n439), .ZN(n349) );
  NOR2_X1 U437 ( .A1(n646), .A2(G902), .ZN(n350) );
  XOR2_X1 U438 ( .A(n692), .B(n691), .Z(n351) );
  NAND2_X1 U439 ( .A1(n362), .A2(n654), .ZN(n361) );
  NAND2_X1 U440 ( .A1(n355), .A2(n654), .ZN(n354) );
  NAND2_X1 U441 ( .A1(n625), .A2(n641), .ZN(n644) );
  AND2_X2 U442 ( .A1(n644), .A2(n643), .ZN(n371) );
  XNOR2_X1 U443 ( .A(n354), .B(n353), .ZN(G60) );
  NAND2_X1 U444 ( .A1(n359), .A2(n510), .ZN(n512) );
  XNOR2_X1 U445 ( .A(n361), .B(n360), .ZN(G51) );
  NOR2_X1 U446 ( .A1(n366), .A2(n554), .ZN(n560) );
  NOR2_X1 U447 ( .A1(n366), .A2(n470), .ZN(n472) );
  NAND2_X1 U448 ( .A1(n618), .A2(n366), .ZN(n537) );
  XNOR2_X2 U449 ( .A(n391), .B(n390), .ZN(n366) );
  NAND2_X1 U450 ( .A1(n457), .A2(G221), .ZN(n369) );
  XNOR2_X2 U451 ( .A(n379), .B(n370), .ZN(n457) );
  AND2_X4 U452 ( .A1(n372), .A2(n371), .ZN(n684) );
  OR2_X1 U453 ( .A1(n718), .A2(G952), .ZN(n654) );
  NOR2_X1 U454 ( .A1(n535), .A2(n573), .ZN(n377) );
  INV_X1 U455 ( .A(KEYINPUT46), .ZN(n582) );
  INV_X1 U456 ( .A(KEYINPUT68), .ZN(n607) );
  BUF_X1 U457 ( .A(n641), .Z(n705) );
  XNOR2_X1 U458 ( .A(n404), .B(n403), .ZN(n405) );
  AND2_X1 U459 ( .A1(n535), .A2(n536), .ZN(n510) );
  XNOR2_X1 U460 ( .A(n640), .B(n639), .ZN(G75) );
  XNOR2_X2 U461 ( .A(n378), .B(G953), .ZN(n718) );
  NAND2_X1 U462 ( .A1(n718), .A2(G234), .ZN(n379) );
  XNOR2_X1 U463 ( .A(n432), .B(n381), .ZN(n385) );
  XOR2_X1 U464 ( .A(KEYINPUT24), .B(KEYINPUT76), .Z(n383) );
  XNOR2_X1 U465 ( .A(G137), .B(KEYINPUT84), .ZN(n382) );
  XNOR2_X1 U466 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U467 ( .A(n385), .B(n384), .Z(n386) );
  NOR2_X1 U468 ( .A1(n694), .A2(G902), .ZN(n391) );
  INV_X1 U469 ( .A(G902), .ZN(n406) );
  XNOR2_X1 U470 ( .A(n406), .B(KEYINPUT15), .ZN(n643) );
  INV_X1 U471 ( .A(n643), .ZN(n387) );
  NAND2_X1 U472 ( .A1(G234), .A2(n387), .ZN(n388) );
  XNOR2_X1 U473 ( .A(KEYINPUT20), .B(n388), .ZN(n392) );
  NAND2_X1 U474 ( .A1(n392), .A2(G217), .ZN(n389) );
  NAND2_X1 U475 ( .A1(G221), .A2(n392), .ZN(n393) );
  XNOR2_X1 U476 ( .A(n393), .B(KEYINPUT21), .ZN(n554) );
  INV_X1 U477 ( .A(n554), .ZN(n470) );
  XNOR2_X2 U478 ( .A(n394), .B(KEYINPUT67), .ZN(n570) );
  XNOR2_X2 U479 ( .A(G143), .B(G128), .ZN(n462) );
  XNOR2_X1 U480 ( .A(n462), .B(n395), .ZN(n425) );
  XNOR2_X1 U481 ( .A(G134), .B(G131), .ZN(n397) );
  INV_X1 U482 ( .A(G137), .ZN(n396) );
  XNOR2_X1 U483 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U484 ( .A(n425), .B(n398), .ZN(n711) );
  XNOR2_X1 U485 ( .A(n711), .B(G146), .ZN(n417) );
  XOR2_X1 U486 ( .A(G140), .B(G107), .Z(n400) );
  AND2_X1 U487 ( .A1(n718), .A2(G227), .ZN(n399) );
  XNOR2_X1 U488 ( .A(n400), .B(n399), .ZN(n404) );
  XNOR2_X1 U489 ( .A(n413), .B(KEYINPUT70), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n401), .B(KEYINPUT77), .ZN(n402) );
  XNOR2_X1 U491 ( .A(n427), .B(n402), .ZN(n403) );
  XNOR2_X1 U492 ( .A(n417), .B(n405), .ZN(n687) );
  NAND2_X1 U493 ( .A1(n687), .A2(n406), .ZN(n407) );
  XNOR2_X2 U494 ( .A(n407), .B(G469), .ZN(n568) );
  NAND2_X1 U495 ( .A1(n570), .A2(n535), .ZN(n408) );
  XNOR2_X1 U496 ( .A(n408), .B(KEYINPUT72), .ZN(n480) );
  NAND2_X1 U497 ( .A1(n440), .A2(G210), .ZN(n409) );
  XNOR2_X1 U498 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U499 ( .A(n411), .B(KEYINPUT5), .Z(n415) );
  XNOR2_X1 U500 ( .A(G116), .B(KEYINPUT69), .ZN(n412) );
  XNOR2_X1 U501 ( .A(n412), .B(KEYINPUT3), .ZN(n436) );
  XNOR2_X1 U502 ( .A(n436), .B(n413), .ZN(n414) );
  XNOR2_X1 U503 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U504 ( .A(n417), .B(n416), .ZN(n651) );
  OR2_X1 U505 ( .A1(n651), .A2(G902), .ZN(n418) );
  XNOR2_X1 U506 ( .A(n418), .B(G472), .ZN(n573) );
  XNOR2_X1 U507 ( .A(n573), .B(KEYINPUT6), .ZN(n536) );
  INV_X1 U508 ( .A(KEYINPUT91), .ZN(n419) );
  XNOR2_X1 U509 ( .A(n419), .B(KEYINPUT33), .ZN(n420) );
  XNOR2_X2 U510 ( .A(n421), .B(n420), .ZN(n517) );
  INV_X1 U511 ( .A(n517), .ZN(n467) );
  XOR2_X1 U512 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n423) );
  NAND2_X1 U513 ( .A1(G224), .A2(n718), .ZN(n422) );
  XNOR2_X1 U514 ( .A(n423), .B(n422), .ZN(n431) );
  XNOR2_X1 U515 ( .A(n424), .B(KEYINPUT92), .ZN(n426) );
  XNOR2_X1 U516 ( .A(n426), .B(n425), .ZN(n429) );
  INV_X1 U517 ( .A(n427), .ZN(n428) );
  XNOR2_X1 U518 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U519 ( .A(n431), .B(n430), .ZN(n437) );
  XOR2_X1 U520 ( .A(n442), .B(KEYINPUT16), .Z(n434) );
  XNOR2_X1 U521 ( .A(n432), .B(n464), .ZN(n433) );
  XNOR2_X1 U522 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U523 ( .A(n436), .B(n435), .ZN(n697) );
  XNOR2_X1 U524 ( .A(n438), .B(KEYINPUT73), .ZN(n439) );
  NAND2_X1 U525 ( .A1(G214), .A2(n439), .ZN(n616) );
  NAND2_X1 U526 ( .A1(G214), .A2(n440), .ZN(n441) );
  XNOR2_X1 U527 ( .A(n441), .B(n712), .ZN(n443) );
  XOR2_X1 U528 ( .A(n443), .B(n442), .Z(n453) );
  XOR2_X1 U529 ( .A(KEYINPUT11), .B(KEYINPUT97), .Z(n445) );
  XNOR2_X1 U530 ( .A(G131), .B(KEYINPUT98), .ZN(n444) );
  XNOR2_X1 U531 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U532 ( .A(KEYINPUT99), .B(KEYINPUT96), .Z(n447) );
  XNOR2_X1 U533 ( .A(KEYINPUT12), .B(KEYINPUT95), .ZN(n446) );
  XNOR2_X1 U534 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U535 ( .A(n449), .B(n448), .Z(n451) );
  XNOR2_X1 U536 ( .A(n453), .B(n452), .ZN(n692) );
  NOR2_X1 U537 ( .A1(G902), .A2(n692), .ZN(n456) );
  XNOR2_X1 U538 ( .A(KEYINPUT100), .B(KEYINPUT13), .ZN(n454) );
  INV_X1 U539 ( .A(n521), .ZN(n466) );
  NAND2_X1 U540 ( .A1(G217), .A2(n457), .ZN(n458) );
  XOR2_X1 U541 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n460) );
  XNOR2_X1 U542 ( .A(G116), .B(G134), .ZN(n459) );
  XNOR2_X1 U543 ( .A(n460), .B(n459), .ZN(n461) );
  INV_X1 U544 ( .A(n462), .ZN(n463) );
  XNOR2_X1 U545 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U546 ( .A(n350), .B(G478), .ZN(n519) );
  NAND2_X1 U547 ( .A1(n466), .A2(n519), .ZN(n494) );
  NOR2_X1 U548 ( .A1(n467), .A2(n565), .ZN(n468) );
  NOR2_X1 U549 ( .A1(n468), .A2(G953), .ZN(n636) );
  XNOR2_X1 U550 ( .A(n469), .B(KEYINPUT14), .ZN(n499) );
  NAND2_X1 U551 ( .A1(G952), .A2(n499), .ZN(n498) );
  XNOR2_X1 U552 ( .A(KEYINPUT49), .B(KEYINPUT114), .ZN(n471) );
  XNOR2_X1 U553 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U554 ( .A(KEYINPUT115), .B(n473), .Z(n477) );
  NOR2_X1 U555 ( .A1(n570), .A2(n535), .ZN(n474) );
  XOR2_X1 U556 ( .A(KEYINPUT116), .B(n474), .Z(n475) );
  XNOR2_X1 U557 ( .A(KEYINPUT50), .B(n475), .ZN(n476) );
  NAND2_X1 U558 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U559 ( .A1(n573), .A2(n478), .ZN(n479) );
  XNOR2_X1 U560 ( .A(KEYINPUT117), .B(n479), .ZN(n481) );
  INV_X1 U561 ( .A(n573), .ZN(n561) );
  OR2_X1 U562 ( .A1(n480), .A2(n561), .ZN(n527) );
  NAND2_X1 U563 ( .A1(n481), .A2(n527), .ZN(n482) );
  XNOR2_X1 U564 ( .A(n482), .B(KEYINPUT51), .ZN(n483) );
  XNOR2_X1 U565 ( .A(n483), .B(KEYINPUT118), .ZN(n484) );
  NOR2_X1 U566 ( .A1(n565), .A2(n484), .ZN(n491) );
  NOR2_X1 U567 ( .A1(n577), .A2(n616), .ZN(n485) );
  NOR2_X1 U568 ( .A1(n494), .A2(n485), .ZN(n488) );
  NOR2_X1 U569 ( .A1(n519), .A2(n521), .ZN(n665) );
  NAND2_X1 U570 ( .A1(n519), .A2(n521), .ZN(n673) );
  INV_X1 U571 ( .A(n673), .ZN(n670) );
  NOR2_X1 U572 ( .A1(n665), .A2(n670), .ZN(n601) );
  NOR2_X1 U573 ( .A1(n486), .A2(n601), .ZN(n487) );
  OR2_X1 U574 ( .A1(n488), .A2(n487), .ZN(n489) );
  AND2_X1 U575 ( .A1(n517), .A2(n489), .ZN(n490) );
  NOR2_X1 U576 ( .A1(n491), .A2(n490), .ZN(n492) );
  XNOR2_X1 U577 ( .A(n492), .B(KEYINPUT52), .ZN(n493) );
  NOR2_X1 U578 ( .A1(n498), .A2(n493), .ZN(n634) );
  NOR2_X1 U579 ( .A1(n554), .A2(n494), .ZN(n495) );
  XNOR2_X1 U580 ( .A(KEYINPUT103), .B(n495), .ZN(n506) );
  NOR2_X1 U581 ( .A1(G953), .A2(n498), .ZN(n558) );
  NAND2_X1 U582 ( .A1(n499), .A2(G902), .ZN(n500) );
  XNOR2_X1 U583 ( .A(KEYINPUT94), .B(n500), .ZN(n555) );
  INV_X1 U584 ( .A(G953), .ZN(n704) );
  NOR2_X1 U585 ( .A1(n704), .A2(G898), .ZN(n501) );
  XNOR2_X1 U586 ( .A(n501), .B(KEYINPUT93), .ZN(n698) );
  NOR2_X1 U587 ( .A1(n555), .A2(n698), .ZN(n502) );
  NOR2_X1 U588 ( .A1(n558), .A2(n502), .ZN(n503) );
  NOR2_X2 U589 ( .A1(n599), .A2(n503), .ZN(n505) );
  INV_X1 U590 ( .A(KEYINPUT0), .ZN(n504) );
  XNOR2_X2 U591 ( .A(n505), .B(n504), .ZN(n531) );
  NOR2_X1 U592 ( .A1(n506), .A2(n531), .ZN(n508) );
  XNOR2_X1 U593 ( .A(KEYINPUT71), .B(KEYINPUT22), .ZN(n507) );
  XNOR2_X1 U594 ( .A(n508), .B(n507), .ZN(n534) );
  INV_X1 U595 ( .A(n728), .ZN(n514) );
  XOR2_X1 U596 ( .A(KEYINPUT78), .B(KEYINPUT32), .Z(n511) );
  XNOR2_X1 U597 ( .A(n512), .B(n511), .ZN(n722) );
  NOR2_X1 U598 ( .A1(n722), .A2(KEYINPUT44), .ZN(n513) );
  NAND2_X1 U599 ( .A1(n514), .A2(n513), .ZN(n515) );
  INV_X1 U600 ( .A(KEYINPUT89), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n515), .A2(n547), .ZN(n526) );
  INV_X1 U602 ( .A(n531), .ZN(n516) );
  NAND2_X1 U603 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U604 ( .A(n518), .B(KEYINPUT34), .ZN(n522) );
  INV_X1 U605 ( .A(n519), .ZN(n520) );
  XNOR2_X1 U606 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n523) );
  XNOR2_X2 U607 ( .A(n524), .B(n523), .ZN(n649) );
  INV_X1 U608 ( .A(n649), .ZN(n525) );
  NAND2_X1 U609 ( .A1(n526), .A2(n525), .ZN(n542) );
  NOR2_X1 U610 ( .A1(n527), .A2(n531), .ZN(n528) );
  XNOR2_X1 U611 ( .A(n528), .B(KEYINPUT31), .ZN(n675) );
  AND2_X1 U612 ( .A1(n561), .A2(n568), .ZN(n529) );
  NAND2_X1 U613 ( .A1(n570), .A2(n529), .ZN(n530) );
  OR2_X1 U614 ( .A1(n531), .A2(n530), .ZN(n662) );
  NAND2_X1 U615 ( .A1(n675), .A2(n662), .ZN(n533) );
  INV_X1 U616 ( .A(n601), .ZN(n532) );
  NAND2_X1 U617 ( .A1(n533), .A2(n532), .ZN(n540) );
  INV_X1 U618 ( .A(n534), .ZN(n539) );
  INV_X1 U619 ( .A(n535), .ZN(n618) );
  INV_X1 U620 ( .A(n536), .ZN(n587) );
  NOR2_X1 U621 ( .A1(n537), .A2(n587), .ZN(n538) );
  NAND2_X1 U622 ( .A1(n539), .A2(n538), .ZN(n658) );
  AND2_X1 U623 ( .A1(n540), .A2(n658), .ZN(n541) );
  AND2_X1 U624 ( .A1(n542), .A2(n541), .ZN(n551) );
  NAND2_X1 U625 ( .A1(n649), .A2(n547), .ZN(n545) );
  INV_X1 U626 ( .A(KEYINPUT44), .ZN(n546) );
  NOR2_X1 U627 ( .A1(n728), .A2(n543), .ZN(n544) );
  NAND2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n549) );
  NAND2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U630 ( .A1(n549), .A2(n548), .ZN(n550) );
  NAND2_X1 U631 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X2 U632 ( .A(n552), .B(KEYINPUT45), .ZN(n641) );
  NOR2_X1 U633 ( .A1(n705), .A2(KEYINPUT2), .ZN(n553) );
  XNOR2_X1 U634 ( .A(n553), .B(KEYINPUT85), .ZN(n632) );
  INV_X1 U635 ( .A(KEYINPUT48), .ZN(n612) );
  XOR2_X1 U636 ( .A(KEYINPUT106), .B(KEYINPUT28), .Z(n563) );
  OR2_X1 U637 ( .A1(n555), .A2(n718), .ZN(n556) );
  NOR2_X1 U638 ( .A1(G900), .A2(n556), .ZN(n557) );
  NOR2_X1 U639 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U640 ( .A(KEYINPUT79), .B(n559), .ZN(n567) );
  NAND2_X1 U641 ( .A1(n560), .A2(n567), .ZN(n585) );
  OR2_X1 U642 ( .A1(n585), .A2(n561), .ZN(n562) );
  XNOR2_X1 U643 ( .A(n563), .B(n562), .ZN(n564) );
  NAND2_X1 U644 ( .A1(n564), .A2(n568), .ZN(n600) );
  XOR2_X1 U645 ( .A(KEYINPUT42), .B(n566), .Z(n725) );
  AND2_X1 U646 ( .A1(n568), .A2(n567), .ZN(n569) );
  NAND2_X1 U647 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U648 ( .A(n572), .B(n571), .ZN(n576) );
  NAND2_X1 U649 ( .A1(n573), .A2(n616), .ZN(n574) );
  XOR2_X1 U650 ( .A(KEYINPUT30), .B(n574), .Z(n575) );
  NAND2_X1 U651 ( .A1(n595), .A2(n577), .ZN(n579) );
  XOR2_X1 U652 ( .A(KEYINPUT88), .B(KEYINPUT39), .Z(n578) );
  XOR2_X1 U653 ( .A(n579), .B(n578), .Z(n613) );
  AND2_X1 U654 ( .A1(n613), .A2(n670), .ZN(n581) );
  XNOR2_X1 U655 ( .A(KEYINPUT107), .B(KEYINPUT40), .ZN(n580) );
  XNOR2_X1 U656 ( .A(n581), .B(n580), .ZN(n727) );
  NAND2_X1 U657 ( .A1(n725), .A2(n727), .ZN(n584) );
  XNOR2_X1 U658 ( .A(n584), .B(n583), .ZN(n610) );
  INV_X1 U659 ( .A(KEYINPUT105), .ZN(n589) );
  NOR2_X1 U660 ( .A1(n585), .A2(n673), .ZN(n586) );
  NAND2_X1 U661 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U662 ( .A(n589), .B(n588), .ZN(n615) );
  NOR2_X1 U663 ( .A1(n615), .A2(n590), .ZN(n592) );
  NOR2_X1 U664 ( .A1(n593), .A2(n618), .ZN(n594) );
  XNOR2_X1 U665 ( .A(n594), .B(KEYINPUT110), .ZN(n723) );
  NAND2_X1 U666 ( .A1(KEYINPUT47), .A2(n601), .ZN(n596) );
  NAND2_X1 U667 ( .A1(n597), .A2(n596), .ZN(n598) );
  XNOR2_X1 U668 ( .A(KEYINPUT81), .B(n598), .ZN(n605) );
  NOR2_X1 U669 ( .A1(n600), .A2(n599), .ZN(n671) );
  XOR2_X1 U670 ( .A(n671), .B(KEYINPUT47), .Z(n603) );
  NAND2_X1 U671 ( .A1(n671), .A2(n601), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n606) );
  NOR2_X1 U674 ( .A1(n723), .A2(n606), .ZN(n608) );
  XNOR2_X1 U675 ( .A(n608), .B(n607), .ZN(n609) );
  NOR2_X1 U676 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U677 ( .A(n612), .B(n611), .ZN(n628) );
  NAND2_X1 U678 ( .A1(n665), .A2(n613), .ZN(n678) );
  NAND2_X1 U679 ( .A1(n678), .A2(KEYINPUT2), .ZN(n614) );
  XOR2_X1 U680 ( .A(n614), .B(KEYINPUT80), .Z(n623) );
  INV_X1 U681 ( .A(n615), .ZN(n617) );
  AND2_X1 U682 ( .A1(n617), .A2(n616), .ZN(n619) );
  NAND2_X1 U683 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U684 ( .A(n620), .B(KEYINPUT43), .ZN(n622) );
  AND2_X1 U685 ( .A1(n622), .A2(n621), .ZN(n679) );
  INV_X1 U686 ( .A(n679), .ZN(n626) );
  NAND2_X1 U687 ( .A1(n623), .A2(n626), .ZN(n624) );
  NOR2_X1 U688 ( .A1(n628), .A2(n624), .ZN(n625) );
  INV_X1 U689 ( .A(n644), .ZN(n630) );
  NAND2_X1 U690 ( .A1(n626), .A2(n678), .ZN(n627) );
  NOR2_X1 U691 ( .A1(KEYINPUT2), .A2(n717), .ZN(n629) );
  NOR2_X1 U692 ( .A1(n630), .A2(n629), .ZN(n631) );
  AND2_X1 U693 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U694 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U695 ( .A1(n636), .A2(n635), .ZN(n640) );
  XOR2_X1 U696 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n638) );
  INV_X1 U697 ( .A(KEYINPUT119), .ZN(n637) );
  XNOR2_X1 U698 ( .A(n638), .B(n637), .ZN(n639) );
  INV_X1 U699 ( .A(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U700 ( .A1(n684), .A2(G478), .ZN(n645) );
  XNOR2_X1 U701 ( .A(n645), .B(KEYINPUT122), .ZN(n647) );
  XNOR2_X1 U702 ( .A(n647), .B(n646), .ZN(n648) );
  INV_X1 U703 ( .A(n654), .ZN(n696) );
  NOR2_X1 U704 ( .A1(n648), .A2(n696), .ZN(G63) );
  XOR2_X1 U705 ( .A(G122), .B(n649), .Z(G24) );
  NAND2_X1 U706 ( .A1(n684), .A2(G472), .ZN(n653) );
  XNOR2_X1 U707 ( .A(KEYINPUT111), .B(KEYINPUT62), .ZN(n650) );
  XNOR2_X1 U708 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U709 ( .A(n653), .B(n652), .ZN(n655) );
  NAND2_X1 U710 ( .A1(n655), .A2(n654), .ZN(n657) );
  XNOR2_X1 U711 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n656) );
  XNOR2_X1 U712 ( .A(n657), .B(n656), .ZN(G57) );
  XNOR2_X1 U713 ( .A(G101), .B(n658), .ZN(G3) );
  NOR2_X1 U714 ( .A1(n673), .A2(n662), .ZN(n659) );
  XOR2_X1 U715 ( .A(G104), .B(n659), .Z(G6) );
  XOR2_X1 U716 ( .A(KEYINPUT27), .B(KEYINPUT112), .Z(n661) );
  XNOR2_X1 U717 ( .A(G107), .B(KEYINPUT26), .ZN(n660) );
  XNOR2_X1 U718 ( .A(n661), .B(n660), .ZN(n664) );
  INV_X1 U719 ( .A(n665), .ZN(n676) );
  NOR2_X1 U720 ( .A1(n676), .A2(n662), .ZN(n663) );
  XOR2_X1 U721 ( .A(n664), .B(n663), .Z(G9) );
  XOR2_X1 U722 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n667) );
  NAND2_X1 U723 ( .A1(n671), .A2(n665), .ZN(n666) );
  XNOR2_X1 U724 ( .A(n667), .B(n666), .ZN(n668) );
  XOR2_X1 U725 ( .A(G128), .B(n668), .Z(G30) );
  XOR2_X1 U726 ( .A(G143), .B(n669), .Z(G45) );
  NAND2_X1 U727 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U728 ( .A(n672), .B(G146), .ZN(G48) );
  NOR2_X1 U729 ( .A1(n673), .A2(n675), .ZN(n674) );
  XOR2_X1 U730 ( .A(G113), .B(n674), .Z(G15) );
  NOR2_X1 U731 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U732 ( .A(G116), .B(n677), .Z(G18) );
  XNOR2_X1 U733 ( .A(G134), .B(n678), .ZN(G36) );
  XOR2_X1 U734 ( .A(G140), .B(n679), .Z(G42) );
  XNOR2_X1 U735 ( .A(KEYINPUT55), .B(KEYINPUT82), .ZN(n682) );
  XNOR2_X1 U736 ( .A(n680), .B(KEYINPUT54), .ZN(n681) );
  XNOR2_X1 U737 ( .A(n682), .B(n681), .ZN(n683) );
  NAND2_X1 U738 ( .A1(n684), .A2(G469), .ZN(n689) );
  XOR2_X1 U739 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n685) );
  XNOR2_X1 U740 ( .A(n685), .B(KEYINPUT121), .ZN(n686) );
  XNOR2_X1 U741 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U742 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U743 ( .A1(n696), .A2(n690), .ZN(G54) );
  INV_X1 U744 ( .A(KEYINPUT59), .ZN(n691) );
  NAND2_X1 U745 ( .A1(n684), .A2(G217), .ZN(n693) );
  XNOR2_X1 U746 ( .A(n694), .B(n693), .ZN(n695) );
  NOR2_X1 U747 ( .A1(n696), .A2(n695), .ZN(G66) );
  XNOR2_X1 U748 ( .A(n697), .B(G101), .ZN(n699) );
  NAND2_X1 U749 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U750 ( .A(n700), .B(KEYINPUT125), .ZN(n710) );
  NAND2_X1 U751 ( .A1(G953), .A2(G224), .ZN(n701) );
  XNOR2_X1 U752 ( .A(KEYINPUT61), .B(n701), .ZN(n702) );
  NAND2_X1 U753 ( .A1(n702), .A2(G898), .ZN(n703) );
  XNOR2_X1 U754 ( .A(KEYINPUT123), .B(n703), .ZN(n708) );
  NAND2_X1 U755 ( .A1(n705), .A2(n704), .ZN(n706) );
  XOR2_X1 U756 ( .A(KEYINPUT124), .B(n706), .Z(n707) );
  NOR2_X1 U757 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U758 ( .A(n710), .B(n709), .Z(G69) );
  XOR2_X1 U759 ( .A(n712), .B(n711), .Z(n716) );
  XOR2_X1 U760 ( .A(n716), .B(G227), .Z(n713) );
  NAND2_X1 U761 ( .A1(n713), .A2(G900), .ZN(n714) );
  XNOR2_X1 U762 ( .A(n714), .B(KEYINPUT126), .ZN(n715) );
  NAND2_X1 U763 ( .A1(n715), .A2(G953), .ZN(n721) );
  XNOR2_X1 U764 ( .A(n717), .B(n716), .ZN(n719) );
  NAND2_X1 U765 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U766 ( .A1(n721), .A2(n720), .ZN(G72) );
  XOR2_X1 U767 ( .A(G119), .B(n722), .Z(G21) );
  XNOR2_X1 U768 ( .A(G125), .B(KEYINPUT37), .ZN(n724) );
  XNOR2_X1 U769 ( .A(n724), .B(n723), .ZN(G27) );
  XOR2_X1 U770 ( .A(G137), .B(n725), .Z(n726) );
  XNOR2_X1 U771 ( .A(KEYINPUT127), .B(n726), .ZN(G39) );
  XNOR2_X1 U772 ( .A(G131), .B(n727), .ZN(G33) );
  XOR2_X1 U773 ( .A(n728), .B(G110), .Z(G12) );
endmodule

