//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:10 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n551,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n606, new_n607, new_n608, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT65), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT66), .Z(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(G125), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n468), .A2(G2105), .ZN(new_n469));
  AND2_X1   g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n463), .A2(G2105), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n470), .B1(new_n471), .B2(G137), .ZN(new_n472));
  AND2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  MUX2_X1   g048(.A(G100), .B(G112), .S(G2105), .Z(new_n474));
  AOI22_X1  g049(.A1(new_n471), .A2(G136), .B1(G2104), .B2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(KEYINPUT3), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(new_n468), .ZN(new_n477));
  NAND2_X1  g052(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT67), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n479), .A2(new_n480), .A3(G2105), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n480), .B1(new_n479), .B2(G2105), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G124), .ZN(new_n485));
  OAI21_X1  g060(.A(new_n475), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XOR2_X1   g061(.A(new_n486), .B(KEYINPUT68), .Z(G162));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n488), .B1(new_n477), .B2(new_n478), .ZN(new_n489));
  AND2_X1   g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  OAI21_X1  g065(.A(G2105), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G2105), .ZN(new_n492));
  NAND2_X1  g067(.A1(KEYINPUT4), .A2(G138), .ZN(new_n493));
  AOI21_X1  g068(.A(new_n493), .B1(new_n477), .B2(new_n478), .ZN(new_n494));
  NAND2_X1  g069(.A1(G102), .A2(G2104), .ZN(new_n495));
  INV_X1    g070(.A(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n492), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  OAI211_X1 g072(.A(G138), .B(new_n492), .C1(new_n461), .C2(new_n462), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n491), .A2(new_n497), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT69), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n491), .A2(new_n497), .A3(new_n503), .A4(new_n500), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(G164));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  OR2_X1    g082(.A1(KEYINPUT5), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g085(.A1(new_n510), .A2(G62), .ZN(new_n511));
  OR2_X1    g086(.A1(new_n511), .A2(KEYINPUT71), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT72), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n514), .B1(new_n511), .B2(KEYINPUT71), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n507), .B1(new_n512), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(G50), .ZN(new_n517));
  NAND2_X1  g092(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n518));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n507), .A2(KEYINPUT6), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n520), .A2(new_n510), .A3(new_n521), .ZN(new_n523));
  INV_X1    g098(.A(G88), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n517), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n516), .A2(new_n525), .ZN(G166));
  NAND4_X1  g101(.A1(new_n520), .A2(G51), .A3(G543), .A4(new_n521), .ZN(new_n527));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  OR2_X1    g103(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(KEYINPUT7), .ZN(new_n530));
  AND2_X1   g105(.A1(G63), .A2(G651), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n529), .A2(new_n530), .B1(new_n510), .B2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G89), .ZN(new_n533));
  OAI211_X1 g108(.A(new_n527), .B(new_n532), .C1(new_n523), .C2(new_n533), .ZN(G286));
  INV_X1    g109(.A(G286), .ZN(G168));
  INV_X1    g110(.A(new_n523), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G90), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n520), .A2(G543), .A3(new_n521), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G52), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n510), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n540), .A2(new_n507), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n537), .A2(new_n539), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  AOI22_X1  g118(.A1(new_n510), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n507), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT73), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n536), .A2(G81), .B1(new_n538), .B2(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g123(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(G153));
  AND3_X1   g125(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G36), .ZN(G176));
  NAND2_X1  g127(.A1(G1), .A2(G3), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT8), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n551), .A2(new_n554), .ZN(G188));
  INV_X1    g130(.A(KEYINPUT9), .ZN(new_n556));
  NAND3_X1  g131(.A1(new_n538), .A2(new_n556), .A3(G53), .ZN(new_n557));
  INV_X1    g132(.A(G53), .ZN(new_n558));
  OAI21_X1  g133(.A(KEYINPUT9), .B1(new_n522), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(new_n510), .ZN(new_n562));
  INV_X1    g137(.A(G65), .ZN(new_n563));
  OAI21_X1  g138(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n536), .A2(G91), .B1(G651), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n560), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G166), .ZN(G303));
  NAND4_X1  g142(.A1(new_n520), .A2(G87), .A3(new_n510), .A4(new_n521), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n520), .A2(G49), .A3(G543), .A4(new_n521), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n570), .A2(KEYINPUT74), .ZN(new_n571));
  NOR2_X1   g146(.A1(new_n570), .A2(KEYINPUT74), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n568), .B(new_n569), .C1(new_n571), .C2(new_n572), .ZN(G288));
  NAND2_X1  g148(.A1(G73), .A2(G543), .ZN(new_n574));
  INV_X1    g149(.A(G61), .ZN(new_n575));
  OAI21_X1  g150(.A(new_n574), .B1(new_n562), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(G651), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n520), .A2(G86), .A3(new_n510), .A4(new_n521), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n520), .A2(G48), .A3(G543), .A4(new_n521), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(G305));
  INV_X1    g155(.A(G47), .ZN(new_n581));
  INV_X1    g156(.A(G85), .ZN(new_n582));
  OAI22_X1  g157(.A1(new_n581), .A2(new_n522), .B1(new_n523), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT75), .ZN(new_n584));
  AND2_X1   g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g160(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n585), .A2(new_n586), .B1(new_n507), .B2(new_n587), .ZN(G290));
  INV_X1    g163(.A(G868), .ZN(new_n589));
  NOR2_X1   g164(.A1(G301), .A2(new_n589), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n536), .A2(G92), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT10), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n562), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n538), .A2(G54), .B1(G651), .B2(new_n595), .ZN(new_n596));
  AND2_X1   g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g172(.A(new_n590), .B1(new_n597), .B2(new_n589), .ZN(G284));
  AOI21_X1  g173(.A(new_n590), .B1(new_n597), .B2(new_n589), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  XNOR2_X1  g175(.A(G299), .B(KEYINPUT76), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(G148));
  NAND3_X1  g180(.A1(new_n597), .A2(new_n604), .A3(G868), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n549), .A2(new_n589), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(KEYINPUT11), .Z(G282));
  INV_X1    g184(.A(new_n608), .ZN(G323));
  NAND2_X1  g185(.A1(new_n471), .A2(G2104), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT12), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT13), .Z(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(new_n614));
  XOR2_X1   g189(.A(KEYINPUT77), .B(G2100), .Z(new_n615));
  NOR2_X1   g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n616), .B(KEYINPUT78), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n614), .A2(new_n615), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT79), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n471), .A2(G135), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT80), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n621), .A2(new_n492), .A3(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n492), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n623), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n620), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(new_n484), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n625), .B1(new_n626), .B2(G123), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n617), .A2(new_n619), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(KEYINPUT15), .B(G2435), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT81), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2430), .ZN(new_n633));
  OR2_X1    g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n632), .A2(new_n633), .ZN(new_n635));
  NAND3_X1  g210(.A1(new_n634), .A2(KEYINPUT14), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT82), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2451), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT16), .ZN(new_n639));
  XNOR2_X1  g214(.A(G2443), .B(G2446), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n637), .B(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G1341), .B(G1348), .Z(new_n643));
  NOR2_X1   g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT84), .Z(new_n645));
  NAND2_X1  g220(.A1(new_n642), .A2(new_n643), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT83), .ZN(new_n647));
  AND3_X1   g222(.A1(new_n645), .A2(G14), .A3(new_n647), .ZN(G401));
  XOR2_X1   g223(.A(G2084), .B(G2090), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G2072), .B(G2078), .Z(new_n651));
  XNOR2_X1  g226(.A(G2067), .B(G2678), .ZN(new_n652));
  INV_X1    g227(.A(new_n652), .ZN(new_n653));
  NOR3_X1   g228(.A1(new_n650), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT18), .ZN(new_n655));
  INV_X1    g230(.A(new_n651), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n656), .A2(KEYINPUT17), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n652), .B1(new_n658), .B2(new_n649), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(new_n650), .B2(new_n657), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n650), .A2(new_n653), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n656), .B1(new_n661), .B2(KEYINPUT17), .ZN(new_n662));
  OAI21_X1  g237(.A(new_n655), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(G2096), .Z(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(G2100), .ZN(G227));
  XOR2_X1   g240(.A(G1971), .B(G1976), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT19), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g245(.A1(new_n668), .A2(new_n669), .ZN(new_n671));
  NOR3_X1   g246(.A1(new_n667), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT20), .Z(new_n674));
  AOI211_X1 g249(.A(new_n672), .B(new_n674), .C1(new_n667), .C2(new_n671), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1991), .B(G1996), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n677), .B(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n682), .A2(G5), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G171), .B2(new_n682), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n684), .A2(G1961), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(KEYINPUT97), .ZN(new_n686));
  OR2_X1    g261(.A1(KEYINPUT30), .A2(G28), .ZN(new_n687));
  NAND2_X1  g262(.A1(KEYINPUT30), .A2(G28), .ZN(new_n688));
  AOI21_X1  g263(.A(G29), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT31), .B(G11), .Z(new_n690));
  AOI211_X1 g265(.A(new_n689), .B(new_n690), .C1(new_n627), .C2(G29), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n691), .B(KEYINPUT96), .Z(new_n692));
  INV_X1    g267(.A(G29), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n693), .A2(G26), .ZN(new_n694));
  XOR2_X1   g269(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  MUX2_X1   g270(.A(G104), .B(G116), .S(G2105), .Z(new_n696));
  AOI22_X1  g271(.A1(new_n471), .A2(G140), .B1(G2104), .B2(new_n696), .ZN(new_n697));
  INV_X1    g272(.A(G128), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n697), .B1(new_n484), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n695), .B1(new_n699), .B2(G29), .ZN(new_n700));
  INV_X1    g275(.A(G2067), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n692), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT24), .B(G34), .Z(new_n704));
  NOR2_X1   g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(G160), .B2(G29), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G2084), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n684), .A2(G1961), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT27), .B(G1996), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n709), .B(KEYINPUT94), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n693), .A2(G32), .ZN(new_n711));
  AOI22_X1  g286(.A1(new_n471), .A2(G141), .B1(G105), .B2(new_n469), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT26), .Z(new_n714));
  NAND2_X1  g289(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n715), .B1(new_n626), .B2(G129), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n711), .B1(new_n716), .B2(new_n693), .ZN(new_n717));
  AOI211_X1 g292(.A(new_n707), .B(new_n708), .C1(new_n710), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n682), .A2(G21), .ZN(new_n719));
  OAI21_X1  g294(.A(new_n719), .B1(G168), .B2(new_n682), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(G1966), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n682), .A2(G20), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT23), .Z(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(G299), .B2(G16), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT100), .B(G1956), .Z(new_n725));
  AOI21_X1  g300(.A(new_n721), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  AND4_X1   g301(.A1(new_n686), .A2(new_n703), .A3(new_n718), .A4(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n693), .A2(G27), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n693), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT99), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT98), .B(G2078), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G4), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(new_n597), .B2(G16), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT90), .B(G1348), .Z(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n734), .A2(new_n736), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n724), .A2(new_n725), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n737), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n693), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n693), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(KEYINPUT29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G2090), .ZN(new_n744));
  NAND4_X1  g319(.A1(new_n727), .A2(new_n732), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  INV_X1    g320(.A(KEYINPUT101), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n682), .A2(G19), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT91), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n748), .B1(new_n548), .B2(G16), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1341), .Z(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G33), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(KEYINPUT93), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n471), .A2(G139), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n469), .A2(G103), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n479), .A2(G127), .ZN(new_n758));
  NAND2_X1  g333(.A1(G115), .A2(G2104), .ZN(new_n759));
  AND2_X1   g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n754), .B(new_n757), .C1(new_n760), .C2(new_n492), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n753), .B1(new_n761), .B2(new_n693), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(G2072), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n706), .A2(G2084), .ZN(new_n764));
  OAI211_X1 g339(.A(new_n763), .B(new_n764), .C1(new_n710), .C2(new_n717), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT95), .ZN(new_n766));
  OAI211_X1 g341(.A(new_n751), .B(new_n766), .C1(new_n743), .C2(G2090), .ZN(new_n767));
  OR3_X1    g342(.A1(new_n745), .A2(new_n746), .A3(new_n767), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n746), .B1(new_n745), .B2(new_n767), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT36), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n471), .A2(G131), .ZN(new_n772));
  AND2_X1   g347(.A1(G107), .A2(G2105), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G95), .B2(new_n492), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n772), .B1(new_n468), .B2(new_n774), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n626), .B2(G119), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(G29), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G25), .B2(G29), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT35), .B(G1991), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(new_n780), .ZN(new_n781));
  OR2_X1    g356(.A1(G16), .A2(G23), .ZN(new_n782));
  NAND2_X1  g357(.A1(G288), .A2(KEYINPUT87), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n570), .B(KEYINPUT74), .ZN(new_n784));
  INV_X1    g359(.A(KEYINPUT87), .ZN(new_n785));
  NAND4_X1  g360(.A1(new_n784), .A2(new_n785), .A3(new_n568), .A4(new_n569), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n783), .A2(new_n786), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n782), .B1(new_n787), .B2(new_n682), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT33), .B(G1976), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n788), .B(new_n789), .Z(new_n790));
  NOR2_X1   g365(.A1(G6), .A2(G16), .ZN(new_n791));
  AND3_X1   g366(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(G16), .ZN(new_n793));
  XOR2_X1   g368(.A(KEYINPUT32), .B(G1981), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n682), .A2(G22), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(KEYINPUT88), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n797), .B1(G303), .B2(G16), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G1971), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n790), .A2(new_n795), .A3(new_n799), .ZN(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT86), .B(KEYINPUT34), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n781), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g377(.A(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT89), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n682), .A2(G24), .ZN(new_n805));
  INV_X1    g380(.A(KEYINPUT85), .ZN(new_n806));
  XNOR2_X1  g381(.A(G290), .B(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n805), .B1(new_n807), .B2(new_n682), .ZN(new_n808));
  INV_X1    g383(.A(G1986), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n810), .A2(new_n811), .B1(new_n800), .B2(new_n801), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n803), .A2(new_n804), .A3(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n804), .B1(new_n803), .B2(new_n812), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n771), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n815), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n817), .A2(KEYINPUT36), .A3(new_n813), .ZN(new_n818));
  AND3_X1   g393(.A1(new_n770), .A2(new_n816), .A3(new_n818), .ZN(G311));
  NAND3_X1  g394(.A1(new_n816), .A2(new_n770), .A3(new_n818), .ZN(G150));
  NAND2_X1  g395(.A1(new_n597), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT38), .ZN(new_n822));
  AOI22_X1  g397(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n823));
  NOR2_X1   g398(.A1(new_n823), .A2(new_n507), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n536), .B2(G93), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n538), .A2(G55), .ZN(new_n826));
  NAND3_X1  g401(.A1(new_n825), .A2(KEYINPUT102), .A3(new_n826), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n548), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n825), .A2(new_n826), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT102), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n831), .A2(new_n548), .A3(new_n827), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n828), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n822), .B(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(KEYINPUT39), .ZN(new_n835));
  AOI21_X1  g410(.A(G860), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n829), .A2(G860), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(KEYINPUT37), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT103), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n837), .A2(KEYINPUT103), .A3(new_n839), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(G145));
  INV_X1    g419(.A(G37), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n776), .B(new_n612), .ZN(new_n846));
  MUX2_X1   g421(.A(G106), .B(G118), .S(G2105), .Z(new_n847));
  AOI22_X1  g422(.A1(new_n471), .A2(G142), .B1(G2104), .B2(new_n847), .ZN(new_n848));
  INV_X1    g423(.A(G130), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n484), .B2(new_n849), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n846), .B(new_n850), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n716), .B(new_n761), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n699), .B(new_n501), .Z(new_n853));
  XNOR2_X1  g428(.A(new_n852), .B(new_n853), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n851), .A2(new_n854), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(G162), .B(G160), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(new_n627), .Z(new_n859));
  OR2_X1    g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT104), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n851), .A2(KEYINPUT104), .A3(new_n854), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n862), .A2(new_n863), .A3(new_n855), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n864), .A2(new_n859), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n865), .A2(KEYINPUT105), .ZN(new_n866));
  INV_X1    g441(.A(KEYINPUT105), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n867), .B1(new_n864), .B2(new_n859), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n845), .B(new_n860), .C1(new_n866), .C2(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g445(.A1(new_n829), .A2(G868), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n597), .A2(new_n604), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(new_n833), .ZN(new_n873));
  INV_X1    g448(.A(G299), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n597), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n874), .B1(new_n592), .B2(new_n596), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(KEYINPUT41), .A3(new_n877), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n592), .A2(new_n596), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(G299), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n881), .B1(new_n883), .B2(new_n876), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n880), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n879), .B1(new_n885), .B2(new_n873), .ZN(new_n886));
  INV_X1    g461(.A(KEYINPUT42), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n886), .A2(new_n887), .ZN(new_n890));
  OR2_X1    g465(.A1(G290), .A2(new_n787), .ZN(new_n891));
  NAND2_X1  g466(.A1(G290), .A2(new_n787), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(G166), .B(G305), .ZN(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n893), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n891), .A2(new_n892), .A3(new_n894), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  OAI22_X1  g473(.A1(new_n889), .A2(new_n890), .B1(KEYINPUT106), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n890), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n898), .A2(KEYINPUT106), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(new_n901), .A3(new_n888), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n871), .B1(new_n903), .B2(G868), .ZN(G295));
  AOI21_X1  g479(.A(new_n871), .B1(new_n903), .B2(G868), .ZN(G331));
  XNOR2_X1  g480(.A(G301), .B(G168), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n833), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n906), .A2(new_n828), .A3(new_n832), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n880), .A2(new_n884), .A3(new_n910), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n908), .A2(new_n875), .A3(new_n877), .A4(new_n909), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n898), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n911), .A2(new_n898), .A3(new_n912), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n845), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT43), .ZN(new_n918));
  NAND4_X1  g493(.A1(new_n914), .A2(new_n918), .A3(new_n845), .A4(new_n915), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT108), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n923), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n915), .A2(new_n845), .ZN(new_n925));
  OAI211_X1 g500(.A(new_n923), .B(KEYINPUT43), .C1(new_n925), .C2(new_n913), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  OAI21_X1  g502(.A(KEYINPUT44), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n919), .B(KEYINPUT107), .ZN(new_n929));
  OAI21_X1  g504(.A(new_n922), .B1(new_n928), .B2(new_n929), .ZN(G397));
  XNOR2_X1  g505(.A(new_n699), .B(new_n701), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n716), .B(G1996), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n776), .A2(new_n779), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n776), .A2(new_n779), .ZN(new_n934));
  AND4_X1   g509(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n501), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n467), .A2(new_n472), .A3(G40), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n941), .ZN(new_n942));
  NOR2_X1   g517(.A1(new_n935), .A2(new_n942), .ZN(new_n943));
  NOR3_X1   g518(.A1(G290), .A2(new_n942), .A3(G1986), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n943), .B1(KEYINPUT48), .B2(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n945), .B1(KEYINPUT48), .B2(new_n944), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n932), .A2(new_n931), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n934), .B1(new_n947), .B2(new_n941), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n699), .A2(G2067), .ZN(new_n949));
  OR3_X1    g524(.A1(new_n948), .A2(KEYINPUT126), .A3(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT126), .B1(new_n948), .B2(new_n949), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n950), .A2(new_n941), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n942), .B1(new_n931), .B2(new_n716), .ZN(new_n953));
  OR3_X1    g528(.A1(new_n942), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT46), .B1(new_n942), .B2(G1996), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT127), .B(KEYINPUT47), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n956), .B(new_n957), .ZN(new_n958));
  AND3_X1   g533(.A1(new_n946), .A2(new_n952), .A3(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT49), .ZN(new_n960));
  INV_X1    g535(.A(G1981), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n961), .B1(new_n577), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n963), .A2(G305), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n963), .A2(G305), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(G8), .ZN(new_n968));
  AND3_X1   g543(.A1(new_n501), .A2(KEYINPUT110), .A3(new_n936), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT110), .B1(new_n501), .B2(new_n936), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n940), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n968), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n577), .A2(new_n962), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n974), .A2(G1981), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(new_n792), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n976), .A2(KEYINPUT49), .A3(new_n964), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n967), .A2(new_n973), .A3(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G288), .A2(G1976), .ZN(new_n979));
  AND2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NOR2_X1   g555(.A1(G305), .A2(G1981), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT113), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n981), .B1(new_n978), .B2(new_n979), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT113), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n973), .A3(new_n985), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n783), .A2(new_n786), .A3(G1976), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n937), .A2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n501), .A2(KEYINPUT110), .A3(new_n936), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n989), .A2(new_n972), .A3(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n987), .A2(G8), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT52), .ZN(new_n993));
  INV_X1    g568(.A(G1976), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT52), .B1(G288), .B2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n973), .A2(new_n987), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n993), .A2(new_n978), .A3(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n493), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(new_n461), .B2(new_n462), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n1000), .A2(new_n495), .ZN(new_n1001));
  AOI22_X1  g576(.A1(new_n1001), .A2(new_n492), .B1(new_n499), .B2(new_n498), .ZN(new_n1002));
  AOI21_X1  g577(.A(G1384), .B1(new_n1002), .B2(new_n491), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n940), .B1(new_n1003), .B2(KEYINPUT45), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1384), .B1(new_n502), .B2(new_n504), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT109), .ZN(new_n1007));
  INV_X1    g582(.A(G1971), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n1004), .B(new_n1009), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1008), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n969), .B2(new_n970), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n503), .B1(new_n1002), .B2(new_n491), .ZN(new_n1014));
  AND4_X1   g589(.A1(new_n503), .A2(new_n491), .A3(new_n497), .A4(new_n500), .ZN(new_n1015));
  OAI211_X1 g590(.A(KEYINPUT50), .B(new_n936), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n940), .B1(new_n1013), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n968), .B1(new_n1011), .B2(new_n1019), .ZN(new_n1020));
  NOR2_X1   g595(.A1(G166), .A2(new_n968), .ZN(new_n1021));
  XOR2_X1   g596(.A(KEYINPUT111), .B(KEYINPUT55), .Z(new_n1022));
  XNOR2_X1  g597(.A(new_n1021), .B(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(new_n1023), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n998), .A2(new_n1020), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n986), .A2(new_n1025), .ZN(new_n1026));
  NOR2_X1   g601(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1027));
  NOR3_X1   g602(.A1(new_n969), .A2(new_n970), .A3(new_n1012), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1018), .B(new_n972), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g604(.A1(new_n1011), .A2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1023), .B1(new_n1030), .B2(new_n968), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n997), .B1(new_n1020), .B2(new_n1024), .ZN(new_n1032));
  INV_X1    g607(.A(G2084), .ZN(new_n1033));
  AOI21_X1  g608(.A(KEYINPUT50), .B1(new_n989), .B2(new_n990), .ZN(new_n1034));
  AOI211_X1 g609(.A(new_n1012), .B(G1384), .C1(new_n502), .C2(new_n504), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1033), .B(new_n972), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n936), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT45), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n989), .A2(new_n938), .A3(new_n990), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n940), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1036), .B1(new_n1040), .B2(G1966), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n1041), .A2(G8), .A3(G168), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1031), .A2(new_n1032), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  OR2_X1    g620(.A1(new_n1020), .A2(new_n1024), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1046), .A2(new_n1032), .A3(KEYINPUT63), .A4(new_n1042), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1026), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT62), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT120), .ZN(new_n1050));
  NAND3_X1  g625(.A1(G286), .A2(new_n1050), .A3(G8), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1050), .B1(G286), .B2(G8), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1041), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1053), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT51), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1055), .A2(new_n1056), .A3(new_n1051), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1057), .B1(new_n1041), .B2(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT121), .B1(new_n1055), .B2(new_n1051), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1052), .A2(new_n1053), .A3(new_n1060), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1059), .A2(new_n1061), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n1041), .B2(G8), .ZN(new_n1063));
  OAI22_X1  g638(.A1(KEYINPUT122), .A2(new_n1058), .B1(new_n1063), .B2(new_n1056), .ZN(new_n1064));
  AND2_X1   g639(.A1(new_n1058), .A2(KEYINPUT122), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1049), .B(new_n1054), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1067));
  INV_X1    g642(.A(G2078), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1040), .A2(KEYINPUT53), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n972), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT115), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1017), .A2(KEYINPUT115), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1070), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1037), .A2(new_n938), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1009), .B1(new_n1078), .B2(new_n1004), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1010), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1068), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(G171), .B1(new_n1077), .B2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1067), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1066), .A2(new_n1086), .ZN(new_n1087));
  OR2_X1    g662(.A1(new_n1058), .A2(KEYINPUT122), .ZN(new_n1088));
  AND2_X1   g663(.A1(new_n1041), .A2(G8), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT51), .B1(new_n1089), .B2(new_n1062), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1058), .A2(KEYINPUT122), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1088), .A2(new_n1090), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1049), .B1(new_n1092), .B2(new_n1054), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1048), .B1(new_n1087), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT54), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1017), .A2(KEYINPUT115), .ZN(new_n1096));
  AOI211_X1 g671(.A(new_n1072), .B(new_n940), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1069), .B1(new_n1098), .B2(new_n1074), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1099), .B2(new_n1083), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1004), .A2(KEYINPUT53), .A3(new_n1068), .A4(new_n939), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT123), .ZN(new_n1102));
  AND4_X1   g677(.A1(G301), .A2(new_n1083), .A3(new_n1076), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1095), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1054), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1067), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT57), .ZN(new_n1108));
  XNOR2_X1  g683(.A(G299), .B(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1109), .ZN(new_n1110));
  XNOR2_X1  g685(.A(KEYINPUT56), .B(G2072), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1004), .B(new_n1111), .C1(new_n1005), .C2(KEYINPUT45), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n972), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1114));
  INV_X1    g689(.A(G1956), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1110), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1073), .A2(new_n735), .A3(new_n1075), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n971), .A2(new_n701), .A3(new_n972), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1121), .B1(new_n882), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(new_n1109), .A3(new_n1112), .ZN(new_n1127));
  XNOR2_X1  g702(.A(new_n1127), .B(KEYINPUT114), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1125), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1116), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT118), .A3(new_n1110), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT118), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n1116), .B2(new_n1109), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1131), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1116), .A2(KEYINPUT119), .A3(new_n1109), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1131), .B1(new_n1127), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1121), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(G1996), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1078), .A2(new_n1142), .A3(new_n1004), .ZN(new_n1143));
  XOR2_X1   g718(.A(KEYINPUT58), .B(G1341), .Z(new_n1144));
  NAND2_X1  g719(.A1(new_n991), .A2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1143), .A2(new_n1145), .A3(KEYINPUT117), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT117), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n549), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n1148), .A2(KEYINPUT59), .ZN(new_n1149));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1150), .B(new_n549), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1151));
  NOR2_X1   g726(.A1(new_n882), .A2(KEYINPUT60), .ZN(new_n1152));
  AOI22_X1  g727(.A1(new_n1149), .A2(new_n1151), .B1(new_n1124), .B2(new_n1152), .ZN(new_n1153));
  AND3_X1   g728(.A1(new_n1122), .A2(new_n882), .A3(new_n1123), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n882), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT60), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g731(.A1(new_n1137), .A2(new_n1141), .A3(new_n1153), .A4(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1107), .B1(new_n1130), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1083), .A2(new_n1076), .A3(new_n1102), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1159), .A2(G171), .ZN(new_n1160));
  XOR2_X1   g735(.A(new_n1160), .B(KEYINPUT125), .Z(new_n1161));
  NOR3_X1   g736(.A1(new_n1077), .A2(new_n1084), .A3(G171), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT124), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1161), .A2(new_n1163), .A3(KEYINPUT54), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1094), .B1(new_n1158), .B2(new_n1164), .ZN(new_n1165));
  XNOR2_X1  g740(.A(G290), .B(new_n809), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n942), .B1(new_n935), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g742(.A(new_n959), .B1(new_n1165), .B2(new_n1167), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g743(.A1(G401), .A2(new_n459), .A3(G227), .A4(G229), .ZN(new_n1170));
  AND3_X1   g744(.A1(new_n1170), .A2(new_n869), .A3(new_n920), .ZN(G308));
  NAND3_X1  g745(.A1(new_n1170), .A2(new_n869), .A3(new_n920), .ZN(G225));
endmodule


