//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 0 0 1 0 1 0 0 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n695, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n925, new_n926, new_n927, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971;
  INV_X1    g000(.A(G137), .ZN(new_n187));
  AND3_X1   g001(.A1(new_n187), .A2(KEYINPUT11), .A3(G134), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT65), .A2(G134), .ZN(new_n189));
  NOR2_X1   g003(.A1(KEYINPUT65), .A2(G134), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(KEYINPUT11), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n188), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  NOR2_X1   g008(.A1(new_n189), .A2(new_n190), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n194), .B1(new_n195), .B2(G137), .ZN(new_n196));
  NOR4_X1   g010(.A1(new_n189), .A2(new_n190), .A3(KEYINPUT66), .A4(new_n187), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n193), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G131), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT67), .ZN(new_n200));
  INV_X1    g014(.A(G131), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n193), .B(new_n201), .C1(new_n196), .C2(new_n197), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  XNOR2_X1  g017(.A(G143), .B(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT0), .A3(G128), .ZN(new_n205));
  XNOR2_X1  g019(.A(KEYINPUT0), .B(G128), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n205), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n198), .A2(KEYINPUT67), .A3(G131), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  OR2_X1    g024(.A1(KEYINPUT65), .A2(G134), .ZN(new_n211));
  NAND2_X1  g025(.A1(KEYINPUT65), .A2(G134), .ZN(new_n212));
  AOI21_X1  g026(.A(G137), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n214));
  OAI22_X1  g028(.A1(new_n213), .A2(new_n214), .B1(G134), .B2(new_n187), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n214), .B(new_n187), .C1(new_n189), .C2(new_n190), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(G131), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G128), .ZN(new_n219));
  INV_X1    g033(.A(G146), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G143), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n219), .B1(new_n221), .B2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n222), .B(new_n204), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n218), .A2(new_n202), .A3(new_n223), .ZN(new_n224));
  AND2_X1   g038(.A1(new_n224), .A2(KEYINPUT30), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n210), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G119), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G116), .ZN(new_n228));
  INV_X1    g042(.A(G116), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G119), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G116), .B(G119), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(KEYINPUT70), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT2), .A2(G113), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(KEYINPUT69), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT69), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT2), .A3(G113), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(KEYINPUT2), .A2(G113), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n233), .B(new_n235), .C1(new_n240), .C2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT2), .ZN(new_n243));
  INV_X1    g057(.A(G113), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n237), .A2(new_n239), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n234), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n226), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT30), .B1(new_n210), .B2(new_n224), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(new_n247), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n210), .A2(new_n251), .A3(new_n224), .ZN(new_n252));
  INV_X1    g066(.A(G210), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n253), .A2(G237), .A3(G953), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n254), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(KEYINPUT26), .B(G101), .ZN(new_n256));
  XOR2_X1   g070(.A(new_n255), .B(new_n256), .Z(new_n257));
  NAND2_X1  g071(.A1(new_n252), .A2(new_n257), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT31), .B1(new_n250), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT28), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n252), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n210), .A2(new_n224), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n247), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n210), .A2(KEYINPUT28), .A3(new_n251), .A4(new_n224), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n261), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(new_n257), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT30), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n251), .B1(new_n210), .B2(new_n225), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(KEYINPUT71), .B(KEYINPUT31), .Z(new_n272));
  NAND4_X1  g086(.A1(new_n271), .A2(new_n252), .A3(new_n257), .A4(new_n272), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n259), .A2(new_n267), .A3(new_n273), .ZN(new_n274));
  NOR2_X1   g088(.A1(G472), .A2(G902), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT72), .B(KEYINPUT32), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n261), .A2(new_n263), .A3(new_n257), .A4(new_n264), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT29), .ZN(new_n281));
  AND3_X1   g095(.A1(new_n210), .A2(new_n251), .A3(new_n224), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n282), .B1(new_n269), .B2(new_n270), .ZN(new_n283));
  OAI211_X1 g097(.A(new_n280), .B(new_n281), .C1(new_n283), .C2(new_n257), .ZN(new_n284));
  INV_X1    g098(.A(G902), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n257), .A2(KEYINPUT29), .ZN(new_n287));
  INV_X1    g101(.A(new_n261), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT73), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n252), .A2(new_n289), .ZN(new_n290));
  NAND4_X1  g104(.A1(new_n210), .A2(KEYINPUT73), .A3(new_n251), .A4(new_n224), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n263), .A3(new_n291), .ZN(new_n292));
  AOI211_X1 g106(.A(new_n287), .B(new_n288), .C1(new_n292), .C2(KEYINPUT28), .ZN(new_n293));
  OAI21_X1  g107(.A(G472), .B1(new_n286), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n279), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT74), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n279), .A2(new_n294), .A3(KEYINPUT74), .A4(new_n295), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G217), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n301), .B1(G234), .B2(new_n285), .ZN(new_n302));
  INV_X1    g116(.A(G140), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G125), .ZN(new_n304));
  INV_X1    g118(.A(G125), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n305), .A2(G140), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n306), .A3(KEYINPUT75), .ZN(new_n307));
  OR3_X1    g121(.A1(new_n305), .A2(KEYINPUT75), .A3(G140), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT16), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n304), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G146), .ZN(new_n313));
  AND2_X1   g127(.A1(new_n304), .A2(new_n306), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n220), .ZN(new_n315));
  XOR2_X1   g129(.A(G119), .B(G128), .Z(new_n316));
  XNOR2_X1  g130(.A(KEYINPUT24), .B(G110), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT23), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n319), .B1(new_n227), .B2(G128), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n219), .A2(KEYINPUT23), .A3(G119), .ZN(new_n321));
  OAI211_X1 g135(.A(new_n320), .B(new_n321), .C1(G119), .C2(new_n219), .ZN(new_n322));
  OAI21_X1  g136(.A(new_n318), .B1(new_n322), .B2(G110), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT77), .ZN(new_n324));
  AND2_X1   g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n323), .A2(new_n324), .ZN(new_n326));
  OAI211_X1 g140(.A(new_n313), .B(new_n315), .C1(new_n325), .C2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT76), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n309), .A2(new_n220), .A3(new_n311), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n313), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n316), .A2(new_n317), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n331), .B1(G110), .B2(new_n322), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n328), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n309), .A2(new_n220), .A3(new_n311), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n220), .B1(new_n309), .B2(new_n311), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n332), .B(new_n328), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n327), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  XNOR2_X1  g152(.A(KEYINPUT22), .B(G137), .ZN(new_n339));
  INV_X1    g153(.A(G953), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n340), .A2(G221), .A3(G234), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n339), .B(new_n341), .Z(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n327), .B(new_n342), .C1(new_n333), .C2(new_n337), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n344), .A2(new_n285), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT79), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT78), .B(KEYINPUT25), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n346), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT25), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n350), .B2(new_n346), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n347), .B1(new_n346), .B2(new_n348), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n302), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n302), .A2(G902), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n344), .A2(new_n345), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n300), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G221), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT9), .B(G234), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n359), .B1(new_n361), .B2(new_n285), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT3), .ZN(new_n363));
  INV_X1    g177(.A(G107), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(G104), .ZN(new_n365));
  INV_X1    g179(.A(G104), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n365), .B1(new_n366), .B2(G107), .ZN(new_n367));
  OR2_X1    g181(.A1(KEYINPUT80), .A2(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(KEYINPUT80), .A2(G107), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n368), .A2(new_n363), .A3(G104), .A4(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(G101), .ZN(new_n372));
  INV_X1    g186(.A(G101), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n370), .A3(new_n373), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(KEYINPUT4), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n373), .B1(new_n367), .B2(new_n370), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n375), .A2(new_n208), .A3(new_n378), .ZN(new_n379));
  AOI21_X1  g193(.A(G104), .B1(new_n368), .B2(new_n369), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n366), .A2(G107), .ZN(new_n381));
  OAI21_X1  g195(.A(G101), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(new_n374), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(KEYINPUT10), .A3(new_n223), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  INV_X1    g200(.A(G143), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G146), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n221), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n222), .B(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n386), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n379), .A2(new_n385), .A3(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT83), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n203), .A2(new_n209), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n379), .A2(new_n385), .A3(KEYINPUT83), .A4(new_n391), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n394), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n395), .A2(KEYINPUT81), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT81), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n203), .A2(new_n400), .A3(new_n209), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n379), .A2(new_n385), .A3(new_n391), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n401), .A3(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G110), .B(G140), .ZN(new_n405));
  INV_X1    g219(.A(G227), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n406), .A2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n405), .B(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n404), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n408), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n403), .A2(KEYINPUT84), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n223), .A2(new_n374), .A3(new_n382), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n383), .A2(new_n390), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n396), .B(new_n414), .C1(new_n415), .C2(KEYINPUT12), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n203), .A2(new_n414), .A3(new_n209), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n203), .A2(new_n415), .A3(new_n209), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT12), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n416), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(KEYINPUT84), .B1(new_n403), .B2(new_n410), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n409), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(G469), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n424), .A2(new_n425), .A3(new_n285), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n417), .B1(new_n419), .B2(new_n418), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n403), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n392), .B1(KEYINPUT81), .B2(new_n395), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n408), .B1(new_n430), .B2(new_n401), .ZN(new_n431));
  AOI22_X1  g245(.A1(new_n429), .A2(new_n408), .B1(new_n431), .B2(new_n398), .ZN(new_n432));
  OAI21_X1  g246(.A(G469), .B1(new_n432), .B2(G902), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n362), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT85), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(G110), .B(G122), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n233), .A2(new_n235), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n440), .A2(KEYINPUT5), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n229), .A2(G119), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT5), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n244), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n441), .A2(new_n444), .B1(new_n245), .B2(new_n234), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n384), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n242), .A2(new_n246), .B1(new_n376), .B2(new_n377), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT86), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n447), .A2(new_n448), .A3(new_n375), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n448), .B1(new_n447), .B2(new_n375), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n439), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n375), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(KEYINPUT86), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n454), .A2(new_n438), .A3(new_n446), .A4(new_n449), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(KEYINPUT6), .A3(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT6), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(new_n439), .C1(new_n450), .C2(new_n451), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n205), .B(G125), .C1(new_n204), .C2(new_n206), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n390), .B2(G125), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n340), .A2(G224), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n460), .B(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n456), .A2(new_n458), .A3(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n444), .B1(new_n443), .B2(new_n231), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n374), .A2(new_n382), .A3(new_n464), .A4(new_n246), .ZN(new_n465));
  OAI211_X1 g279(.A(KEYINPUT87), .B(new_n465), .C1(new_n445), .C2(new_n384), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n465), .A2(KEYINPUT87), .ZN(new_n467));
  XOR2_X1   g281(.A(new_n438), .B(KEYINPUT8), .Z(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT88), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n461), .A2(KEYINPUT7), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n223), .A2(new_n305), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n470), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n461), .A2(KEYINPUT88), .A3(KEYINPUT7), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n473), .A2(new_n459), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n466), .A2(new_n469), .B1(new_n472), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(new_n455), .ZN(new_n478));
  AOI21_X1  g292(.A(KEYINPUT89), .B1(new_n478), .B2(new_n285), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n480));
  AOI211_X1 g294(.A(new_n480), .B(G902), .C1(new_n477), .C2(new_n455), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n463), .B1(new_n479), .B2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n463), .B(new_n483), .C1(new_n479), .C2(new_n481), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(G214), .B1(G237), .B2(G902), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI211_X1 g304(.A(KEYINPUT85), .B(new_n362), .C1(new_n426), .C2(new_n433), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NOR2_X1   g306(.A1(G475), .A2(G902), .ZN(new_n493));
  INV_X1    g307(.A(G237), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n340), .A3(G214), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(KEYINPUT90), .A3(new_n387), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT90), .B1(new_n495), .B2(new_n387), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n494), .A2(new_n340), .A3(G143), .A4(G214), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n501));
  XNOR2_X1  g315(.A(new_n500), .B(new_n501), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(KEYINPUT18), .A2(G131), .ZN(new_n504));
  AND2_X1   g318(.A1(new_n307), .A2(new_n308), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(G146), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n503), .A2(new_n504), .B1(new_n315), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n498), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n496), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n500), .B(KEYINPUT91), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n201), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n511), .A2(KEYINPUT18), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n507), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT94), .B(G104), .ZN(new_n515));
  XOR2_X1   g329(.A(new_n514), .B(new_n515), .Z(new_n516));
  NOR3_X1   g330(.A1(new_n499), .A2(new_n502), .A3(G131), .ZN(new_n517));
  NOR3_X1   g331(.A1(new_n517), .A2(new_n511), .A3(KEYINPUT17), .ZN(new_n518));
  OAI21_X1  g332(.A(G131), .B1(new_n499), .B2(new_n502), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n329), .B(new_n313), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n513), .B(new_n516), .C1(new_n518), .C2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT93), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n524), .A2(KEYINPUT19), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(KEYINPUT19), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n314), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(KEYINPUT92), .B1(new_n505), .B2(KEYINPUT19), .ZN(new_n528));
  AND4_X1   g342(.A1(KEYINPUT92), .A2(new_n307), .A3(KEYINPUT19), .A4(new_n308), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n220), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n530), .B(new_n313), .C1(new_n511), .C2(new_n517), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n516), .B1(new_n531), .B2(new_n513), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n493), .B1(new_n523), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT20), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT20), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n535), .B(new_n493), .C1(new_n523), .C2(new_n532), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n518), .A2(new_n521), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n516), .B1(new_n538), .B2(new_n513), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n285), .B1(new_n539), .B2(new_n523), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(G475), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(G952), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G953), .ZN(new_n544));
  NAND2_X1  g358(.A1(G234), .A2(G237), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XOR2_X1   g360(.A(KEYINPUT21), .B(G898), .Z(new_n547));
  NAND3_X1  g361(.A1(new_n545), .A2(G902), .A3(G953), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT99), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT97), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT95), .ZN(new_n553));
  INV_X1    g367(.A(G122), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n553), .B1(new_n554), .B2(G116), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n229), .A2(KEYINPUT95), .A3(G122), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT14), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n554), .A2(G116), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT14), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n555), .A2(new_n561), .A3(new_n556), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n558), .B(new_n559), .C1(new_n560), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n560), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  OAI21_X1  g379(.A(G107), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  NAND4_X1  g380(.A1(new_n557), .A2(new_n368), .A3(new_n369), .A4(new_n559), .ZN(new_n567));
  XNOR2_X1  g381(.A(G128), .B(G143), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n195), .B(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n557), .A2(new_n559), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n368), .A2(new_n369), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g387(.A1(new_n573), .A2(new_n567), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n195), .A2(new_n568), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n568), .A2(KEYINPUT13), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n387), .A2(G128), .ZN(new_n577));
  OAI21_X1  g391(.A(G134), .B1(new_n577), .B2(KEYINPUT13), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n575), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n574), .A2(new_n579), .ZN(new_n580));
  NOR3_X1   g394(.A1(new_n360), .A2(new_n301), .A3(G953), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n570), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n581), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n569), .A2(new_n567), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n562), .A2(new_n560), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n585), .A2(new_n559), .A3(new_n564), .A4(new_n558), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n586), .B2(G107), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n574), .A2(new_n579), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n583), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n582), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n552), .B1(new_n590), .B2(new_n285), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(G478), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n593), .A2(KEYINPUT15), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n552), .A3(new_n285), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n594), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n590), .A2(new_n285), .A3(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT98), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n590), .A2(KEYINPUT98), .A3(new_n285), .A4(new_n597), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NOR3_X1   g417(.A1(new_n542), .A2(new_n551), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n437), .A2(new_n490), .A3(new_n492), .A4(new_n604), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n358), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(new_n373), .ZN(G3));
  NOR2_X1   g421(.A1(new_n436), .A2(new_n491), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n274), .A2(new_n285), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(G472), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n610), .A2(new_n276), .ZN(new_n611));
  NOR2_X1   g425(.A1(new_n611), .A2(new_n356), .ZN(new_n612));
  AND2_X1   g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(new_n488), .ZN(new_n614));
  INV_X1    g428(.A(new_n486), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT100), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n485), .A2(KEYINPUT100), .A3(new_n486), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n621));
  AND2_X1   g435(.A1(new_n590), .A2(KEYINPUT33), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n590), .A2(KEYINPUT33), .ZN(new_n623));
  OAI211_X1 g437(.A(G478), .B(new_n285), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AND3_X1   g439(.A1(new_n542), .A2(new_n625), .A3(new_n550), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n613), .A2(new_n620), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n627), .B(KEYINPUT101), .ZN(new_n628));
  XNOR2_X1  g442(.A(KEYINPUT34), .B(G104), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  AND4_X1   g444(.A1(new_n550), .A2(new_n603), .A3(new_n541), .A4(new_n537), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n613), .A2(new_n620), .A3(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n343), .A2(KEYINPUT36), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n338), .B(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n354), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n353), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n604), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n639), .A2(new_n611), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n608), .A2(new_n490), .A3(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT37), .B(G110), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(KEYINPUT102), .B(KEYINPUT103), .ZN(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  AOI21_X1  g459(.A(new_n619), .B1(new_n298), .B2(new_n299), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n546), .B1(G900), .B2(new_n548), .ZN(new_n647));
  AND4_X1   g461(.A1(new_n541), .A2(new_n603), .A3(new_n537), .A4(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n638), .A2(new_n648), .ZN(new_n649));
  NOR3_X1   g463(.A1(new_n436), .A2(new_n491), .A3(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT104), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n646), .A2(KEYINPUT104), .A3(new_n650), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  XNOR2_X1  g469(.A(new_n647), .B(KEYINPUT39), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n608), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n657), .A2(KEYINPUT40), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(KEYINPUT40), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n274), .A2(KEYINPUT32), .A3(new_n275), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n283), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n257), .ZN(new_n664));
  OAI211_X1 g478(.A(new_n664), .B(new_n285), .C1(new_n292), .C2(new_n257), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n665), .A2(G472), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n662), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n487), .B(KEYINPUT38), .Z(new_n668));
  AND2_X1   g482(.A1(new_n353), .A2(new_n637), .ZN(new_n669));
  AOI22_X1  g483(.A1(new_n537), .A2(new_n541), .B1(new_n596), .B2(new_n602), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n488), .A3(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n658), .A2(new_n659), .A3(new_n667), .A4(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT105), .B(G143), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G45));
  NOR3_X1   g489(.A1(new_n436), .A2(new_n491), .A3(new_n669), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n542), .A2(new_n625), .A3(new_n647), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(KEYINPUT106), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n646), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G146), .ZN(G48));
  NAND2_X1  g495(.A1(new_n424), .A2(new_n285), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(G469), .ZN(new_n683));
  INV_X1    g497(.A(new_n362), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n683), .A2(new_n684), .A3(new_n426), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n685), .A2(new_n619), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(new_n626), .ZN(new_n687));
  OAI21_X1  g501(.A(KEYINPUT107), .B1(new_n358), .B2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n356), .B1(new_n298), .B2(new_n299), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n689), .A2(new_n686), .A3(new_n690), .A4(new_n626), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n688), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n692), .B(new_n693), .ZN(G15));
  NAND4_X1  g508(.A1(new_n300), .A2(new_n357), .A3(new_n631), .A4(new_n686), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G116), .ZN(G18));
  NOR2_X1   g510(.A1(new_n639), .A2(new_n685), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n646), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G119), .ZN(G21));
  NAND3_X1  g513(.A1(new_n617), .A2(new_n618), .A3(new_n670), .ZN(new_n700));
  NOR3_X1   g514(.A1(new_n700), .A2(new_n685), .A3(new_n551), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n356), .B(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n610), .A2(KEYINPUT108), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n609), .A2(new_n705), .A3(G472), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n288), .B1(new_n292), .B2(KEYINPUT28), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n259), .B(new_n273), .C1(new_n707), .C2(new_n257), .ZN(new_n708));
  AOI22_X1  g522(.A1(new_n704), .A2(new_n706), .B1(new_n275), .B2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n701), .A2(new_n703), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND2_X1  g525(.A1(new_n708), .A2(new_n275), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n705), .B1(new_n609), .B2(G472), .ZN(new_n713));
  INV_X1    g527(.A(G472), .ZN(new_n714));
  AOI211_X1 g528(.A(KEYINPUT108), .B(new_n714), .C1(new_n274), .C2(new_n285), .ZN(new_n715));
  OAI211_X1 g529(.A(new_n712), .B(new_n638), .C1(new_n713), .C2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(KEYINPUT110), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(KEYINPUT110), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n679), .B(new_n686), .C1(new_n718), .C2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G125), .ZN(G27));
  INV_X1    g535(.A(KEYINPUT32), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n276), .A2(new_n722), .ZN(new_n723));
  NAND3_X1  g537(.A1(new_n723), .A2(new_n294), .A3(new_n295), .ZN(new_n724));
  AND2_X1   g538(.A1(new_n703), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n426), .A2(new_n433), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(new_n684), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n485), .A2(new_n488), .A3(new_n486), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n725), .A2(KEYINPUT42), .A3(new_n679), .A4(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT42), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT74), .B1(new_n662), .B2(new_n294), .ZN(new_n732));
  AND4_X1   g546(.A1(KEYINPUT74), .A2(new_n279), .A3(new_n294), .A4(new_n295), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n357), .B(new_n729), .C1(new_n732), .C2(new_n733), .ZN(new_n734));
  OAI21_X1  g548(.A(new_n731), .B1(new_n734), .B2(new_n678), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G131), .ZN(G33));
  INV_X1    g551(.A(new_n648), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT111), .B1(new_n734), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT111), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n689), .A2(new_n740), .A3(new_n648), .A4(new_n729), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G134), .ZN(G36));
  INV_X1    g557(.A(KEYINPUT43), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n537), .A2(new_n541), .ZN(new_n745));
  AOI21_X1  g559(.A(new_n744), .B1(new_n745), .B2(new_n625), .ZN(new_n746));
  INV_X1    g560(.A(new_n625), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n747), .A2(new_n542), .A3(KEYINPUT43), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n749), .A2(new_n611), .A3(new_n638), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n751));
  OR2_X1    g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n728), .B1(new_n750), .B2(new_n751), .ZN(new_n753));
  OR2_X1    g567(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n432), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT46), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(new_n426), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n761));
  AOI21_X1  g575(.A(new_n362), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n752), .A2(new_n753), .A3(new_n656), .A4(new_n762), .ZN(new_n763));
  XOR2_X1   g577(.A(KEYINPUT112), .B(G137), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n763), .B(new_n764), .ZN(G39));
  INV_X1    g579(.A(new_n300), .ZN(new_n766));
  INV_X1    g580(.A(new_n728), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n766), .A2(new_n356), .A3(new_n679), .A4(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n768), .A2(KEYINPUT113), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n762), .B(KEYINPUT47), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n768), .A2(KEYINPUT113), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G140), .ZN(G42));
  NAND3_X1  g587(.A1(new_n668), .A2(new_n745), .A3(new_n625), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n683), .A2(new_n426), .ZN(new_n775));
  AOI211_X1 g589(.A(new_n667), .B(new_n774), .C1(KEYINPUT49), .C2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n703), .A2(new_n488), .A3(new_n684), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT114), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n775), .A2(KEYINPUT49), .ZN(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT115), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n776), .A2(new_n778), .A3(new_n780), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n646), .A2(KEYINPUT104), .A3(new_n650), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n720), .B1(new_n782), .B2(new_n651), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT117), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g599(.A(new_n720), .B(KEYINPUT117), .C1(new_n782), .C2(new_n651), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n353), .A2(new_n637), .A3(new_n647), .ZN(new_n787));
  OAI21_X1  g601(.A(KEYINPUT118), .B1(new_n727), .B2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT118), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n669), .A2(new_n434), .A3(new_n789), .A4(new_n647), .ZN(new_n790));
  INV_X1    g604(.A(new_n700), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n788), .A2(new_n790), .A3(new_n667), .A4(new_n791), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT119), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n700), .B1(new_n662), .B2(new_n666), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n795), .A2(KEYINPUT119), .A3(new_n790), .A4(new_n788), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n797), .A2(KEYINPUT52), .A3(new_n680), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n785), .A2(new_n786), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT52), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n680), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n783), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  OR2_X1    g617(.A1(new_n716), .A2(KEYINPUT110), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n678), .B1(new_n804), .B2(new_n717), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n542), .A2(new_n603), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n767), .A2(new_n806), .A3(new_n647), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n807), .B1(new_n298), .B2(new_n299), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n805), .A2(new_n729), .B1(new_n676), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n736), .A3(new_n742), .ZN(new_n810));
  OAI211_X1 g624(.A(new_n641), .B(new_n710), .C1(new_n358), .C2(new_n605), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n745), .A2(new_n550), .A3(new_n603), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n814), .B2(new_n489), .ZN(new_n815));
  NAND4_X1  g629(.A1(new_n631), .A2(KEYINPUT116), .A3(new_n488), .A4(new_n487), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n626), .A2(new_n488), .A3(new_n487), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n818), .A2(new_n608), .A3(new_n612), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n698), .A2(new_n695), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n812), .A2(new_n692), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n810), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(KEYINPUT53), .B1(new_n803), .B2(new_n822), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n646), .A2(new_n679), .ZN(new_n824));
  AOI22_X1  g638(.A1(new_n824), .A2(new_n676), .B1(new_n794), .B2(new_n796), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n825), .A2(new_n654), .A3(KEYINPUT52), .A4(new_n720), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n802), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n827), .A2(new_n822), .A3(KEYINPUT53), .ZN(new_n828));
  OAI21_X1  g642(.A(KEYINPUT54), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT54), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT53), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n831), .B1(new_n803), .B2(new_n822), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n827), .A2(new_n822), .A3(new_n831), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n746), .A2(new_n748), .A3(new_n546), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n703), .A2(new_n709), .A3(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n685), .ZN(new_n837));
  AND3_X1   g651(.A1(new_n668), .A2(new_n614), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT50), .Z(new_n840));
  NOR2_X1   g654(.A1(new_n775), .A2(new_n684), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n767), .B(new_n836), .C1(new_n770), .C2(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n667), .A2(new_n356), .A3(new_n546), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n685), .A2(new_n728), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR3_X1   g659(.A1(new_n845), .A2(new_n542), .A3(new_n625), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n835), .A2(new_n844), .ZN(new_n847));
  XOR2_X1   g661(.A(new_n847), .B(KEYINPUT120), .Z(new_n848));
  NAND2_X1  g662(.A1(new_n804), .A2(new_n717), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n846), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n840), .A2(new_n842), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n836), .A2(new_n686), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n542), .A2(new_n625), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n854), .B(new_n544), .C1(new_n855), .C2(new_n845), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n848), .A2(new_n725), .ZN(new_n857));
  OR2_X1    g671(.A1(new_n857), .A2(KEYINPUT48), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(KEYINPUT48), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n840), .A2(new_n842), .A3(KEYINPUT51), .A4(new_n850), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n853), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n829), .A2(new_n834), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n864));
  AND2_X1   g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n829), .A2(new_n834), .A3(new_n862), .A4(KEYINPUT121), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n543), .A2(new_n340), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n781), .B1(new_n865), .B2(new_n868), .ZN(G75));
  NAND2_X1  g683(.A1(new_n456), .A2(new_n458), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(new_n462), .ZN(new_n871));
  XOR2_X1   g685(.A(new_n871), .B(KEYINPUT55), .Z(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(KEYINPUT56), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n827), .A2(new_n822), .A3(new_n831), .ZN(new_n874));
  AOI22_X1  g688(.A1(new_n735), .A2(new_n730), .B1(new_n739), .B2(new_n741), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n698), .A2(new_n695), .A3(new_n819), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n811), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(new_n692), .A3(new_n877), .A4(new_n809), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n878), .B1(new_n799), .B2(new_n802), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n874), .B(G902), .C1(new_n879), .C2(new_n831), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n873), .B1(new_n880), .B2(new_n253), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n340), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OR3_X1    g698(.A1(new_n880), .A2(KEYINPUT122), .A3(new_n253), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT56), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT122), .B1(new_n880), .B2(new_n253), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n884), .B1(new_n888), .B2(new_n872), .ZN(G51));
  OAI211_X1 g703(.A(new_n874), .B(KEYINPUT54), .C1(new_n879), .C2(new_n831), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n834), .A2(new_n890), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n757), .B(KEYINPUT57), .Z(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n424), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n880), .A2(new_n756), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n882), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NOR2_X1   g710(.A1(new_n523), .A2(new_n532), .ZN(new_n897));
  NAND2_X1  g711(.A1(KEYINPUT58), .A2(G475), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n897), .B1(new_n880), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n899), .A2(new_n883), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n880), .A2(new_n897), .A3(new_n898), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n900), .A2(new_n901), .ZN(G60));
  OR2_X1    g716(.A1(new_n622), .A2(new_n623), .ZN(new_n903));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XNOR2_X1  g718(.A(new_n904), .B(KEYINPUT59), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n891), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n883), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n829), .A2(new_n834), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n903), .B1(new_n908), .B2(new_n905), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n909), .ZN(G63));
  INV_X1    g724(.A(KEYINPUT61), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n911), .A2(KEYINPUT123), .ZN(new_n913));
  NAND2_X1  g727(.A1(G217), .A2(G902), .ZN(new_n914));
  XOR2_X1   g728(.A(new_n914), .B(KEYINPUT60), .Z(new_n915));
  OAI211_X1 g729(.A(new_n874), .B(new_n915), .C1(new_n879), .C2(new_n831), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n344), .A2(new_n345), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n882), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n803), .A2(new_n822), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT53), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n920), .A2(new_n636), .A3(new_n874), .A4(new_n915), .ZN(new_n921));
  AOI211_X1 g735(.A(new_n912), .B(new_n913), .C1(new_n918), .C2(new_n921), .ZN(new_n922));
  AND4_X1   g736(.A1(KEYINPUT123), .A2(new_n918), .A3(new_n911), .A4(new_n921), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(G66));
  AOI21_X1  g738(.A(new_n340), .B1(new_n547), .B2(G224), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n821), .B2(new_n340), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n870), .B1(G898), .B2(new_n340), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n926), .B(new_n927), .Z(G69));
  NAND2_X1  g742(.A1(new_n269), .A2(new_n226), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n929), .B(new_n930), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT124), .Z(new_n932));
  NAND2_X1  g746(.A1(new_n745), .A2(new_n603), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT125), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n933), .A2(new_n934), .A3(new_n855), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n934), .B1(new_n933), .B2(new_n855), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n935), .A2(new_n936), .A3(new_n728), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n689), .A2(new_n937), .A3(new_n608), .A4(new_n656), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n763), .A2(KEYINPUT126), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT126), .B1(new_n763), .B2(new_n938), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n772), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n785), .A2(new_n673), .A3(new_n680), .A4(new_n786), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(KEYINPUT62), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n943), .B1(KEYINPUT62), .B2(new_n942), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n932), .B1(new_n944), .B2(new_n340), .ZN(new_n945));
  INV_X1    g759(.A(G900), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n931), .B1(new_n946), .B2(new_n340), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n725), .A2(new_n762), .A3(new_n656), .A4(new_n791), .ZN(new_n948));
  AND4_X1   g762(.A1(new_n763), .A2(new_n772), .A3(new_n875), .A4(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n785), .A2(new_n786), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n949), .A2(new_n680), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n947), .B1(new_n951), .B2(new_n340), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n340), .B1(G227), .B2(G900), .ZN(new_n953));
  OR3_X1    g767(.A1(new_n945), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n945), .B2(new_n952), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(G72));
  NAND2_X1  g770(.A1(G472), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT63), .Z(new_n958));
  NAND2_X1  g772(.A1(new_n283), .A2(new_n266), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n664), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n960), .B1(new_n823), .B2(new_n828), .ZN(new_n961));
  INV_X1    g775(.A(new_n958), .ZN(new_n962));
  INV_X1    g776(.A(new_n821), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n962), .B1(new_n951), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n883), .B(new_n961), .C1(new_n964), .C2(new_n959), .ZN(new_n965));
  OAI211_X1 g779(.A(KEYINPUT127), .B(new_n958), .C1(new_n944), .C2(new_n821), .ZN(new_n966));
  INV_X1    g780(.A(new_n664), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n958), .B1(new_n944), .B2(new_n821), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT127), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n965), .B1(new_n968), .B2(new_n971), .ZN(G57));
endmodule


