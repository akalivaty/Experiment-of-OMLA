//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 0 0 1 1 1 1 0 0 1 0 0 1 1 0 0 0 1 1 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n546, new_n547, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n559, new_n560, new_n561, new_n563,
    new_n564, new_n565, new_n566, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n588,
    new_n591, new_n593, new_n594, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1128, new_n1129, new_n1130,
    new_n1131;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT65), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT66), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  NAND2_X1  g032(.A1(G113), .A2(G2104), .ZN(new_n458));
  AND2_X1   g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NOR2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OAI21_X1  g037(.A(new_n458), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  AOI21_X1  g043(.A(G2105), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n466), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n469), .A2(G137), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n464), .A2(new_n471), .ZN(new_n472));
  XOR2_X1   g047(.A(new_n472), .B(KEYINPUT67), .Z(G160));
  NAND2_X1  g048(.A1(new_n469), .A2(G136), .ZN(new_n474));
  INV_X1    g049(.A(G2105), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n475), .B1(new_n467), .B2(new_n468), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n475), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n474), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  INV_X1    g056(.A(G138), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(new_n483), .B1(new_n459), .B2(new_n460), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT68), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n467), .A2(new_n468), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n486), .A2(new_n487), .A3(new_n483), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n485), .A2(new_n488), .A3(KEYINPUT4), .ZN(new_n489));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n484), .A2(KEYINPUT68), .A3(new_n490), .ZN(new_n491));
  OAI211_X1 g066(.A(G126), .B(G2105), .C1(new_n459), .C2(new_n460), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(G2105), .ZN(new_n495));
  NAND3_X1  g070(.A1(new_n493), .A2(new_n495), .A3(G2104), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n489), .A2(new_n491), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G50), .ZN(new_n501));
  NAND2_X1  g076(.A1(KEYINPUT69), .A2(G651), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT6), .ZN(new_n503));
  XNOR2_X1  g078(.A(new_n502), .B(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT5), .B(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n501), .A2(new_n505), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  AOI22_X1  g084(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n510));
  INV_X1    g085(.A(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  OR2_X1    g087(.A1(new_n509), .A2(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  INV_X1    g089(.A(new_n507), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G89), .ZN(new_n516));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n519), .B1(new_n505), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n516), .B(new_n518), .C1(new_n521), .C2(KEYINPUT70), .ZN(new_n522));
  AND2_X1   g097(.A1(new_n521), .A2(KEYINPUT70), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(G168));
  NAND2_X1  g099(.A1(G77), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(new_n506), .ZN(new_n526));
  INV_X1    g101(.A(G64), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n511), .B1(new_n528), .B2(KEYINPUT71), .ZN(new_n529));
  OAI21_X1  g104(.A(new_n529), .B1(KEYINPUT71), .B2(new_n528), .ZN(new_n530));
  INV_X1    g105(.A(new_n505), .ZN(new_n531));
  AOI22_X1  g106(.A1(G52), .A2(new_n531), .B1(new_n515), .B2(G90), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n530), .A2(new_n532), .ZN(G301));
  INV_X1    g108(.A(G301), .ZN(G171));
  AOI22_X1  g109(.A1(new_n506), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n535), .A2(new_n511), .ZN(new_n536));
  INV_X1    g111(.A(G81), .ZN(new_n537));
  XOR2_X1   g112(.A(KEYINPUT72), .B(G43), .Z(new_n538));
  OAI22_X1  g113(.A1(new_n537), .A2(new_n507), .B1(new_n505), .B2(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(KEYINPUT73), .ZN(new_n540));
  OR2_X1    g115(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n539), .A2(new_n540), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n536), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G860), .ZN(G153));
  NAND4_X1  g119(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT8), .ZN(new_n547));
  NAND4_X1  g122(.A1(G319), .A2(G483), .A3(G661), .A4(new_n547), .ZN(G188));
  INV_X1    g123(.A(G53), .ZN(new_n549));
  OR3_X1    g124(.A1(new_n505), .A2(KEYINPUT9), .A3(new_n549), .ZN(new_n550));
  OAI21_X1  g125(.A(KEYINPUT9), .B1(new_n505), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(G78), .A2(G543), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n526), .B2(new_n554), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n515), .A2(G91), .B1(new_n555), .B2(G651), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n552), .A2(new_n556), .ZN(G299));
  INV_X1    g132(.A(G168), .ZN(G286));
  NAND2_X1  g133(.A1(new_n531), .A2(G49), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n515), .A2(G87), .ZN(new_n560));
  OAI21_X1  g135(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(G288));
  NAND2_X1  g137(.A1(new_n515), .A2(G86), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n531), .A2(G48), .ZN(new_n564));
  AOI22_X1  g139(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n565), .A2(new_n511), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n563), .A2(new_n564), .A3(new_n566), .ZN(G305));
  NAND2_X1  g142(.A1(G72), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G60), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n526), .B2(new_n569), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n515), .A2(G85), .B1(new_n570), .B2(G651), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n531), .A2(G47), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n571), .A2(new_n572), .ZN(G290));
  INV_X1    g148(.A(G868), .ZN(new_n574));
  NOR2_X1   g149(.A1(G301), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n515), .A2(G92), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT10), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n576), .B(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n506), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n511), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(new_n581), .B1(new_n580), .B2(new_n579), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n531), .A2(G54), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n578), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g159(.A(new_n584), .B(KEYINPUT75), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n575), .B1(new_n585), .B2(new_n574), .ZN(G284));
  AOI21_X1  g161(.A(new_n575), .B1(new_n585), .B2(new_n574), .ZN(G321));
  NAND2_X1  g162(.A1(G299), .A2(new_n574), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(G168), .B2(new_n574), .ZN(G297));
  OAI21_X1  g164(.A(new_n588), .B1(G168), .B2(new_n574), .ZN(G280));
  INV_X1    g165(.A(G559), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n585), .B1(new_n591), .B2(G860), .ZN(G148));
  NAND2_X1  g167(.A1(new_n585), .A2(new_n591), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G868), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n594), .B1(G868), .B2(new_n543), .ZN(G323));
  XNOR2_X1  g170(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g171(.A1(new_n486), .A2(new_n470), .ZN(new_n597));
  XNOR2_X1  g172(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n598));
  XOR2_X1   g173(.A(new_n597), .B(new_n598), .Z(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT13), .ZN(new_n600));
  INV_X1    g175(.A(G2100), .ZN(new_n601));
  OR2_X1    g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n600), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n469), .A2(G135), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n476), .A2(G123), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n475), .A2(G111), .ZN(new_n606));
  OAI21_X1  g181(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  XOR2_X1   g183(.A(new_n608), .B(G2096), .Z(new_n609));
  NAND3_X1  g184(.A1(new_n602), .A2(new_n603), .A3(new_n609), .ZN(G156));
  XNOR2_X1  g185(.A(KEYINPUT15), .B(G2435), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT77), .B(G2438), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g188(.A(G2427), .B(G2430), .ZN(new_n614));
  OR2_X1    g189(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n613), .A2(new_n614), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n615), .A2(KEYINPUT14), .A3(new_n616), .ZN(new_n617));
  XOR2_X1   g192(.A(G2443), .B(G2446), .Z(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(G2451), .B(G2454), .Z(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT16), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT78), .Z(new_n622));
  XNOR2_X1  g197(.A(new_n619), .B(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(G1341), .B(G1348), .Z(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT79), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g201(.A(new_n626), .B(KEYINPUT80), .Z(new_n627));
  OAI211_X1 g202(.A(new_n627), .B(G14), .C1(new_n625), .C2(new_n623), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(G401));
  XOR2_X1   g204(.A(G2084), .B(G2090), .Z(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2072), .B(G2078), .Z(new_n632));
  XNOR2_X1  g207(.A(G2067), .B(G2678), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  NOR3_X1   g209(.A1(new_n631), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT81), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT18), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n632), .B(KEYINPUT17), .Z(new_n638));
  NOR3_X1   g213(.A1(new_n638), .A2(new_n633), .A3(new_n631), .ZN(new_n639));
  XOR2_X1   g214(.A(new_n639), .B(KEYINPUT82), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n633), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n630), .B1(new_n634), .B2(new_n632), .ZN(new_n642));
  AOI211_X1 g217(.A(new_n637), .B(new_n640), .C1(new_n641), .C2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2096), .B(G2100), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(G227));
  XOR2_X1   g220(.A(G1956), .B(G2474), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT84), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1961), .B(G1966), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G1971), .B(G1976), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT20), .Z(new_n655));
  OR3_X1    g230(.A1(new_n647), .A2(new_n653), .A3(new_n649), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT85), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n647), .A2(new_n649), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n658), .A2(new_n653), .A3(new_n650), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n655), .A2(new_n657), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1991), .B(G1996), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1981), .B(G1986), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(G229));
  INV_X1    g242(.A(G29), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G25), .ZN(new_n669));
  INV_X1    g244(.A(G95), .ZN(new_n670));
  AND3_X1   g245(.A1(new_n670), .A2(new_n475), .A3(KEYINPUT86), .ZN(new_n671));
  AOI21_X1  g246(.A(KEYINPUT86), .B1(new_n670), .B2(new_n475), .ZN(new_n672));
  OAI221_X1 g247(.A(G2104), .B1(G107), .B2(new_n475), .C1(new_n671), .C2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n469), .A2(G131), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n476), .A2(G119), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g251(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n669), .B1(new_n677), .B2(new_n668), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT35), .B(G1991), .Z(new_n679));
  XOR2_X1   g254(.A(new_n678), .B(new_n679), .Z(new_n680));
  MUX2_X1   g255(.A(G24), .B(G290), .S(G16), .Z(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT87), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(KEYINPUT90), .ZN(new_n684));
  AOI211_X1 g259(.A(new_n680), .B(new_n683), .C1(new_n684), .C2(KEYINPUT36), .ZN(new_n685));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G22), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n687), .B1(G166), .B2(new_n686), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1971), .ZN(new_n689));
  MUX2_X1   g264(.A(G23), .B(G288), .S(G16), .Z(new_n690));
  XNOR2_X1  g265(.A(KEYINPUT33), .B(G1976), .ZN(new_n691));
  XOR2_X1   g266(.A(new_n690), .B(new_n691), .Z(new_n692));
  INV_X1    g267(.A(KEYINPUT89), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n686), .A2(G6), .ZN(new_n694));
  INV_X1    g269(.A(G305), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n694), .B1(new_n695), .B2(new_n686), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT32), .B(G1981), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n697), .B(KEYINPUT88), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n696), .B(new_n698), .ZN(new_n699));
  AOI211_X1 g274(.A(new_n689), .B(new_n692), .C1(new_n693), .C2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(new_n693), .B2(new_n699), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n685), .B1(new_n701), .B2(KEYINPUT34), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(KEYINPUT34), .B2(new_n701), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n703), .A2(new_n684), .A3(KEYINPUT36), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n703), .B1(new_n684), .B2(KEYINPUT36), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n686), .A2(G4), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n585), .B2(new_n686), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT91), .B(G1348), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT92), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n707), .B(new_n709), .ZN(new_n710));
  NOR2_X1   g285(.A1(G171), .A2(new_n686), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G5), .B2(new_n686), .ZN(new_n712));
  INV_X1    g287(.A(G1961), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n686), .A2(G20), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT23), .ZN(new_n715));
  INV_X1    g290(.A(G299), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n715), .B1(new_n716), .B2(new_n686), .ZN(new_n717));
  OAI22_X1  g292(.A1(new_n712), .A2(new_n713), .B1(G1956), .B2(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n668), .A2(G32), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n476), .A2(G129), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n470), .A2(G105), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n722), .B1(G141), .B2(new_n469), .ZN(new_n723));
  NAND3_X1  g298(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(KEYINPUT95), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT26), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n723), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n719), .B1(new_n728), .B2(new_n668), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT27), .ZN(new_n730));
  INV_X1    g305(.A(G1996), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n730), .B(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(G160), .A2(G29), .ZN(new_n733));
  INV_X1    g308(.A(G34), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n734), .A2(KEYINPUT24), .ZN(new_n735));
  AOI21_X1  g310(.A(G29), .B1(new_n734), .B2(KEYINPUT24), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n735), .B1(new_n736), .B2(KEYINPUT94), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(KEYINPUT94), .B2(new_n736), .ZN(new_n738));
  AND2_X1   g313(.A1(new_n733), .A2(new_n738), .ZN(new_n739));
  AOI211_X1 g314(.A(new_n718), .B(new_n732), .C1(G2084), .C2(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n469), .A2(G140), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n476), .A2(G128), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n475), .A2(G116), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n745), .A2(G29), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n668), .A2(G26), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT28), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT93), .ZN(new_n750));
  INV_X1    g325(.A(G2067), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G19), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n543), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1341), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n686), .A2(G21), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n756), .B1(G168), .B2(new_n686), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT96), .B(G1966), .Z(new_n758));
  INV_X1    g333(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g334(.A(new_n752), .B(new_n755), .C1(new_n757), .C2(new_n759), .ZN(new_n760));
  OR2_X1    g335(.A1(new_n739), .A2(G2084), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n712), .A2(new_n713), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n717), .A2(G1956), .ZN(new_n763));
  NOR2_X1   g338(.A1(G29), .A2(G35), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(G162), .B2(G29), .ZN(new_n765));
  XNOR2_X1  g340(.A(KEYINPUT29), .B(G2090), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n765), .B(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n668), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n475), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  NAND2_X1  g345(.A1(new_n469), .A2(G139), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI22_X1  g347(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n773));
  NOR2_X1   g348(.A1(new_n773), .A2(new_n475), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n768), .B1(new_n775), .B2(new_n668), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G2072), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n767), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g353(.A1(new_n761), .A2(new_n762), .A3(new_n763), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g354(.A1(new_n757), .A2(new_n759), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n668), .A2(G27), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT97), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G164), .B2(new_n668), .ZN(new_n783));
  OR2_X1    g358(.A1(new_n783), .A2(G2078), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(G2078), .ZN(new_n785));
  XNOR2_X1  g360(.A(KEYINPUT30), .B(G28), .ZN(new_n786));
  OR2_X1    g361(.A1(KEYINPUT31), .A2(G11), .ZN(new_n787));
  NAND2_X1  g362(.A1(KEYINPUT31), .A2(G11), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n786), .A2(new_n668), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(new_n608), .B2(new_n668), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n776), .B2(G2072), .ZN(new_n791));
  NAND3_X1  g366(.A1(new_n784), .A2(new_n785), .A3(new_n791), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n779), .A2(new_n780), .A3(new_n792), .ZN(new_n793));
  AND4_X1   g368(.A1(new_n710), .A2(new_n740), .A3(new_n760), .A4(new_n793), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n704), .A2(new_n705), .A3(new_n794), .ZN(G150));
  INV_X1    g370(.A(G150), .ZN(G311));
  AOI22_X1  g371(.A1(G55), .A2(new_n531), .B1(new_n515), .B2(G93), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n506), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n798), .A2(new_n511), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g376(.A1(new_n799), .A2(KEYINPUT99), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G860), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n805), .B(KEYINPUT37), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n585), .A2(G559), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(new_n803), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT100), .ZN(new_n811));
  NOR2_X1   g386(.A1(new_n543), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g387(.A1(new_n539), .A2(new_n540), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n539), .A2(new_n540), .ZN(new_n814));
  OAI22_X1  g389(.A1(new_n813), .A2(new_n814), .B1(new_n511), .B2(new_n535), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n810), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n543), .A2(new_n811), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n815), .A2(KEYINPUT100), .ZN(new_n819));
  NAND3_X1  g394(.A1(new_n818), .A2(new_n819), .A3(new_n803), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n817), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n809), .B(new_n821), .ZN(new_n822));
  AND2_X1   g397(.A1(new_n822), .A2(KEYINPUT39), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n804), .B1(new_n822), .B2(KEYINPUT39), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n806), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(G145));
  OAI21_X1  g402(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n828));
  INV_X1    g403(.A(G118), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n828), .B1(new_n829), .B2(G2105), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n476), .A2(G130), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT104), .ZN(new_n832));
  AOI211_X1 g407(.A(new_n830), .B(new_n832), .C1(G142), .C2(new_n469), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n599), .B(new_n676), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n833), .B(new_n834), .Z(new_n835));
  XNOR2_X1  g410(.A(new_n727), .B(G164), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n745), .B(KEYINPUT102), .Z(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OR3_X1    g413(.A1(new_n838), .A2(KEYINPUT103), .A3(new_n775), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n775), .B(KEYINPUT103), .Z(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n835), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT105), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n839), .A2(new_n835), .A3(new_n841), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n842), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n845), .B1(new_n843), .B2(new_n844), .ZN(new_n846));
  XNOR2_X1  g421(.A(G160), .B(new_n608), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(G162), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n846), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT106), .B(G37), .Z(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n842), .A2(new_n848), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n851), .B1(new_n852), .B2(new_n844), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n849), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g430(.A(new_n593), .B(new_n821), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n584), .B(new_n716), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n857), .B(KEYINPUT41), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(new_n857), .B2(new_n856), .ZN(new_n860));
  OR2_X1    g435(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n861));
  XOR2_X1   g436(.A(G303), .B(G288), .Z(new_n862));
  XNOR2_X1  g437(.A(new_n695), .B(G290), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n862), .B(new_n863), .Z(new_n864));
  NAND2_X1  g439(.A1(new_n860), .A2(KEYINPUT42), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n861), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n864), .B1(new_n861), .B2(new_n865), .ZN(new_n867));
  OAI21_X1  g442(.A(G868), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n810), .A2(new_n574), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(G295));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n869), .ZN(G331));
  INV_X1    g446(.A(KEYINPUT44), .ZN(new_n872));
  INV_X1    g447(.A(new_n820), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n803), .B1(new_n818), .B2(new_n819), .ZN(new_n874));
  NOR3_X1   g449(.A1(new_n873), .A2(G171), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(G301), .B1(new_n817), .B2(new_n820), .ZN(new_n876));
  OAI21_X1  g451(.A(G286), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(G171), .B1(new_n873), .B2(new_n874), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n817), .A2(G301), .A3(new_n820), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n878), .A2(G168), .A3(new_n879), .ZN(new_n880));
  AND3_X1   g455(.A1(new_n877), .A2(new_n857), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g456(.A(new_n858), .B1(new_n877), .B2(new_n880), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n864), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(G37), .ZN(new_n884));
  XNOR2_X1  g459(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n885));
  INV_X1    g460(.A(new_n858), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n875), .A2(new_n876), .A3(G286), .ZN(new_n887));
  AOI21_X1  g462(.A(G168), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n886), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n864), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n877), .A2(new_n857), .A3(new_n880), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n883), .A2(new_n884), .A3(new_n885), .A4(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n872), .B1(new_n893), .B2(KEYINPUT108), .ZN(new_n894));
  NOR3_X1   g469(.A1(new_n881), .A2(new_n882), .A3(new_n864), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n890), .B1(new_n889), .B2(new_n891), .ZN(new_n896));
  NOR2_X1   g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT108), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n884), .A4(new_n885), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n883), .A2(new_n850), .A3(new_n892), .ZN(new_n900));
  AND2_X1   g475(.A1(new_n900), .A2(KEYINPUT109), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT109), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n883), .A2(new_n902), .A3(new_n850), .A4(new_n892), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT43), .ZN(new_n904));
  OAI211_X1 g479(.A(new_n894), .B(new_n899), .C1(new_n901), .C2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n885), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n897), .A2(new_n884), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n900), .A2(new_n885), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n872), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n905), .A2(new_n909), .ZN(G397));
  INV_X1    g485(.A(G1384), .ZN(new_n911));
  AND3_X1   g486(.A1(new_n485), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n491), .A2(new_n496), .A3(new_n492), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT45), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n464), .A2(G40), .A3(new_n471), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n918), .A2(G1986), .A3(G290), .ZN(new_n919));
  NOR2_X1   g494(.A1(G290), .A2(G1986), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n918), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XOR2_X1   g497(.A(new_n922), .B(KEYINPUT110), .Z(new_n923));
  XNOR2_X1  g498(.A(new_n727), .B(new_n731), .ZN(new_n924));
  XNOR2_X1  g499(.A(new_n745), .B(new_n751), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g501(.A(new_n676), .B(new_n679), .Z(new_n927));
  OAI21_X1  g502(.A(new_n918), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n923), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n917), .B1(new_n914), .B2(KEYINPUT50), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT50), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n499), .A2(new_n931), .A3(new_n911), .ZN(new_n932));
  XOR2_X1   g507(.A(KEYINPUT116), .B(G2084), .Z(new_n933));
  NAND3_X1  g508(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT115), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n915), .A2(G1384), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n917), .B1(new_n499), .B2(new_n936), .ZN(new_n937));
  AOI211_X1 g512(.A(new_n935), .B(new_n759), .C1(new_n916), .C2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n917), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n936), .B1(new_n912), .B2(new_n913), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n487), .B1(new_n486), .B2(new_n483), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n497), .B1(new_n490), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G1384), .B1(new_n942), .B2(new_n489), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n939), .B(new_n940), .C1(new_n943), .C2(KEYINPUT45), .ZN(new_n944));
  AOI21_X1  g519(.A(KEYINPUT115), .B1(new_n944), .B2(new_n758), .ZN(new_n945));
  OAI211_X1 g520(.A(G168), .B(new_n934), .C1(new_n938), .C2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G8), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT51), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(KEYINPUT118), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n948), .A2(KEYINPUT118), .ZN(new_n950));
  INV_X1    g525(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n934), .B1(new_n938), .B2(new_n945), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n953), .A2(G8), .A3(G286), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n951), .B1(new_n946), .B2(new_n949), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT119), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT62), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n946), .A2(new_n949), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n950), .ZN(new_n960));
  INV_X1    g535(.A(KEYINPUT119), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n960), .A2(new_n961), .A3(new_n954), .A4(new_n952), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n957), .A2(new_n958), .A3(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n914), .A2(KEYINPUT50), .ZN(new_n964));
  INV_X1    g539(.A(G2090), .ZN(new_n965));
  NAND4_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n932), .A4(new_n939), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT112), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n930), .A2(new_n968), .A3(new_n965), .A4(new_n932), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n940), .A2(new_n939), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT111), .B1(new_n943), .B2(KEYINPUT45), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT111), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n914), .A2(new_n972), .A3(new_n915), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  OAI211_X1 g549(.A(new_n967), .B(new_n969), .C1(G1971), .C2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(G303), .A2(G8), .ZN(new_n976));
  XNOR2_X1  g551(.A(new_n976), .B(KEYINPUT55), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n975), .A2(new_n978), .A3(G8), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n943), .A2(KEYINPUT111), .A3(KEYINPUT45), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n972), .B1(new_n914), .B2(new_n915), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n937), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(G1971), .ZN(new_n983));
  AND3_X1   g558(.A1(new_n964), .A2(new_n932), .A3(new_n939), .ZN(new_n984));
  AOI22_X1  g559(.A1(new_n982), .A2(new_n983), .B1(new_n984), .B2(new_n965), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n977), .B1(new_n985), .B2(new_n947), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n943), .A2(new_n939), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(G8), .ZN(new_n988));
  NAND4_X1  g563(.A1(new_n560), .A2(new_n559), .A3(G1976), .A4(new_n561), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g565(.A(KEYINPUT52), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1976), .ZN(new_n992));
  AOI21_X1  g567(.A(KEYINPUT52), .B1(G288), .B2(new_n992), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n993), .A2(G8), .A3(new_n987), .A4(new_n989), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n991), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT113), .B(G1981), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n563), .A2(new_n564), .A3(new_n566), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT114), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n996), .A2(KEYINPUT114), .A3(KEYINPUT49), .A4(new_n998), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT49), .B1(new_n996), .B2(new_n998), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(new_n988), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n995), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n979), .A2(new_n986), .A3(new_n1006), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n964), .A2(new_n932), .A3(new_n939), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(new_n713), .ZN(new_n1009));
  INV_X1    g584(.A(new_n944), .ZN(new_n1010));
  INV_X1    g585(.A(G2078), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n1011), .ZN(new_n1012));
  AOI211_X1 g587(.A(G2078), .B(new_n970), .C1(new_n971), .C2(new_n973), .ZN(new_n1013));
  OAI211_X1 g588(.A(new_n1009), .B(new_n1012), .C1(new_n1013), .C2(KEYINPUT53), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1014), .A2(G171), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1007), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n963), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT122), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n963), .A2(KEYINPUT122), .A3(new_n1016), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n957), .A2(new_n962), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(KEYINPUT62), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1019), .A2(new_n1020), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT57), .ZN(new_n1024));
  XNOR2_X1  g599(.A(G299), .B(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT56), .B(G2072), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n974), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1956), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1008), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(G1348), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1008), .A2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n987), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1033), .A2(new_n751), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n584), .B1(new_n1032), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1027), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1030), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT61), .ZN(new_n1038));
  AND3_X1   g613(.A1(new_n1027), .A2(new_n1025), .A3(new_n1029), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1038), .B1(new_n1039), .B2(new_n1030), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1025), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1026), .ZN(new_n1042));
  NOR2_X1   g617(.A1(new_n982), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(new_n1029), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1041), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT61), .A3(new_n1036), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1040), .A2(new_n1046), .ZN(new_n1047));
  AND3_X1   g622(.A1(new_n1032), .A2(new_n584), .A3(new_n1034), .ZN(new_n1048));
  OAI21_X1  g623(.A(KEYINPUT60), .B1(new_n1048), .B2(new_n1035), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT59), .ZN(new_n1050));
  XNOR2_X1  g625(.A(KEYINPUT58), .B(G1341), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1033), .A2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n974), .B2(new_n731), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1050), .B1(new_n1053), .B2(new_n815), .ZN(new_n1054));
  NOR2_X1   g629(.A1(new_n584), .A2(KEYINPUT60), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1055), .A2(new_n1034), .A3(new_n1032), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n982), .A2(G1996), .ZN(new_n1057));
  OAI211_X1 g632(.A(KEYINPUT59), .B(new_n543), .C1(new_n1057), .C2(new_n1052), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n1049), .A2(new_n1054), .A3(new_n1056), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1037), .B1(new_n1047), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n1061));
  XNOR2_X1  g636(.A(KEYINPUT120), .B(G2078), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1010), .A2(KEYINPUT53), .A3(new_n1062), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n1009), .B(new_n1063), .C1(new_n1013), .C2(KEYINPUT53), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1064), .B2(G171), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1014), .A2(G171), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1066), .A2(KEYINPUT121), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT121), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1014), .A2(new_n1068), .A3(G171), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1065), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1015), .B1(new_n1064), .B2(G171), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1007), .B1(new_n1071), .B2(new_n1061), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1021), .A2(new_n1060), .A3(new_n1070), .A4(new_n1072), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n979), .A2(new_n1006), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n930), .A2(new_n932), .A3(new_n933), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT45), .B1(new_n499), .B2(new_n911), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n758), .B1(new_n970), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n935), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n944), .A2(KEYINPUT115), .A3(new_n758), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NOR3_X1   g655(.A1(new_n1080), .A2(new_n947), .A3(G286), .ZN(new_n1081));
  INV_X1    g656(.A(new_n975), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n977), .B1(new_n1082), .B2(new_n947), .ZN(new_n1083));
  NAND4_X1  g658(.A1(new_n1074), .A2(KEYINPUT63), .A3(new_n1081), .A4(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1081), .A2(new_n979), .A3(new_n986), .A4(new_n1006), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n1085), .A2(KEYINPUT117), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1087), .B1(new_n1085), .B2(KEYINPUT117), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1084), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g664(.A(G1976), .B(G288), .C1(new_n1003), .C2(new_n1005), .ZN(new_n1090));
  INV_X1    g665(.A(new_n998), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(new_n988), .ZN(new_n1093));
  INV_X1    g668(.A(new_n979), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1006), .ZN(new_n1095));
  AND3_X1   g670(.A1(new_n1073), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n929), .B1(new_n1023), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n728), .A2(new_n925), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n918), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT125), .Z(new_n1100));
  NAND2_X1  g675(.A1(new_n918), .A2(new_n731), .ZN(new_n1101));
  XNOR2_X1  g676(.A(new_n1101), .B(KEYINPUT46), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g678(.A(new_n1103), .B(KEYINPUT47), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n921), .B(KEYINPUT126), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT48), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1105), .A2(new_n1106), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n928), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n677), .A2(new_n679), .ZN(new_n1110));
  XOR2_X1   g685(.A(new_n1110), .B(KEYINPUT123), .Z(new_n1111));
  INV_X1    g686(.A(new_n1111), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n926), .B2(new_n918), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n745), .A2(G2067), .ZN(new_n1114));
  OR3_X1    g689(.A1(new_n1113), .A2(KEYINPUT124), .A3(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(KEYINPUT124), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1115), .A2(new_n918), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1104), .A2(new_n1109), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(KEYINPUT127), .B1(new_n1097), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT127), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1118), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1073), .A2(new_n1089), .A3(new_n1095), .ZN(new_n1122));
  AOI22_X1  g697(.A1(new_n1017), .A2(new_n1018), .B1(KEYINPUT62), .B2(new_n1021), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(new_n1020), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1120), .B(new_n1121), .C1(new_n1124), .C2(new_n929), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1119), .A2(new_n1125), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g701(.A(G319), .ZN(new_n1128));
  NOR2_X1   g702(.A1(G227), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g703(.A1(new_n666), .A2(new_n628), .A3(new_n1129), .ZN(new_n1130));
  AOI21_X1  g704(.A(new_n1130), .B1(new_n853), .B2(new_n849), .ZN(new_n1131));
  AND3_X1   g705(.A1(new_n1131), .A2(new_n908), .A3(new_n907), .ZN(G308));
  NAND3_X1  g706(.A1(new_n1131), .A2(new_n908), .A3(new_n907), .ZN(G225));
endmodule


