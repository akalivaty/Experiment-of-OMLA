//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:14 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n597, new_n598, new_n601, new_n603, new_n604, new_n605,
    new_n606, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1233,
    new_n1234, new_n1235;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  XOR2_X1   g004(.A(KEYINPUT64), .B(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT65), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  XNOR2_X1  g033(.A(KEYINPUT3), .B(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G125), .ZN(new_n460));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  AOI21_X1  g036(.A(new_n458), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND3_X1  g037(.A1(new_n459), .A2(G137), .A3(new_n458), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n458), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(G101), .ZN(new_n465));
  OR3_X1    g040(.A1(new_n464), .A2(KEYINPUT66), .A3(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(KEYINPUT66), .B1(new_n464), .B2(new_n465), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT67), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g045(.A1(new_n463), .A2(new_n466), .A3(KEYINPUT67), .A4(new_n467), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n459), .A2(new_n458), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G136), .ZN(new_n475));
  AND2_X1   g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NOR2_X1   g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n478), .A2(new_n458), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n475), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND3_X1  g059(.A1(new_n459), .A2(G138), .A3(new_n458), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT68), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n459), .A2(KEYINPUT68), .A3(G138), .A4(new_n458), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n487), .A2(KEYINPUT4), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n478), .B2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G2104), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n492), .A2(G2105), .B1(G102), .B2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n485), .A2(new_n486), .A3(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n489), .A2(new_n495), .A3(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(new_n498), .ZN(G164));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n502));
  OAI21_X1  g077(.A(KEYINPUT69), .B1(new_n502), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT69), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(new_n500), .A3(KEYINPUT5), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n501), .B1(new_n503), .B2(new_n505), .ZN(new_n506));
  AOI22_X1  g081(.A1(new_n506), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G651), .ZN(new_n508));
  NOR2_X1   g083(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g084(.A(KEYINPUT6), .B(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n510), .A2(G543), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n511), .A2(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n509), .A2(new_n515), .ZN(G166));
  AND3_X1   g091(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT70), .ZN(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT7), .ZN(new_n520));
  INV_X1    g095(.A(new_n511), .ZN(new_n521));
  INV_X1    g096(.A(new_n514), .ZN(new_n522));
  AOI22_X1  g097(.A1(new_n521), .A2(G89), .B1(new_n522), .B2(G51), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n518), .A2(new_n520), .A3(new_n523), .ZN(G286));
  INV_X1    g099(.A(G286), .ZN(G168));
  AOI22_X1  g100(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n508), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  OAI22_X1  g104(.A1(new_n511), .A2(new_n528), .B1(new_n529), .B2(new_n514), .ZN(new_n530));
  OR2_X1    g105(.A1(new_n527), .A2(new_n530), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  AND3_X1   g107(.A1(new_n506), .A2(G81), .A3(new_n510), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n522), .A2(G43), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT71), .ZN(new_n536));
  NAND2_X1  g111(.A1(G68), .A2(G543), .ZN(new_n537));
  INV_X1    g112(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n506), .B2(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n536), .B1(new_n539), .B2(new_n508), .ZN(new_n540));
  INV_X1    g115(.A(new_n501), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n504), .B1(KEYINPUT5), .B2(new_n500), .ZN(new_n542));
  NOR3_X1   g117(.A1(new_n502), .A2(KEYINPUT69), .A3(G543), .ZN(new_n543));
  OAI211_X1 g118(.A(G56), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(new_n537), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n545), .A2(KEYINPUT71), .A3(G651), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n533), .B(new_n535), .C1(new_n540), .C2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G860), .ZN(G153));
  AND3_X1   g123(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G36), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT73), .ZN(new_n552));
  XOR2_X1   g127(.A(KEYINPUT72), .B(KEYINPUT8), .Z(new_n553));
  XNOR2_X1  g128(.A(new_n552), .B(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n549), .A2(new_n554), .ZN(G188));
  NAND3_X1  g130(.A1(new_n506), .A2(G91), .A3(new_n510), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT75), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n556), .B(new_n557), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT74), .B(KEYINPUT9), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n522), .A2(G53), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  INV_X1    g136(.A(G53), .ZN(new_n562));
  OAI211_X1 g137(.A(KEYINPUT74), .B(new_n561), .C1(new_n514), .C2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n506), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI211_X1 g139(.A(new_n560), .B(new_n563), .C1(new_n564), .C2(new_n508), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n558), .A2(new_n565), .ZN(G299));
  INV_X1    g141(.A(G166), .ZN(G303));
  OAI21_X1  g142(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n506), .A2(G87), .A3(new_n510), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n510), .A2(G49), .A3(G543), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(G288));
  NAND2_X1  g146(.A1(new_n522), .A2(G48), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n506), .A2(G86), .A3(new_n510), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n506), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n574));
  OAI211_X1 g149(.A(new_n572), .B(new_n573), .C1(new_n574), .C2(new_n508), .ZN(G305));
  AOI22_X1  g150(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n576), .A2(new_n508), .ZN(new_n577));
  INV_X1    g152(.A(G85), .ZN(new_n578));
  INV_X1    g153(.A(G47), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n511), .A2(new_n578), .B1(new_n579), .B2(new_n514), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n577), .A2(new_n580), .ZN(G290));
  NAND2_X1  g156(.A1(G301), .A2(G868), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n506), .A2(G66), .ZN(new_n583));
  INV_X1    g158(.A(G79), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n584), .B2(new_n500), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n522), .A2(G54), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT76), .B(KEYINPUT10), .Z(new_n588));
  NAND4_X1  g163(.A1(new_n506), .A2(G92), .A3(new_n510), .A4(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n588), .ZN(new_n590));
  INV_X1    g165(.A(G92), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n511), .B2(new_n591), .ZN(new_n592));
  NAND4_X1  g167(.A1(new_n586), .A2(new_n587), .A3(new_n589), .A4(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n582), .B1(new_n594), .B2(G868), .ZN(G284));
  OAI21_X1  g170(.A(new_n582), .B1(new_n594), .B2(G868), .ZN(G321));
  INV_X1    g171(.A(G868), .ZN(new_n597));
  NAND2_X1  g172(.A1(G299), .A2(new_n597), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G297));
  OAI21_X1  g174(.A(new_n598), .B1(G168), .B2(new_n597), .ZN(G280));
  INV_X1    g175(.A(G559), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n594), .B1(new_n601), .B2(G860), .ZN(G148));
  NAND2_X1  g177(.A1(new_n594), .A2(new_n601), .ZN(new_n603));
  INV_X1    g178(.A(new_n603), .ZN(new_n604));
  OR3_X1    g179(.A1(new_n604), .A2(KEYINPUT77), .A3(new_n597), .ZN(new_n605));
  OAI21_X1  g180(.A(KEYINPUT77), .B1(new_n604), .B2(new_n597), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n605), .B(new_n606), .C1(G868), .C2(new_n547), .ZN(G323));
  XNOR2_X1  g182(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g183(.A1(new_n459), .A2(new_n494), .ZN(new_n609));
  XOR2_X1   g184(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2100), .ZN(new_n611));
  XOR2_X1   g186(.A(KEYINPUT78), .B(KEYINPUT13), .Z(new_n612));
  XNOR2_X1  g187(.A(new_n611), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n474), .A2(G135), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n479), .A2(G123), .ZN(new_n615));
  NOR2_X1   g190(.A1(G99), .A2(G2105), .ZN(new_n616));
  OAI21_X1  g191(.A(G2104), .B1(new_n458), .B2(G111), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n614), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  XOR2_X1   g193(.A(new_n618), .B(G2096), .Z(new_n619));
  NAND2_X1  g194(.A1(new_n613), .A2(new_n619), .ZN(G156));
  XOR2_X1   g195(.A(G1341), .B(G1348), .Z(new_n621));
  INV_X1    g196(.A(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(G2451), .B(G2454), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT16), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2446), .ZN(new_n625));
  INV_X1    g200(.A(new_n625), .ZN(new_n626));
  INV_X1    g201(.A(G2443), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT15), .B(G2435), .ZN(new_n628));
  INV_X1    g203(.A(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(G2427), .B(G2430), .Z(new_n631));
  OAI21_X1  g206(.A(KEYINPUT14), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT79), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n630), .A2(new_n631), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n627), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n633), .A2(new_n627), .A3(new_n634), .ZN(new_n637));
  AOI21_X1  g212(.A(new_n626), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g213(.A(new_n637), .ZN(new_n639));
  NOR3_X1   g214(.A1(new_n639), .A2(new_n635), .A3(new_n625), .ZN(new_n640));
  OAI21_X1  g215(.A(new_n622), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n625), .B1(new_n639), .B2(new_n635), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n636), .A2(new_n637), .A3(new_n626), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n643), .A3(new_n621), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(G14), .A3(new_n644), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  INV_X1    g222(.A(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2067), .B(G2678), .Z(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n650), .A2(new_n651), .A3(KEYINPUT17), .ZN(new_n652));
  INV_X1    g227(.A(KEYINPUT18), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2072), .B(G2078), .Z(new_n655));
  AOI21_X1  g230(.A(new_n655), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2096), .B(G2100), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT80), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(G227));
  XNOR2_X1  g236(.A(G1971), .B(G1976), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT19), .ZN(new_n663));
  XOR2_X1   g238(.A(G1956), .B(G2474), .Z(new_n664));
  XOR2_X1   g239(.A(G1961), .B(G1966), .Z(new_n665));
  OR2_X1    g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n664), .A2(new_n665), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT81), .B(KEYINPUT20), .Z(new_n670));
  AOI21_X1  g245(.A(new_n667), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n663), .A2(new_n666), .A3(new_n668), .ZN(new_n672));
  OAI211_X1 g247(.A(new_n671), .B(new_n672), .C1(new_n669), .C2(new_n670), .ZN(new_n673));
  XOR2_X1   g248(.A(G1991), .B(G1996), .Z(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n678), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n679), .A2(new_n680), .ZN(G229));
  INV_X1    g256(.A(G16), .ZN(new_n682));
  AND2_X1   g257(.A1(new_n682), .A2(G6), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n683), .B1(G305), .B2(G16), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n686), .A2(G1981), .A3(new_n687), .ZN(new_n688));
  INV_X1    g263(.A(G1981), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  AOI211_X1 g265(.A(KEYINPUT32), .B(new_n683), .C1(G305), .C2(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n682), .A2(G23), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n694), .B1(G288), .B2(G16), .ZN(new_n695));
  INV_X1    g270(.A(KEYINPUT33), .ZN(new_n696));
  OR2_X1    g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  AOI211_X1 g272(.A(KEYINPUT33), .B(new_n694), .C1(G288), .C2(G16), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AOI21_X1  g274(.A(G1976), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  INV_X1    g276(.A(G1976), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n701), .A2(new_n698), .A3(new_n702), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g279(.A(KEYINPUT83), .B(G16), .Z(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n706), .A2(G22), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(G166), .B2(new_n706), .ZN(new_n708));
  XNOR2_X1  g283(.A(KEYINPUT84), .B(G1971), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  OAI211_X1 g286(.A(new_n709), .B(new_n707), .C1(G166), .C2(new_n706), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(new_n713), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n693), .A2(new_n704), .A3(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT85), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n713), .B1(new_n688), .B2(new_n692), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n718), .A2(KEYINPUT85), .A3(new_n704), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n717), .A2(KEYINPUT34), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(KEYINPUT34), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  INV_X1    g296(.A(G29), .ZN(new_n722));
  AND2_X1   g297(.A1(new_n722), .A2(G25), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n479), .A2(G119), .ZN(new_n724));
  OR2_X1    g299(.A1(new_n724), .A2(KEYINPUT82), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(KEYINPUT82), .ZN(new_n726));
  AOI22_X1  g301(.A1(new_n725), .A2(new_n726), .B1(G131), .B2(new_n474), .ZN(new_n727));
  OR2_X1    g302(.A1(G95), .A2(G2105), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n728), .B(G2104), .C1(G107), .C2(new_n458), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n723), .B1(new_n730), .B2(G29), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT35), .B(G1991), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n731), .B(new_n733), .ZN(new_n734));
  MUX2_X1   g309(.A(G24), .B(G290), .S(new_n705), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1986), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT86), .ZN(new_n739));
  NOR3_X1   g314(.A1(new_n721), .A2(new_n738), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT34), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n718), .A2(KEYINPUT85), .A3(new_n704), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT85), .B1(new_n718), .B2(new_n704), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g319(.A(KEYINPUT86), .B1(new_n744), .B2(new_n737), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n720), .B1(new_n740), .B2(new_n745), .ZN(new_n746));
  XOR2_X1   g321(.A(KEYINPUT87), .B(KEYINPUT36), .Z(new_n747));
  INV_X1    g322(.A(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT97), .ZN(new_n750));
  INV_X1    g325(.A(G35), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n750), .B1(new_n751), .B2(G29), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(G29), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n483), .B2(G29), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n752), .B1(new_n754), .B2(new_n750), .ZN(new_n755));
  XOR2_X1   g330(.A(KEYINPUT98), .B(KEYINPUT29), .Z(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n757), .A2(G2090), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n722), .A2(G27), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G164), .B2(new_n722), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n758), .B1(G2078), .B2(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(G2067), .ZN(new_n762));
  INV_X1    g337(.A(KEYINPUT28), .ZN(new_n763));
  INV_X1    g338(.A(G26), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n763), .B1(new_n764), .B2(G29), .ZN(new_n765));
  NOR2_X1   g340(.A1(new_n764), .A2(G29), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n474), .A2(G140), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n479), .A2(G128), .ZN(new_n768));
  NOR2_X1   g343(.A1(G104), .A2(G2105), .ZN(new_n769));
  OAI21_X1  g344(.A(G2104), .B1(new_n458), .B2(G116), .ZN(new_n770));
  OAI211_X1 g345(.A(new_n767), .B(new_n768), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(G29), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n765), .B1(new_n772), .B2(new_n763), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n773), .B(KEYINPUT91), .ZN(new_n774));
  AOI21_X1  g349(.A(new_n761), .B1(new_n762), .B2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(G5), .A2(G16), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G171), .B2(G16), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT96), .ZN(new_n778));
  XOR2_X1   g353(.A(new_n778), .B(G1961), .Z(new_n779));
  NOR2_X1   g354(.A1(new_n757), .A2(G2090), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT99), .ZN(new_n781));
  NOR2_X1   g356(.A1(new_n774), .A2(new_n762), .ZN(new_n782));
  AND2_X1   g357(.A1(new_n760), .A2(G2078), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n682), .A2(G4), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(new_n594), .B2(new_n682), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT88), .B(G1348), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR3_X1   g362(.A1(new_n782), .A2(new_n783), .A3(new_n787), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n775), .A2(new_n779), .A3(new_n781), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(G29), .A2(G32), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n479), .A2(G129), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n494), .A2(G105), .ZN(new_n792));
  INV_X1    g367(.A(G141), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n473), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT93), .B(KEYINPUT26), .ZN(new_n795));
  NAND3_X1  g370(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(new_n794), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n790), .B1(new_n798), .B2(G29), .ZN(new_n799));
  XOR2_X1   g374(.A(KEYINPUT27), .B(G1996), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n706), .A2(G19), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n547), .B2(new_n706), .ZN(new_n803));
  MUX2_X1   g378(.A(new_n802), .B(new_n803), .S(KEYINPUT89), .Z(new_n804));
  XNOR2_X1  g379(.A(KEYINPUT90), .B(G1341), .ZN(new_n805));
  XNOR2_X1  g380(.A(new_n804), .B(new_n805), .ZN(new_n806));
  NOR2_X1   g381(.A1(G29), .A2(G33), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n494), .A2(G103), .ZN(new_n808));
  XOR2_X1   g383(.A(new_n808), .B(KEYINPUT25), .Z(new_n809));
  NAND2_X1  g384(.A1(new_n474), .A2(G139), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n459), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n811));
  OAI211_X1 g386(.A(new_n809), .B(new_n810), .C1(new_n458), .C2(new_n811), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT92), .ZN(new_n813));
  AOI21_X1  g388(.A(new_n807), .B1(new_n813), .B2(G29), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n814), .A2(G2072), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n682), .A2(G21), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(G168), .B2(new_n682), .ZN(new_n817));
  NOR2_X1   g392(.A1(new_n817), .A2(G1966), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  OR2_X1    g394(.A1(KEYINPUT24), .A2(G34), .ZN(new_n820));
  NAND2_X1  g395(.A1(KEYINPUT24), .A2(G34), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(new_n722), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(G160), .B2(new_n722), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2084), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(G2072), .B2(new_n814), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n706), .A2(G20), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT100), .B(KEYINPUT23), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n828), .B1(G299), .B2(G16), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n829), .B(G1956), .ZN(new_n830));
  XOR2_X1   g405(.A(KEYINPUT31), .B(G11), .Z(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT94), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT30), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n833), .A2(G28), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n833), .A2(G28), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n834), .A2(new_n835), .A3(new_n722), .ZN(new_n836));
  OAI211_X1 g411(.A(new_n832), .B(new_n836), .C1(new_n618), .C2(new_n722), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(KEYINPUT95), .Z(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(new_n817), .B2(G1966), .ZN(new_n839));
  NAND4_X1  g414(.A1(new_n819), .A2(new_n825), .A3(new_n830), .A4(new_n839), .ZN(new_n840));
  NOR4_X1   g415(.A1(new_n789), .A2(new_n801), .A3(new_n806), .A4(new_n840), .ZN(new_n841));
  OAI211_X1 g416(.A(new_n720), .B(new_n747), .C1(new_n740), .C2(new_n745), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n749), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(G311));
  INV_X1    g419(.A(KEYINPUT101), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND4_X1  g421(.A1(new_n749), .A2(new_n841), .A3(KEYINPUT101), .A4(new_n842), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n846), .A2(new_n847), .ZN(G150));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n849));
  INV_X1    g424(.A(G67), .ZN(new_n850));
  AOI211_X1 g425(.A(new_n850), .B(new_n501), .C1(new_n503), .C2(new_n505), .ZN(new_n851));
  NAND2_X1  g426(.A1(G80), .A2(G543), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n849), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g429(.A(G67), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n855), .A2(KEYINPUT102), .A3(new_n852), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n854), .A2(G651), .A3(new_n856), .ZN(new_n857));
  INV_X1    g432(.A(G93), .ZN(new_n858));
  INV_X1    g433(.A(G55), .ZN(new_n859));
  OAI22_X1  g434(.A1(new_n511), .A2(new_n858), .B1(new_n859), .B2(new_n514), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n857), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n862), .A2(G860), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n863), .B(KEYINPUT37), .Z(new_n864));
  NOR2_X1   g439(.A1(new_n593), .A2(new_n601), .ZN(new_n865));
  XNOR2_X1  g440(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n865), .B(new_n866), .ZN(new_n867));
  AOI211_X1 g442(.A(new_n849), .B(new_n853), .C1(new_n506), .C2(G67), .ZN(new_n868));
  AOI21_X1  g443(.A(KEYINPUT102), .B1(new_n855), .B2(new_n852), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n868), .A2(new_n869), .A3(new_n508), .ZN(new_n870));
  OAI21_X1  g445(.A(KEYINPUT103), .B1(new_n870), .B2(new_n860), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT103), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n857), .A2(new_n872), .A3(new_n861), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n871), .A2(new_n547), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n533), .ZN(new_n875));
  NOR3_X1   g450(.A1(new_n539), .A2(new_n536), .A3(new_n508), .ZN(new_n876));
  AOI21_X1  g451(.A(KEYINPUT71), .B1(new_n545), .B2(G651), .ZN(new_n877));
  OAI211_X1 g452(.A(new_n875), .B(new_n534), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n878), .A2(KEYINPUT103), .A3(new_n862), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n874), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n867), .B(new_n880), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n864), .B1(new_n881), .B2(G860), .ZN(G145));
  XNOR2_X1  g457(.A(G160), .B(new_n618), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(G162), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n479), .A2(G130), .ZN(new_n885));
  OR2_X1    g460(.A1(G106), .A2(G2105), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n886), .B(G2104), .C1(G118), .C2(new_n458), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n474), .A2(G142), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(new_n890), .B1(new_n727), .B2(new_n729), .ZN(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT104), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n727), .A2(new_n729), .A3(new_n890), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  AND3_X1   g470(.A1(new_n727), .A2(new_n729), .A3(new_n890), .ZN(new_n896));
  OAI21_X1  g471(.A(KEYINPUT104), .B1(new_n896), .B2(new_n891), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n610), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n895), .A2(new_n897), .A3(new_n610), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n900), .A2(KEYINPUT105), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT105), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n610), .B1(new_n895), .B2(new_n897), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n798), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n813), .A2(new_n771), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n813), .A2(new_n771), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n908), .A2(new_n498), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n498), .B1(new_n908), .B2(new_n909), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n907), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n908), .A2(new_n909), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n913), .A2(G164), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n498), .A3(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n914), .A2(new_n798), .A3(new_n915), .ZN(new_n916));
  AND4_X1   g491(.A1(new_n902), .A2(new_n906), .A3(new_n912), .A4(new_n916), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n916), .A2(new_n912), .B1(new_n906), .B2(new_n902), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n884), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n912), .A2(new_n916), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(new_n904), .B2(new_n905), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n906), .A2(new_n912), .A3(new_n916), .A4(new_n902), .ZN(new_n922));
  INV_X1    g497(.A(new_n884), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(G37), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n919), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g502(.A(KEYINPUT107), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT106), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n880), .B(new_n603), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n558), .A2(new_n565), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n593), .ZN(new_n932));
  AND2_X1   g507(.A1(new_n592), .A2(new_n589), .ZN(new_n933));
  AOI22_X1  g508(.A1(new_n585), .A2(G651), .B1(G54), .B2(new_n522), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n933), .B(new_n934), .C1(new_n558), .C2(new_n565), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n932), .A2(KEYINPUT41), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT41), .B1(new_n932), .B2(new_n935), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n930), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n932), .A2(new_n935), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n930), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n929), .B1(new_n940), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n929), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n928), .B1(new_n943), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G166), .B(G288), .ZN(new_n947));
  INV_X1    g522(.A(G305), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n947), .A2(new_n948), .ZN(new_n950));
  OR3_X1    g525(.A1(new_n949), .A2(new_n950), .A3(G290), .ZN(new_n951));
  OAI21_X1  g526(.A(G290), .B1(new_n949), .B2(new_n950), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g528(.A(new_n953), .B(KEYINPUT42), .ZN(new_n954));
  INV_X1    g529(.A(new_n942), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT106), .B1(new_n955), .B2(new_n939), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n956), .A2(KEYINPUT107), .A3(new_n944), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n946), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n954), .ZN(new_n959));
  NAND4_X1  g534(.A1(new_n959), .A2(KEYINPUT107), .A3(new_n956), .A4(new_n944), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n958), .A2(G868), .A3(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(KEYINPUT108), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n862), .A2(new_n597), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n958), .A2(new_n964), .A3(G868), .A4(new_n960), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(G295));
  NAND3_X1  g541(.A1(new_n962), .A2(new_n963), .A3(new_n965), .ZN(G331));
  INV_X1    g542(.A(new_n953), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT109), .ZN(new_n969));
  NAND2_X1  g544(.A1(G171), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(G301), .A2(KEYINPUT109), .ZN(new_n971));
  NAND2_X1  g546(.A1(G286), .A2(new_n971), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n874), .A2(new_n972), .A3(new_n879), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n972), .B1(new_n874), .B2(new_n879), .ZN(new_n974));
  OAI21_X1  g549(.A(new_n970), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(new_n972), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n857), .A2(new_n872), .A3(new_n861), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n872), .B1(new_n857), .B2(new_n861), .ZN(new_n978));
  NOR3_X1   g553(.A1(new_n977), .A2(new_n978), .A3(new_n878), .ZN(new_n979));
  INV_X1    g554(.A(new_n879), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n976), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(new_n970), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n874), .A2(new_n972), .A3(new_n879), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n981), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AND3_X1   g559(.A1(new_n975), .A2(new_n984), .A3(new_n941), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n938), .B1(new_n975), .B2(new_n984), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n968), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(new_n938), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n973), .A2(new_n974), .A3(new_n970), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n982), .B1(new_n981), .B2(new_n983), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n975), .A2(new_n984), .A3(new_n941), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n991), .A2(new_n953), .A3(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n987), .A2(new_n993), .A3(new_n925), .ZN(new_n994));
  INV_X1    g569(.A(KEYINPUT43), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n997));
  NOR3_X1   g572(.A1(new_n936), .A2(new_n937), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n937), .A2(new_n997), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  AOI211_X1 g575(.A(new_n998), .B(new_n1000), .C1(new_n975), .C2(new_n984), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n968), .B1(new_n1001), .B2(new_n985), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1002), .A2(KEYINPUT43), .A3(new_n925), .A4(new_n993), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n996), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT44), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n985), .A2(new_n986), .ZN(new_n1007));
  AOI21_X1  g582(.A(G37), .B1(new_n1007), .B2(new_n953), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n995), .B1(new_n1008), .B2(new_n987), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n993), .A2(new_n925), .ZN(new_n1010));
  INV_X1    g585(.A(new_n998), .ZN(new_n1011));
  OAI211_X1 g586(.A(new_n1011), .B(new_n999), .C1(new_n989), .C2(new_n990), .ZN(new_n1012));
  AOI21_X1  g587(.A(new_n953), .B1(new_n1012), .B2(new_n992), .ZN(new_n1013));
  NOR3_X1   g588(.A1(new_n1010), .A2(new_n1013), .A3(KEYINPUT43), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1006), .B1(new_n1009), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT111), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1005), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1006), .B1(new_n996), .B2(new_n1003), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1002), .A2(new_n995), .A3(new_n925), .A4(new_n993), .ZN(new_n1020));
  AOI21_X1  g595(.A(KEYINPUT44), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1021));
  OAI21_X1  g596(.A(KEYINPUT111), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1017), .A2(new_n1022), .ZN(G397));
  INV_X1    g598(.A(KEYINPUT61), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n931), .B(KEYINPUT57), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  INV_X1    g601(.A(G1384), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n498), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(KEYINPUT119), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT119), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n498), .A2(new_n1030), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1029), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(G160), .A2(G40), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n498), .A2(new_n1027), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1033), .B1(KEYINPUT50), .B2(new_n1034), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G1956), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(G40), .ZN(new_n1039));
  AOI211_X1 g614(.A(new_n1039), .B(new_n462), .C1(new_n470), .C2(new_n471), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT45), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1034), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n498), .A2(KEYINPUT45), .A3(new_n1027), .ZN(new_n1043));
  XNOR2_X1  g618(.A(KEYINPUT56), .B(G2072), .ZN(new_n1044));
  AND4_X1   g619(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .A4(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1025), .B1(new_n1038), .B2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(G1956), .B1(new_n1032), .B2(new_n1035), .ZN(new_n1048));
  XNOR2_X1  g623(.A(G299), .B(KEYINPUT57), .ZN(new_n1049));
  NOR3_X1   g624(.A1(new_n1048), .A2(new_n1049), .A3(new_n1045), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1024), .B1(new_n1047), .B2(new_n1050), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(new_n762), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1034), .A2(KEYINPUT50), .ZN(new_n1054));
  AND3_X1   g629(.A1(new_n1054), .A2(new_n1040), .A3(new_n1028), .ZN(new_n1055));
  OAI211_X1 g630(.A(KEYINPUT60), .B(new_n1053), .C1(new_n1055), .C2(new_n786), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT123), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1056), .A2(new_n1057), .A3(new_n593), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1040), .A3(new_n1028), .ZN(new_n1059));
  INV_X1    g634(.A(new_n786), .ZN(new_n1060));
  AOI22_X1  g635(.A1(new_n1059), .A2(new_n1060), .B1(new_n762), .B2(new_n1052), .ZN(new_n1061));
  OR2_X1    g636(.A1(new_n1061), .A2(KEYINPUT60), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n594), .A2(KEYINPUT123), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n593), .A2(new_n1057), .ZN(new_n1064));
  NAND4_X1  g639(.A1(new_n1061), .A2(KEYINPUT60), .A3(new_n1063), .A4(new_n1064), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1058), .A2(new_n1062), .A3(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1038), .A2(new_n1025), .A3(new_n1046), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1049), .B1(new_n1048), .B2(new_n1045), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1067), .A2(KEYINPUT61), .A3(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1051), .A2(new_n1066), .A3(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1043), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT45), .B1(new_n498), .B2(new_n1027), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1071), .A2(new_n1033), .A3(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT121), .ZN(new_n1074));
  INV_X1    g649(.A(G1996), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1042), .A2(new_n1040), .A3(new_n1043), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT121), .B1(new_n1077), .B2(G1996), .ZN(new_n1078));
  XNOR2_X1  g653(.A(KEYINPUT122), .B(G1341), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT58), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1076), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n547), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1082), .A2(KEYINPUT59), .A3(new_n547), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1053), .B1(new_n1055), .B2(new_n786), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1088), .A2(new_n594), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1089), .A2(new_n1068), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT120), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1090), .A2(new_n1091), .A3(new_n1067), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1090), .B2(new_n1067), .ZN(new_n1093));
  OAI22_X1  g668(.A1(new_n1070), .A2(new_n1087), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT124), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n1097));
  INV_X1    g672(.A(G2078), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1042), .A2(new_n1098), .A3(new_n1040), .A4(new_n1043), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1099), .A2(KEYINPUT53), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(KEYINPUT53), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  XNOR2_X1  g677(.A(KEYINPUT125), .B(G1961), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1104), .B1(new_n1035), .B2(new_n1028), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1105), .ZN(new_n1106));
  AOI21_X1  g681(.A(G301), .B1(new_n1102), .B2(new_n1106), .ZN(new_n1107));
  AOI211_X1 g682(.A(G171), .B(new_n1105), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1097), .B1(new_n1107), .B2(new_n1108), .ZN(new_n1109));
  OAI221_X1 g684(.A(G8), .B1(new_n702), .B2(G288), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1110));
  INV_X1    g685(.A(G288), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1111), .A2(G1976), .ZN(new_n1112));
  OR3_X1    g687(.A1(new_n1110), .A2(KEYINPUT52), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n574), .ZN(new_n1114));
  AOI22_X1  g689(.A1(new_n1114), .A2(G651), .B1(G48), .B2(new_n522), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT118), .B(G86), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n521), .A2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n689), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT49), .ZN(new_n1119));
  NOR2_X1   g694(.A1(G305), .A2(G1981), .ZN(new_n1120));
  OR3_X1    g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(G8), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1052), .A2(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1119), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1121), .A2(new_n1123), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT117), .ZN(new_n1126));
  AND3_X1   g701(.A1(new_n1110), .A2(new_n1126), .A3(KEYINPUT52), .ZN(new_n1127));
  AOI21_X1  g702(.A(new_n1126), .B1(new_n1110), .B2(KEYINPUT52), .ZN(new_n1128));
  OAI211_X1 g703(.A(new_n1113), .B(new_n1125), .C1(new_n1127), .C2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(G303), .A2(G8), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT55), .ZN(new_n1132));
  XNOR2_X1  g707(.A(new_n1131), .B(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1133), .A2(KEYINPUT116), .ZN(new_n1134));
  XNOR2_X1  g709(.A(new_n1131), .B(KEYINPUT55), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT116), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1134), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G1971), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1077), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1140), .A2(KEYINPUT114), .ZN(new_n1141));
  INV_X1    g716(.A(G2090), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1055), .A2(KEYINPUT115), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1059), .B2(G2090), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT114), .ZN(new_n1146));
  NAND3_X1  g721(.A1(new_n1077), .A2(new_n1146), .A3(new_n1139), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1141), .A2(new_n1143), .A3(new_n1145), .A4(new_n1147), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1138), .A2(new_n1148), .A3(G8), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1140), .B1(new_n1036), .B2(G2090), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1133), .B1(new_n1150), .B2(G8), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1109), .A2(new_n1130), .A3(new_n1149), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1102), .A2(new_n1106), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G171), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1102), .A2(G301), .A3(new_n1106), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1155), .A2(KEYINPUT54), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(G2084), .ZN(new_n1158));
  INV_X1    g733(.A(G1966), .ZN(new_n1159));
  AOI22_X1  g734(.A1(new_n1055), .A2(new_n1158), .B1(new_n1077), .B2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(G286), .A2(G8), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(KEYINPUT51), .ZN(new_n1163));
  OAI211_X1 g738(.A(new_n1163), .B(new_n1161), .C1(new_n1160), .C2(new_n1122), .ZN(new_n1164));
  OAI22_X1  g739(.A1(new_n1073), .A2(G1966), .B1(new_n1059), .B2(G2084), .ZN(new_n1165));
  OAI211_X1 g740(.A(KEYINPUT51), .B(G8), .C1(new_n1165), .C2(G286), .ZN(new_n1166));
  AOI21_X1  g741(.A(new_n1162), .B1(new_n1164), .B2(new_n1166), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1157), .A2(new_n1168), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1153), .A2(new_n1169), .ZN(new_n1170));
  NOR2_X1   g745(.A1(new_n1061), .A2(new_n593), .ZN(new_n1171));
  OAI21_X1  g746(.A(new_n1067), .B1(new_n1047), .B2(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1172), .A2(KEYINPUT120), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1090), .A2(new_n1091), .A3(new_n1067), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1175), .B(KEYINPUT124), .C1(new_n1070), .C2(new_n1087), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1096), .A2(new_n1170), .A3(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(KEYINPUT62), .ZN(new_n1178));
  OAI21_X1  g753(.A(new_n1107), .B1(new_n1167), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g754(.A(KEYINPUT62), .B(new_n1162), .C1(new_n1164), .C2(new_n1166), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1130), .A2(new_n1149), .A3(new_n1152), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1138), .A2(new_n1148), .A3(G8), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT63), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1165), .A2(new_n1184), .A3(G8), .A4(G168), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1151), .A2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g761(.A(new_n1130), .B1(new_n1183), .B2(new_n1186), .ZN(new_n1187));
  AND3_X1   g762(.A1(new_n1125), .A2(new_n702), .A3(new_n1111), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n1123), .B1(new_n1188), .B2(new_n1120), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1133), .B1(new_n1148), .B2(G8), .ZN(new_n1190));
  NAND3_X1  g765(.A1(new_n1165), .A2(G8), .A3(G168), .ZN(new_n1191));
  NOR3_X1   g766(.A1(new_n1190), .A2(new_n1129), .A3(new_n1191), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1187), .B(new_n1189), .C1(new_n1192), .C2(new_n1184), .ZN(new_n1193));
  NOR2_X1   g768(.A1(new_n1182), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1177), .A2(new_n1194), .ZN(new_n1195));
  NOR2_X1   g770(.A1(new_n1042), .A2(new_n1033), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1196), .A2(new_n1075), .ZN(new_n1197));
  XOR2_X1   g772(.A(new_n1197), .B(KEYINPUT113), .Z(new_n1198));
  XNOR2_X1  g773(.A(new_n771), .B(new_n762), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1199), .B1(new_n798), .B2(new_n1075), .ZN(new_n1200));
  AOI22_X1  g775(.A1(new_n1198), .A2(new_n798), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NOR2_X1   g776(.A1(new_n730), .A2(new_n732), .ZN(new_n1202));
  AOI21_X1  g777(.A(new_n733), .B1(new_n727), .B2(new_n729), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1196), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  AND2_X1   g779(.A1(new_n1201), .A2(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(new_n1196), .ZN(new_n1206));
  OR3_X1    g781(.A1(new_n1206), .A2(G1986), .A3(G290), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1196), .A2(G1986), .A3(G290), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  XNOR2_X1  g784(.A(new_n1209), .B(KEYINPUT112), .ZN(new_n1210));
  AND2_X1   g785(.A1(new_n1205), .A2(new_n1210), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1195), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT46), .ZN(new_n1213));
  XNOR2_X1  g788(.A(new_n1198), .B(new_n1213), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1199), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1196), .B1(new_n1215), .B2(new_n907), .ZN(new_n1216));
  NAND2_X1  g791(.A1(new_n1214), .A2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g792(.A(new_n1217), .B(KEYINPUT47), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1219));
  OAI21_X1  g794(.A(new_n1219), .B1(G2067), .B2(new_n771), .ZN(new_n1220));
  XNOR2_X1  g795(.A(new_n1207), .B(KEYINPUT48), .ZN(new_n1221));
  AOI22_X1  g796(.A1(new_n1220), .A2(new_n1196), .B1(new_n1205), .B2(new_n1221), .ZN(new_n1222));
  AND2_X1   g797(.A1(new_n1218), .A2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g798(.A1(new_n1212), .A2(new_n1223), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g799(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1226));
  NAND3_X1  g800(.A1(new_n645), .A2(G319), .A3(new_n660), .ZN(new_n1227));
  INV_X1    g801(.A(KEYINPUT126), .ZN(new_n1228));
  OAI22_X1  g802(.A1(new_n1227), .A2(new_n1228), .B1(new_n679), .B2(new_n680), .ZN(new_n1229));
  AND2_X1   g803(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1230));
  NOR2_X1   g804(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g805(.A1(new_n1226), .A2(new_n926), .A3(new_n1231), .ZN(G225));
  NAND2_X1  g806(.A1(G225), .A2(KEYINPUT127), .ZN(new_n1233));
  INV_X1    g807(.A(KEYINPUT127), .ZN(new_n1234));
  NAND4_X1  g808(.A1(new_n1226), .A2(new_n926), .A3(new_n1231), .A4(new_n1234), .ZN(new_n1235));
  NAND2_X1  g809(.A1(new_n1233), .A2(new_n1235), .ZN(G308));
endmodule


