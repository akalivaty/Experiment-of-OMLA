//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n576, new_n577, new_n579, new_n580, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n598, new_n599, new_n600, new_n602, new_n603,
    new_n604, new_n605, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n660, new_n661, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n869, new_n870,
    new_n871, new_n872, new_n873, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053, new_n1054, new_n1055,
    new_n1056, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1156, new_n1157, new_n1158, new_n1159,
    new_n1160, new_n1161, new_n1162, new_n1163, new_n1164, new_n1165,
    new_n1166, new_n1167, new_n1168, new_n1169, new_n1170, new_n1171,
    new_n1172, new_n1173, new_n1174, new_n1175, new_n1176, new_n1177,
    new_n1178, new_n1179, new_n1180, new_n1181, new_n1182, new_n1183,
    new_n1184, new_n1185, new_n1186, new_n1187, new_n1188, new_n1189,
    new_n1190, new_n1191, new_n1192, new_n1193, new_n1194, new_n1195,
    new_n1196, new_n1197, new_n1198, new_n1199, new_n1200, new_n1201,
    new_n1202, new_n1203, new_n1204, new_n1205, new_n1206, new_n1207,
    new_n1208, new_n1209, new_n1210, new_n1211, new_n1212, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1217, new_n1218, new_n1219,
    new_n1220, new_n1221, new_n1222, new_n1223, new_n1224, new_n1225,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1230, new_n1231,
    new_n1232, new_n1233, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1243,
    new_n1244, new_n1245, new_n1246, new_n1247, new_n1248, new_n1249,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1254, new_n1255,
    new_n1256, new_n1257, new_n1258, new_n1259, new_n1260, new_n1261,
    new_n1262, new_n1263, new_n1264, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1270, new_n1271, new_n1272, new_n1273,
    new_n1274, new_n1275, new_n1276, new_n1277, new_n1278, new_n1279,
    new_n1280, new_n1281, new_n1282, new_n1283, new_n1284, new_n1285,
    new_n1286, new_n1287, new_n1288, new_n1289, new_n1290, new_n1291,
    new_n1292, new_n1293, new_n1294, new_n1295, new_n1296, new_n1297,
    new_n1298, new_n1299, new_n1300, new_n1301, new_n1302, new_n1303,
    new_n1304, new_n1305, new_n1306, new_n1307, new_n1308, new_n1309,
    new_n1310, new_n1311, new_n1312, new_n1313, new_n1314, new_n1315,
    new_n1316, new_n1317, new_n1318, new_n1319, new_n1320, new_n1321,
    new_n1324, new_n1325, new_n1326, new_n1327, new_n1329;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  INV_X1    g017(.A(G2072), .ZN(new_n443));
  INV_X1    g018(.A(G2078), .ZN(new_n444));
  NOR2_X1   g019(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND3_X1  g020(.A1(new_n445), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  NOR4_X1   g030(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT67), .Z(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n455), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n455), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND3_X1   g037(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(KEYINPUT3), .B1(KEYINPUT68), .B2(G2104), .ZN(new_n464));
  OAI211_X1 g039(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n465));
  NAND3_X1  g040(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  AND2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n469));
  OAI21_X1  g044(.A(G125), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(new_n462), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n467), .A2(new_n472), .ZN(G160));
  NOR2_X1   g048(.A1(new_n462), .A2(G112), .ZN(new_n474));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT68), .A2(G2104), .ZN(new_n477));
  INV_X1    g052(.A(KEYINPUT3), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g054(.A1(KEYINPUT68), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n480));
  AOI21_X1  g055(.A(G2105), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  AOI21_X1  g056(.A(new_n476), .B1(new_n481), .B2(G136), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n462), .B1(new_n479), .B2(new_n480), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G124), .ZN(new_n485));
  INV_X1    g060(.A(KEYINPUT69), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n484), .A2(KEYINPUT69), .A3(G124), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(G162));
  OR2_X1    g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR3_X1   g068(.A1(new_n493), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n462), .A2(G138), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n496), .B1(new_n479), .B2(new_n480), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n462), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g077(.A(new_n502), .B1(new_n484), .B2(G126), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(G164));
  XNOR2_X1  g080(.A(KEYINPUT6), .B(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  NOR2_X1   g083(.A1(KEYINPUT5), .A2(G543), .ZN(new_n509));
  AND2_X1   g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n509), .A2(new_n510), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G88), .ZN(new_n514));
  OAI22_X1  g089(.A1(new_n507), .A2(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g094(.A1(KEYINPUT5), .A2(G543), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G62), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  AOI21_X1  g098(.A(new_n516), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n515), .A2(new_n524), .ZN(G166));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OR2_X1    g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  NAND2_X1  g102(.A1(KEYINPUT6), .A2(G651), .ZN(new_n528));
  AOI21_X1  g103(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n518), .B1(new_n527), .B2(new_n528), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT70), .B(G51), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT7), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(KEYINPUT71), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT71), .ZN(new_n538));
  NAND4_X1  g113(.A1(new_n538), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n539));
  AOI21_X1  g114(.A(new_n535), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AND3_X1   g115(.A1(new_n537), .A2(new_n535), .A3(new_n539), .ZN(new_n541));
  OAI211_X1 g116(.A(new_n531), .B(new_n534), .C1(new_n540), .C2(new_n541), .ZN(G286));
  INV_X1    g117(.A(G286), .ZN(G168));
  NAND3_X1  g118(.A1(new_n521), .A2(new_n506), .A3(G90), .ZN(new_n544));
  OAI211_X1 g119(.A(G52), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n544), .A2(KEYINPUT73), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  AOI21_X1  g122(.A(KEYINPUT73), .B1(new_n544), .B2(new_n545), .ZN(new_n548));
  OAI21_X1  g123(.A(G64), .B1(new_n510), .B2(new_n509), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(KEYINPUT72), .B1(new_n551), .B2(G651), .ZN(new_n552));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n553));
  AOI211_X1 g128(.A(new_n553), .B(new_n516), .C1(new_n549), .C2(new_n550), .ZN(new_n554));
  OAI22_X1  g129(.A1(new_n547), .A2(new_n548), .B1(new_n552), .B2(new_n554), .ZN(G301));
  INV_X1    g130(.A(G301), .ZN(G171));
  OAI211_X1 g131(.A(G43), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n557));
  XNOR2_X1  g132(.A(KEYINPUT74), .B(G81), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n557), .B1(new_n513), .B2(new_n558), .ZN(new_n559));
  OAI21_X1  g134(.A(G56), .B1(new_n510), .B2(new_n509), .ZN(new_n560));
  NAND2_X1  g135(.A1(G68), .A2(G543), .ZN(new_n561));
  AOI21_X1  g136(.A(new_n516), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI21_X1  g137(.A(KEYINPUT75), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(G56), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n564), .B1(new_n519), .B2(new_n520), .ZN(new_n565));
  INV_X1    g140(.A(new_n561), .ZN(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  XOR2_X1   g143(.A(KEYINPUT74), .B(G81), .Z(new_n569));
  NAND3_X1  g144(.A1(new_n569), .A2(new_n521), .A3(new_n506), .ZN(new_n570));
  NAND4_X1  g145(.A1(new_n567), .A2(new_n568), .A3(new_n570), .A4(new_n557), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n563), .A2(new_n571), .ZN(new_n572));
  INV_X1    g147(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G860), .ZN(G153));
  NAND4_X1  g149(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g150(.A1(G1), .A2(G3), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT8), .ZN(new_n577));
  NAND4_X1  g152(.A1(G319), .A2(G483), .A3(G661), .A4(new_n577), .ZN(G188));
  AOI22_X1  g153(.A1(new_n521), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n579), .A2(new_n516), .ZN(new_n580));
  OAI211_X1 g155(.A(G53), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n581));
  OAI21_X1  g156(.A(KEYINPUT77), .B1(new_n581), .B2(KEYINPUT9), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT9), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n532), .A2(new_n583), .A3(new_n584), .A4(G53), .ZN(new_n585));
  AND2_X1   g160(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n581), .A2(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n587), .A2(KEYINPUT76), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT76), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n581), .A2(new_n589), .A3(KEYINPUT9), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n580), .B1(new_n586), .B2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT78), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n513), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g169(.A1(new_n521), .A2(new_n506), .A3(KEYINPUT78), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n594), .A2(G91), .A3(new_n595), .ZN(new_n596));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g173(.A1(new_n594), .A2(KEYINPUT79), .A3(G91), .A4(new_n595), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n592), .A2(new_n600), .ZN(G299));
  NAND2_X1  g176(.A1(new_n522), .A2(new_n523), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  AOI22_X1  g178(.A1(new_n527), .A2(new_n528), .B1(new_n519), .B2(new_n520), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G88), .B1(new_n532), .B2(G50), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n605), .ZN(G303));
  NAND3_X1  g181(.A1(new_n506), .A2(G49), .A3(G543), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n532), .A2(KEYINPUT80), .A3(G49), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND3_X1  g186(.A1(new_n594), .A2(G87), .A3(new_n595), .ZN(new_n612));
  OAI21_X1  g187(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(G288));
  NAND2_X1  g189(.A1(G73), .A2(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(KEYINPUT81), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n615), .A2(KEYINPUT81), .ZN(new_n617));
  NOR2_X1   g192(.A1(new_n510), .A2(new_n509), .ZN(new_n618));
  INV_X1    g193(.A(G61), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n620), .A2(G651), .B1(G48), .B2(new_n532), .ZN(new_n621));
  NAND3_X1  g196(.A1(new_n594), .A2(G86), .A3(new_n595), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n621), .A2(new_n622), .ZN(G305));
  AOI22_X1  g198(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n624), .A2(new_n516), .ZN(new_n625));
  INV_X1    g200(.A(G47), .ZN(new_n626));
  INV_X1    g201(.A(G85), .ZN(new_n627));
  OAI22_X1  g202(.A1(new_n507), .A2(new_n626), .B1(new_n513), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g203(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g204(.A(new_n629), .ZN(G290));
  NAND2_X1  g205(.A1(G301), .A2(G868), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n594), .A2(G92), .A3(new_n595), .ZN(new_n632));
  INV_X1    g207(.A(KEYINPUT10), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g209(.A1(new_n594), .A2(KEYINPUT10), .A3(G92), .A4(new_n595), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n637));
  INV_X1    g212(.A(G66), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n638), .A2(KEYINPUT82), .ZN(new_n639));
  INV_X1    g214(.A(KEYINPUT82), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G66), .ZN(new_n641));
  OAI211_X1 g216(.A(new_n639), .B(new_n641), .C1(new_n510), .C2(new_n509), .ZN(new_n642));
  NAND2_X1  g217(.A1(G79), .A2(G543), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n516), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n506), .A2(G54), .A3(G543), .ZN(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n637), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(KEYINPUT82), .B(G66), .ZN(new_n648));
  AOI22_X1  g223(.A1(new_n521), .A2(new_n648), .B1(G79), .B2(G543), .ZN(new_n649));
  OAI211_X1 g224(.A(KEYINPUT83), .B(new_n645), .C1(new_n649), .C2(new_n516), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n636), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT84), .ZN(new_n653));
  AOI22_X1  g228(.A1(new_n634), .A2(new_n635), .B1(new_n647), .B2(new_n650), .ZN(new_n654));
  INV_X1    g229(.A(KEYINPUT84), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  AND2_X1   g231(.A1(new_n653), .A2(new_n656), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n631), .B1(new_n657), .B2(G868), .ZN(G284));
  XNOR2_X1  g233(.A(G284), .B(KEYINPUT85), .ZN(G321));
  INV_X1    g234(.A(G868), .ZN(new_n660));
  NAND2_X1  g235(.A1(G299), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g236(.A(new_n661), .B1(new_n660), .B2(G168), .ZN(G297));
  OAI21_X1  g237(.A(new_n661), .B1(new_n660), .B2(G168), .ZN(G280));
  INV_X1    g238(.A(G559), .ZN(new_n664));
  OAI21_X1  g239(.A(new_n657), .B1(new_n664), .B2(G860), .ZN(G148));
  NAND3_X1  g240(.A1(new_n653), .A2(new_n664), .A3(new_n656), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n666), .A2(KEYINPUT86), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  INV_X1    g243(.A(KEYINPUT86), .ZN(new_n669));
  NAND4_X1  g244(.A1(new_n653), .A2(new_n656), .A3(new_n669), .A4(new_n664), .ZN(new_n670));
  INV_X1    g245(.A(new_n670), .ZN(new_n671));
  OAI21_X1  g246(.A(G868), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g247(.A(new_n672), .B1(G868), .B2(new_n573), .ZN(G323));
  XNOR2_X1  g248(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g249(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT12), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n676), .B(KEYINPUT13), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G2100), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n481), .A2(G135), .ZN(new_n679));
  NAND2_X1  g254(.A1(new_n484), .A2(G123), .ZN(new_n680));
  NOR2_X1   g255(.A1(new_n462), .A2(G111), .ZN(new_n681));
  OAI21_X1  g256(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n682));
  OAI211_X1 g257(.A(new_n679), .B(new_n680), .C1(new_n681), .C2(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(new_n683), .B(G2096), .Z(new_n684));
  NAND2_X1  g259(.A1(new_n678), .A2(new_n684), .ZN(G156));
  XNOR2_X1  g260(.A(KEYINPUT15), .B(G2435), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT87), .B(G2438), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G2427), .B(G2430), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n689), .ZN(new_n691));
  NAND3_X1  g266(.A1(new_n690), .A2(KEYINPUT14), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2451), .B(G2454), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT16), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1341), .B(G1348), .ZN(new_n695));
  XOR2_X1   g270(.A(new_n694), .B(new_n695), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n692), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G2443), .B(G2446), .ZN(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  AND2_X1   g274(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(G14), .B1(new_n697), .B2(new_n699), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(new_n701), .ZN(G401));
  XOR2_X1   g277(.A(G2084), .B(G2090), .Z(new_n703));
  XNOR2_X1  g278(.A(G2072), .B(G2078), .ZN(new_n704));
  XNOR2_X1  g279(.A(G2067), .B(G2678), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n706), .B(KEYINPUT18), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n704), .B(KEYINPUT17), .Z(new_n708));
  INV_X1    g283(.A(new_n703), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n709), .A2(new_n705), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n707), .B1(new_n708), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n705), .B1(new_n704), .B2(KEYINPUT88), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(KEYINPUT88), .B2(new_n704), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n713), .A2(KEYINPUT89), .A3(new_n709), .ZN(new_n714));
  INV_X1    g289(.A(new_n705), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n708), .ZN(new_n716));
  AOI21_X1  g291(.A(KEYINPUT89), .B1(new_n713), .B2(new_n709), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  XOR2_X1   g293(.A(G2096), .B(G2100), .Z(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(G227));
  XNOR2_X1  g295(.A(G1981), .B(G1986), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1971), .B(G1976), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT19), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  XOR2_X1   g300(.A(G1956), .B(G2474), .Z(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT90), .ZN(new_n727));
  XOR2_X1   g302(.A(G1961), .B(G1966), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT20), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n731));
  OR2_X1    g306(.A1(new_n727), .A2(new_n728), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI211_X1 g308(.A(new_n730), .B(new_n733), .C1(new_n724), .C2(new_n732), .ZN(new_n734));
  XOR2_X1   g309(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT91), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n734), .B(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(G1991), .B(G1996), .Z(new_n738));
  INV_X1    g313(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n737), .A2(new_n739), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n722), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n737), .A2(new_n739), .ZN(new_n744));
  NAND3_X1  g319(.A1(new_n744), .A2(new_n721), .A3(new_n740), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  INV_X1    g321(.A(new_n746), .ZN(G229));
  NAND2_X1  g322(.A1(G301), .A2(G16), .ZN(new_n748));
  INV_X1    g323(.A(G16), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G5), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G1961), .ZN(new_n752));
  NOR2_X1   g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n749), .A2(G21), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G168), .B2(new_n749), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n755), .A2(G1966), .ZN(new_n756));
  INV_X1    g331(.A(G28), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n757), .A2(KEYINPUT30), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(KEYINPUT30), .ZN(new_n759));
  OR2_X1    g334(.A1(KEYINPUT31), .A2(G11), .ZN(new_n760));
  NAND2_X1  g335(.A1(KEYINPUT31), .A2(G11), .ZN(new_n761));
  AOI22_X1  g336(.A1(new_n758), .A2(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g337(.A(G29), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n762), .B1(new_n683), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n755), .B2(G1966), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n756), .A2(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(KEYINPUT104), .B1(new_n753), .B2(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(new_n751), .A2(new_n752), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT104), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n768), .A2(new_n769), .A3(new_n756), .A4(new_n765), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n492), .A2(G127), .ZN(new_n771));
  AND2_X1   g346(.A1(G115), .A2(G2104), .ZN(new_n772));
  OAI21_X1  g347(.A(G2105), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n481), .A2(G139), .ZN(new_n774));
  NAND3_X1  g349(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT25), .Z(new_n776));
  AND3_X1   g351(.A1(new_n774), .A2(new_n776), .A3(KEYINPUT100), .ZN(new_n777));
  AOI21_X1  g352(.A(KEYINPUT100), .B1(new_n776), .B2(new_n774), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n773), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n779), .A2(G29), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n763), .A2(G33), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n780), .A2(new_n443), .A3(new_n781), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n443), .B1(new_n780), .B2(new_n781), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n763), .A2(G27), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G164), .B2(new_n763), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n785), .B(G2078), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT101), .B(KEYINPUT24), .ZN(new_n787));
  INV_X1    g362(.A(G34), .ZN(new_n788));
  AND2_X1   g363(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n763), .B1(new_n787), .B2(new_n788), .ZN(new_n790));
  OAI22_X1  g365(.A1(G160), .A2(new_n763), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2084), .ZN(new_n792));
  NOR3_X1   g367(.A1(new_n783), .A2(new_n786), .A3(new_n792), .ZN(new_n793));
  AND4_X1   g368(.A1(new_n767), .A2(new_n770), .A3(new_n782), .A4(new_n793), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n487), .A2(new_n488), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n763), .B1(new_n795), .B2(new_n482), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n763), .A2(G35), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(KEYINPUT29), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT29), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n800), .B(new_n797), .C1(G162), .C2(new_n763), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n802), .A2(G2090), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n749), .A2(G20), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(KEYINPUT23), .Z(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G299), .B2(G16), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n806), .A2(G1956), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(G1956), .ZN(new_n808));
  OAI21_X1  g383(.A(new_n803), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT105), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  OAI211_X1 g386(.A(KEYINPUT105), .B(new_n803), .C1(new_n807), .C2(new_n808), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(KEYINPUT99), .B(KEYINPUT28), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n763), .A2(G26), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  OAI21_X1  g391(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n817));
  INV_X1    g392(.A(G116), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n817), .B1(new_n818), .B2(G2105), .ZN(new_n819));
  AOI21_X1  g394(.A(new_n819), .B1(new_n484), .B2(G128), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n481), .A2(G140), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g397(.A(new_n816), .B1(new_n822), .B2(G29), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G2067), .ZN(new_n824));
  NAND3_X1  g399(.A1(new_n748), .A2(new_n752), .A3(new_n750), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n749), .A2(G19), .ZN(new_n826));
  XNOR2_X1  g401(.A(KEYINPUT98), .B(G1341), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n826), .B(new_n827), .C1(new_n573), .C2(new_n749), .ZN(new_n828));
  INV_X1    g403(.A(new_n827), .ZN(new_n829));
  AOI21_X1  g404(.A(new_n749), .B1(new_n563), .B2(new_n571), .ZN(new_n830));
  INV_X1    g405(.A(new_n826), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AND4_X1   g407(.A1(new_n824), .A2(new_n825), .A3(new_n828), .A4(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(KEYINPUT103), .A2(KEYINPUT26), .ZN(new_n834));
  NAND2_X1  g409(.A1(KEYINPUT103), .A2(KEYINPUT26), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n837));
  INV_X1    g412(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n834), .A2(new_n837), .A3(new_n835), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n484), .A2(G129), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n462), .A2(G105), .A3(G2104), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n841), .A2(new_n842), .A3(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n481), .A2(G141), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n846), .A2(KEYINPUT102), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT102), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n481), .A2(new_n848), .A3(G141), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n847), .A2(new_n849), .ZN(new_n850));
  AOI21_X1  g425(.A(new_n763), .B1(new_n845), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n763), .A2(G32), .ZN(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(KEYINPUT27), .B1(new_n851), .B2(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(KEYINPUT27), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n844), .B1(new_n847), .B2(new_n849), .ZN(new_n856));
  OAI211_X1 g431(.A(new_n855), .B(new_n852), .C1(new_n856), .C2(new_n763), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n854), .A2(new_n857), .A3(G1996), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n854), .A2(new_n857), .ZN(new_n859));
  INV_X1    g434(.A(G1996), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G2090), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n799), .A2(new_n862), .A3(new_n801), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n833), .A2(new_n858), .A3(new_n861), .A4(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n749), .A2(G4), .ZN(new_n865));
  OAI21_X1  g440(.A(new_n865), .B1(new_n657), .B2(new_n749), .ZN(new_n866));
  XNOR2_X1  g441(.A(KEYINPUT97), .B(G1348), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  OAI211_X1 g444(.A(new_n869), .B(new_n865), .C1(new_n657), .C2(new_n749), .ZN(new_n870));
  AOI21_X1  g445(.A(new_n864), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n794), .A2(new_n813), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(KEYINPUT95), .A2(KEYINPUT36), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT96), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n749), .A2(G24), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n875), .B1(new_n629), .B2(new_n749), .ZN(new_n876));
  XOR2_X1   g451(.A(new_n876), .B(G1986), .Z(new_n877));
  OR2_X1    g452(.A1(G25), .A2(G29), .ZN(new_n878));
  XOR2_X1   g453(.A(KEYINPUT35), .B(G1991), .Z(new_n879));
  INV_X1    g454(.A(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n481), .A2(G131), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n484), .A2(G119), .ZN(new_n882));
  OR2_X1    g457(.A1(G95), .A2(G2105), .ZN(new_n883));
  OAI211_X1 g458(.A(new_n883), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n881), .A2(new_n882), .A3(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(KEYINPUT92), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n878), .B(new_n880), .C1(new_n886), .C2(new_n763), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n878), .B1(new_n886), .B2(new_n763), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n888), .A2(new_n879), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n877), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  XOR2_X1   g465(.A(KEYINPUT32), .B(G1981), .Z(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(KEYINPUT93), .ZN(new_n893));
  INV_X1    g468(.A(new_n622), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n615), .B(KEYINPUT81), .ZN(new_n895));
  AOI21_X1  g470(.A(new_n619), .B1(new_n519), .B2(new_n520), .ZN(new_n896));
  OAI21_X1  g471(.A(G651), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n532), .A2(G48), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  OAI21_X1  g474(.A(G16), .B1(new_n894), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n749), .A2(G6), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n893), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n749), .B1(new_n621), .B2(new_n622), .ZN(new_n903));
  INV_X1    g478(.A(new_n901), .ZN(new_n904));
  NOR3_X1   g479(.A1(new_n903), .A2(KEYINPUT93), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n892), .B1(new_n902), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n900), .A2(new_n893), .A3(new_n901), .ZN(new_n907));
  OAI21_X1  g482(.A(KEYINPUT93), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n908), .A3(new_n891), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n906), .A2(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G1971), .ZN(new_n911));
  OAI21_X1  g486(.A(G16), .B1(new_n515), .B2(new_n524), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT94), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n749), .A2(G22), .ZN(new_n914));
  AND3_X1   g489(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n911), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(G288), .A2(G16), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n749), .A2(G23), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  XNOR2_X1  g495(.A(KEYINPUT33), .B(G1976), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n749), .B1(new_n603), .B2(new_n605), .ZN(new_n925));
  INV_X1    g500(.A(new_n914), .ZN(new_n926));
  OAI21_X1  g501(.A(KEYINPUT94), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n928), .A3(G1971), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n917), .A2(new_n923), .A3(new_n924), .A4(new_n929), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n910), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT34), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n890), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT34), .B1(new_n910), .B2(new_n930), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n874), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(new_n930), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n907), .A2(new_n908), .A3(new_n891), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n891), .B1(new_n907), .B2(new_n908), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n932), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n890), .ZN(new_n941));
  AND4_X1   g516(.A1(new_n874), .A2(new_n940), .A3(new_n934), .A4(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n873), .B1(new_n935), .B2(new_n942), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n940), .A2(new_n934), .A3(new_n941), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n944), .A2(KEYINPUT96), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n933), .A2(new_n874), .A3(new_n934), .ZN(new_n946));
  INV_X1    g521(.A(new_n873), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n872), .B1(new_n943), .B2(new_n948), .ZN(G311));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n943), .A2(new_n948), .ZN(new_n951));
  INV_X1    g526(.A(new_n872), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n950), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI211_X1 g528(.A(KEYINPUT106), .B(new_n872), .C1(new_n943), .C2(new_n948), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(G150));
  OAI211_X1 g530(.A(G55), .B(G543), .C1(new_n511), .C2(new_n512), .ZN(new_n956));
  INV_X1    g531(.A(G93), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n956), .B1(new_n513), .B2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n959));
  INV_X1    g534(.A(G67), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n519), .B2(new_n520), .ZN(new_n961));
  AND2_X1   g536(.A1(G80), .A2(G543), .ZN(new_n962));
  OAI21_X1  g537(.A(G651), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n958), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  OAI211_X1 g539(.A(KEYINPUT107), .B(G651), .C1(new_n961), .C2(new_n962), .ZN(new_n965));
  AOI22_X1  g540(.A1(new_n964), .A2(new_n965), .B1(new_n563), .B2(new_n571), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n963), .A2(new_n959), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n604), .A2(G93), .B1(new_n532), .B2(G55), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n967), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n559), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(new_n567), .ZN(new_n971));
  NOR2_X1   g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(new_n966), .A2(new_n972), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n973), .B(KEYINPUT38), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n657), .A2(G559), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n974), .A2(G559), .A3(new_n657), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT39), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n979), .A2(G860), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n977), .A2(KEYINPUT39), .A3(new_n978), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g558(.A1(new_n981), .A2(new_n982), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n980), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n969), .A2(G860), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n986), .B(KEYINPUT37), .ZN(new_n987));
  INV_X1    g562(.A(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT109), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n985), .A2(KEYINPUT109), .A3(new_n988), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(G145));
  AOI22_X1  g568(.A1(G130), .A2(new_n484), .B1(new_n481), .B2(G142), .ZN(new_n994));
  OAI21_X1  g569(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n995));
  INV_X1    g570(.A(G118), .ZN(new_n996));
  AOI22_X1  g571(.A1(new_n995), .A2(KEYINPUT111), .B1(new_n996), .B2(G2105), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n997), .B1(KEYINPUT111), .B2(new_n995), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n994), .A2(new_n998), .ZN(new_n999));
  XOR2_X1   g574(.A(new_n999), .B(new_n676), .Z(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n856), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1002), .A2(new_n779), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1002), .A2(new_n779), .ZN(new_n1005));
  NOR3_X1   g580(.A1(new_n1001), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(new_n1006), .ZN(new_n1007));
  XNOR2_X1  g582(.A(new_n504), .B(new_n822), .ZN(new_n1008));
  XNOR2_X1  g583(.A(new_n1008), .B(new_n886), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n1001), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1009), .ZN(new_n1012));
  INV_X1    g587(.A(new_n1010), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1012), .B1(new_n1013), .B2(new_n1006), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(G160), .B(KEYINPUT110), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(new_n683), .ZN(new_n1017));
  XNOR2_X1  g592(.A(new_n1017), .B(G162), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(G37), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1015), .A2(new_n1018), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1019), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT40), .ZN(G395));
  AOI21_X1  g598(.A(new_n973), .B1(new_n667), .B2(new_n670), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n667), .A2(new_n670), .A3(new_n973), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G299), .A2(new_n652), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT41), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n654), .A2(new_n600), .A3(new_n592), .ZN(new_n1029));
  AND3_X1   g604(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1028), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1031));
  OAI211_X1 g606(.A(new_n1025), .B(new_n1026), .C1(new_n1030), .C2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1026), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n1034), .B1(new_n1035), .B2(new_n1024), .ZN(new_n1036));
  XNOR2_X1  g611(.A(G288), .B(G305), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n629), .B(G166), .ZN(new_n1038));
  XNOR2_X1  g613(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  XNOR2_X1  g614(.A(new_n1039), .B(KEYINPUT42), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1032), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1040), .B1(new_n1032), .B2(new_n1036), .ZN(new_n1042));
  OAI21_X1  g617(.A(G868), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n969), .A2(new_n660), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(G295));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1043), .A2(new_n1046), .A3(new_n1044), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1040), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1033), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1035), .A2(new_n1024), .A3(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1048), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1032), .A2(new_n1036), .A3(new_n1040), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n660), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1044), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT112), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1047), .A2(new_n1056), .ZN(G331));
  XOR2_X1   g632(.A(KEYINPUT113), .B(KEYINPUT44), .Z(new_n1058));
  INV_X1    g633(.A(G90), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n545), .B1(new_n513), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT73), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n546), .ZN(new_n1063));
  INV_X1    g638(.A(new_n550), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1064), .B1(new_n521), .B2(G64), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n553), .B1(new_n1065), .B2(new_n516), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n551), .A2(KEYINPUT72), .A3(G651), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AND3_X1   g643(.A1(new_n1063), .A2(G286), .A3(new_n1068), .ZN(new_n1069));
  AOI21_X1  g644(.A(G286), .B1(new_n1063), .B2(new_n1068), .ZN(new_n1070));
  OAI22_X1  g645(.A1(new_n1069), .A2(new_n1070), .B1(new_n966), .B2(new_n972), .ZN(new_n1071));
  NAND2_X1  g646(.A1(G301), .A2(G168), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n572), .A2(new_n969), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n964), .A2(new_n567), .A3(new_n970), .A4(new_n965), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1063), .A2(new_n1068), .A3(G286), .ZN(new_n1075));
  NAND4_X1  g650(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1077), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1071), .A2(new_n1076), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1034), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1078), .A2(new_n1039), .A3(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1033), .B1(new_n1076), .B2(new_n1071), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1079), .B1(new_n1030), .B2(KEYINPUT115), .ZN(new_n1083));
  NOR2_X1   g658(.A1(G299), .A2(new_n652), .ZN(new_n1084));
  AOI22_X1  g659(.A1(new_n592), .A2(new_n600), .B1(new_n636), .B2(new_n651), .ZN(new_n1085));
  OAI21_X1  g660(.A(KEYINPUT41), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT115), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1027), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1082), .B1(new_n1083), .B2(new_n1089), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1020), .B(new_n1081), .C1(new_n1090), .C2(new_n1039), .ZN(new_n1091));
  OAI21_X1  g666(.A(KEYINPUT116), .B1(new_n1091), .B2(KEYINPUT43), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1039), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1079), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1094), .B2(new_n1082), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n1081), .A3(new_n1020), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1096), .A2(KEYINPUT43), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT114), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1092), .A2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1089), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1077), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1101));
  OAI21_X1  g676(.A(new_n1080), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1102), .A2(new_n1093), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n1081), .A2(new_n1020), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT116), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT43), .ZN(new_n1106));
  NAND4_X1  g681(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT114), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1096), .A2(new_n1108), .A3(KEYINPUT43), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1058), .B1(new_n1099), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1091), .A2(KEYINPUT43), .ZN(new_n1112));
  OAI211_X1 g687(.A(new_n1112), .B(KEYINPUT44), .C1(KEYINPUT43), .C2(new_n1096), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(G397));
  AOI21_X1  g689(.A(G1384), .B1(new_n499), .B2(new_n503), .ZN(new_n1115));
  INV_X1    g690(.A(G125), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1116), .B1(new_n490), .B2(new_n491), .ZN(new_n1117));
  INV_X1    g692(.A(new_n471), .ZN(new_n1118));
  OAI21_X1  g693(.A(G2105), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1119), .A2(G40), .A3(new_n465), .A4(new_n466), .ZN(new_n1120));
  NOR3_X1   g695(.A1(new_n1115), .A2(new_n1120), .A3(KEYINPUT45), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1002), .A2(G1996), .A3(new_n1121), .ZN(new_n1122));
  XOR2_X1   g697(.A(new_n1122), .B(KEYINPUT118), .Z(new_n1123));
  NAND2_X1  g698(.A1(new_n822), .A2(G2067), .ZN(new_n1124));
  INV_X1    g699(.A(G2067), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n820), .A2(new_n1125), .A3(new_n821), .ZN(new_n1126));
  AND2_X1   g701(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1123), .B1(new_n1121), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1121), .A2(new_n860), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1130), .A2(new_n1002), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT117), .Z(new_n1132));
  INV_X1    g707(.A(new_n1121), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n886), .B(new_n880), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT119), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1133), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1136), .B1(new_n1135), .B2(new_n1134), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1129), .A2(new_n1132), .A3(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n629), .B(G1986), .Z(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1121), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT122), .B(KEYINPUT57), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1141), .ZN(new_n1142));
  AND2_X1   g717(.A1(new_n598), .A2(new_n599), .ZN(new_n1143));
  INV_X1    g718(.A(new_n590), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n589), .B1(new_n581), .B2(KEYINPUT9), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n582), .A2(new_n585), .ZN(new_n1147));
  OAI22_X1  g722(.A1(new_n1146), .A2(new_n1147), .B1(new_n516), .B2(new_n579), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1142), .B1(new_n1143), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g724(.A(G1956), .ZN(new_n1150));
  INV_X1    g725(.A(G40), .ZN(new_n1151));
  NOR3_X1   g726(.A1(new_n467), .A2(new_n472), .A3(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT50), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1152), .B1(new_n1115), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(G1384), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n493), .A2(G2105), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1156), .B1(new_n463), .B2(new_n464), .ZN(new_n1157));
  AOI22_X1  g732(.A1(new_n1157), .A2(KEYINPUT4), .B1(new_n492), .B2(new_n494), .ZN(new_n1158));
  OAI211_X1 g733(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n1159));
  OR2_X1    g734(.A1(new_n500), .A2(new_n501), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  OAI211_X1 g736(.A(new_n1153), .B(new_n1155), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1162), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1150), .B1(new_n1154), .B2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n592), .A2(new_n600), .A3(new_n1141), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1155), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1166));
  INV_X1    g741(.A(KEYINPUT45), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1120), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  OAI211_X1 g743(.A(KEYINPUT45), .B(new_n1155), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1169));
  XNOR2_X1  g744(.A(KEYINPUT56), .B(G2072), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NAND4_X1  g746(.A1(new_n1149), .A2(new_n1164), .A3(new_n1165), .A4(new_n1171), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1149), .A2(new_n1165), .B1(new_n1164), .B2(new_n1171), .ZN(new_n1173));
  OAI21_X1  g748(.A(new_n867), .B1(new_n1154), .B2(new_n1163), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1115), .A2(new_n1152), .A3(new_n1125), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n652), .B1(new_n1174), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1172), .B1(new_n1173), .B2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1149), .A2(new_n1165), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1164), .A2(new_n1171), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g755(.A1(new_n1180), .A2(KEYINPUT61), .A3(new_n1172), .ZN(new_n1181));
  AND3_X1   g756(.A1(new_n1174), .A2(new_n652), .A3(new_n1175), .ZN(new_n1182));
  OAI21_X1  g757(.A(KEYINPUT60), .B1(new_n1182), .B2(new_n1176), .ZN(new_n1183));
  XOR2_X1   g758(.A(KEYINPUT58), .B(G1341), .Z(new_n1184));
  OAI21_X1  g759(.A(new_n1184), .B1(new_n1166), .B2(new_n1120), .ZN(new_n1185));
  OR2_X1    g760(.A1(new_n1185), .A2(KEYINPUT123), .ZN(new_n1186));
  NAND3_X1  g761(.A1(new_n1168), .A2(new_n860), .A3(new_n1169), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1185), .A2(KEYINPUT123), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1186), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g764(.A(KEYINPUT59), .ZN(new_n1190));
  AND3_X1   g765(.A1(new_n1189), .A2(new_n1190), .A3(new_n573), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1190), .B1(new_n1189), .B2(new_n573), .ZN(new_n1192));
  OAI211_X1 g767(.A(new_n1181), .B(new_n1183), .C1(new_n1191), .C2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n1194));
  AND4_X1   g769(.A1(new_n1165), .A2(new_n1149), .A3(new_n1164), .A4(new_n1171), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1194), .B1(new_n1195), .B2(new_n1173), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT60), .ZN(new_n1197));
  NAND4_X1  g772(.A1(new_n1174), .A2(new_n1197), .A3(new_n654), .A4(new_n1175), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n1177), .B1(new_n1193), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n1201));
  NOR3_X1   g776(.A1(new_n1154), .A2(G2084), .A3(new_n1163), .ZN(new_n1202));
  AOI21_X1  g777(.A(G1966), .B1(new_n1168), .B2(new_n1169), .ZN(new_n1203));
  OAI21_X1  g778(.A(new_n1201), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g779(.A(G1966), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1152), .B1(new_n1115), .B2(KEYINPUT45), .ZN(new_n1206));
  INV_X1    g781(.A(new_n1169), .ZN(new_n1207));
  OAI21_X1  g782(.A(new_n1205), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1120), .B1(new_n1166), .B2(KEYINPUT50), .ZN(new_n1209));
  INV_X1    g784(.A(G2084), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1209), .A2(new_n1210), .A3(new_n1162), .ZN(new_n1211));
  NAND3_X1  g786(.A1(new_n1208), .A2(KEYINPUT124), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g787(.A(G286), .B1(new_n1204), .B2(new_n1212), .ZN(new_n1213));
  INV_X1    g788(.A(KEYINPUT51), .ZN(new_n1214));
  INV_X1    g789(.A(G8), .ZN(new_n1215));
  NOR2_X1   g790(.A1(new_n1214), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1216), .ZN(new_n1217));
  AOI21_X1  g792(.A(new_n1215), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1218));
  OAI21_X1  g793(.A(new_n1214), .B1(G168), .B2(new_n1215), .ZN(new_n1219));
  OAI22_X1  g794(.A1(new_n1213), .A2(new_n1217), .B1(new_n1218), .B2(new_n1219), .ZN(new_n1220));
  NOR2_X1   g795(.A1(G168), .A2(new_n1215), .ZN(new_n1221));
  NAND3_X1  g796(.A1(new_n1204), .A2(new_n1212), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1222), .A2(KEYINPUT125), .ZN(new_n1223));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1204), .A2(new_n1212), .A3(new_n1224), .A4(new_n1221), .ZN(new_n1225));
  NAND3_X1  g800(.A1(new_n1220), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  NOR2_X1   g801(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1227));
  NAND2_X1  g802(.A1(new_n1209), .A2(new_n1162), .ZN(new_n1228));
  OAI22_X1  g803(.A1(new_n1227), .A2(G1971), .B1(new_n1228), .B2(G2090), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1229), .A2(G8), .ZN(new_n1230));
  NAND3_X1  g805(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1231), .ZN(new_n1232));
  AOI21_X1  g807(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1233));
  NOR2_X1   g808(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1230), .A2(new_n1234), .ZN(new_n1235));
  AND2_X1   g810(.A1(new_n604), .A2(G86), .ZN(new_n1236));
  OAI21_X1  g811(.A(G1981), .B1(new_n899), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g812(.A(G1981), .ZN(new_n1238));
  NAND3_X1  g813(.A1(new_n621), .A2(new_n1238), .A3(new_n622), .ZN(new_n1239));
  OR2_X1    g814(.A1(KEYINPUT121), .A2(KEYINPUT49), .ZN(new_n1240));
  NAND2_X1  g815(.A1(KEYINPUT121), .A2(KEYINPUT49), .ZN(new_n1241));
  AOI22_X1  g816(.A1(new_n1237), .A2(new_n1239), .B1(new_n1240), .B2(new_n1241), .ZN(new_n1242));
  AND2_X1   g817(.A1(new_n1237), .A2(new_n1239), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1242), .B1(new_n1243), .B2(new_n1240), .ZN(new_n1244));
  OAI21_X1  g819(.A(G8), .B1(new_n1166), .B2(new_n1120), .ZN(new_n1245));
  NAND2_X1  g820(.A1(new_n1245), .A2(KEYINPUT120), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT120), .ZN(new_n1247));
  OAI211_X1 g822(.A(new_n1247), .B(G8), .C1(new_n1166), .C2(new_n1120), .ZN(new_n1248));
  NAND2_X1  g823(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  INV_X1    g824(.A(G1976), .ZN(new_n1250));
  NOR2_X1   g825(.A1(G288), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g826(.A(new_n1251), .B1(new_n1246), .B2(new_n1248), .ZN(new_n1252));
  AOI21_X1  g827(.A(KEYINPUT52), .B1(G288), .B2(new_n1250), .ZN(new_n1253));
  AOI22_X1  g828(.A1(new_n1244), .A2(new_n1249), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g829(.A(new_n1249), .ZN(new_n1255));
  OAI21_X1  g830(.A(KEYINPUT52), .B1(new_n1255), .B2(new_n1251), .ZN(new_n1256));
  INV_X1    g831(.A(new_n1234), .ZN(new_n1257));
  NAND3_X1  g832(.A1(new_n1229), .A2(G8), .A3(new_n1257), .ZN(new_n1258));
  NAND4_X1  g833(.A1(new_n1235), .A2(new_n1254), .A3(new_n1256), .A4(new_n1258), .ZN(new_n1259));
  INV_X1    g834(.A(new_n1259), .ZN(new_n1260));
  NAND2_X1  g835(.A1(new_n1228), .A2(new_n752), .ZN(new_n1261));
  NAND4_X1  g836(.A1(new_n1168), .A2(KEYINPUT53), .A3(new_n444), .A4(new_n1169), .ZN(new_n1262));
  AND2_X1   g837(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g838(.A(KEYINPUT53), .ZN(new_n1264));
  NAND2_X1  g839(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1265));
  OAI21_X1  g840(.A(new_n1264), .B1(new_n1265), .B2(G2078), .ZN(new_n1266));
  NAND2_X1  g841(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g842(.A1(new_n1267), .A2(G171), .ZN(new_n1268));
  AND4_X1   g843(.A1(G301), .A2(new_n1266), .A3(new_n1261), .A4(new_n1262), .ZN(new_n1269));
  INV_X1    g844(.A(new_n1269), .ZN(new_n1270));
  INV_X1    g845(.A(KEYINPUT54), .ZN(new_n1271));
  NAND3_X1  g846(.A1(new_n1268), .A2(new_n1270), .A3(new_n1271), .ZN(new_n1272));
  AOI21_X1  g847(.A(G301), .B1(new_n1263), .B2(new_n1266), .ZN(new_n1273));
  OAI21_X1  g848(.A(KEYINPUT54), .B1(new_n1273), .B2(new_n1269), .ZN(new_n1274));
  NAND2_X1  g849(.A1(new_n1272), .A2(new_n1274), .ZN(new_n1275));
  NAND4_X1  g850(.A1(new_n1200), .A2(new_n1226), .A3(new_n1260), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g851(.A1(new_n1223), .A2(new_n1225), .ZN(new_n1277));
  NOR2_X1   g852(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1278));
  AND3_X1   g853(.A1(new_n1208), .A2(KEYINPUT124), .A3(new_n1211), .ZN(new_n1279));
  AOI21_X1  g854(.A(KEYINPUT124), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1280));
  OAI21_X1  g855(.A(G168), .B1(new_n1279), .B2(new_n1280), .ZN(new_n1281));
  AOI21_X1  g856(.A(new_n1278), .B1(new_n1281), .B2(new_n1216), .ZN(new_n1282));
  OAI21_X1  g857(.A(KEYINPUT62), .B1(new_n1277), .B2(new_n1282), .ZN(new_n1283));
  INV_X1    g858(.A(KEYINPUT62), .ZN(new_n1284));
  NAND4_X1  g859(.A1(new_n1220), .A2(new_n1284), .A3(new_n1223), .A4(new_n1225), .ZN(new_n1285));
  NOR2_X1   g860(.A1(new_n1259), .A2(new_n1268), .ZN(new_n1286));
  NAND4_X1  g861(.A1(new_n1283), .A2(new_n1285), .A3(KEYINPUT126), .A4(new_n1286), .ZN(new_n1287));
  NAND2_X1  g862(.A1(new_n1254), .A2(new_n1256), .ZN(new_n1288));
  INV_X1    g863(.A(new_n1239), .ZN(new_n1289));
  NAND2_X1  g864(.A1(new_n1244), .A2(new_n1249), .ZN(new_n1290));
  NOR2_X1   g865(.A1(G288), .A2(G1976), .ZN(new_n1291));
  AOI21_X1  g866(.A(new_n1289), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI22_X1  g867(.A1(new_n1288), .A2(new_n1258), .B1(new_n1292), .B2(new_n1255), .ZN(new_n1293));
  INV_X1    g868(.A(KEYINPUT63), .ZN(new_n1294));
  NAND2_X1  g869(.A1(new_n1218), .A2(G168), .ZN(new_n1295));
  OAI21_X1  g870(.A(new_n1294), .B1(new_n1259), .B2(new_n1295), .ZN(new_n1296));
  INV_X1    g871(.A(new_n1288), .ZN(new_n1297));
  AND3_X1   g872(.A1(new_n1229), .A2(G8), .A3(new_n1257), .ZN(new_n1298));
  AOI21_X1  g873(.A(new_n1257), .B1(new_n1229), .B2(G8), .ZN(new_n1299));
  NOR2_X1   g874(.A1(new_n1298), .A2(new_n1299), .ZN(new_n1300));
  INV_X1    g875(.A(new_n1295), .ZN(new_n1301));
  NAND4_X1  g876(.A1(new_n1297), .A2(new_n1300), .A3(KEYINPUT63), .A4(new_n1301), .ZN(new_n1302));
  AOI21_X1  g877(.A(new_n1293), .B1(new_n1296), .B2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g878(.A1(new_n1276), .A2(new_n1287), .A3(new_n1303), .ZN(new_n1304));
  NAND3_X1  g879(.A1(new_n1297), .A2(new_n1300), .A3(new_n1273), .ZN(new_n1305));
  AOI21_X1  g880(.A(new_n1305), .B1(KEYINPUT62), .B2(new_n1226), .ZN(new_n1306));
  AOI21_X1  g881(.A(KEYINPUT126), .B1(new_n1306), .B2(new_n1285), .ZN(new_n1307));
  OAI21_X1  g882(.A(new_n1140), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  AOI21_X1  g883(.A(new_n1133), .B1(new_n1127), .B2(new_n856), .ZN(new_n1309));
  OR2_X1    g884(.A1(new_n1130), .A2(KEYINPUT46), .ZN(new_n1310));
  NAND2_X1  g885(.A1(new_n1130), .A2(KEYINPUT46), .ZN(new_n1311));
  AOI21_X1  g886(.A(new_n1309), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  XOR2_X1   g887(.A(new_n1312), .B(KEYINPUT47), .Z(new_n1313));
  NOR3_X1   g888(.A1(new_n1133), .A2(G1986), .A3(G290), .ZN(new_n1314));
  XOR2_X1   g889(.A(KEYINPUT127), .B(KEYINPUT48), .Z(new_n1315));
  XNOR2_X1  g890(.A(new_n1314), .B(new_n1315), .ZN(new_n1316));
  OAI21_X1  g891(.A(new_n1313), .B1(new_n1138), .B2(new_n1316), .ZN(new_n1317));
  NOR2_X1   g892(.A1(new_n886), .A2(new_n880), .ZN(new_n1318));
  NAND3_X1  g893(.A1(new_n1129), .A2(new_n1132), .A3(new_n1318), .ZN(new_n1319));
  AOI21_X1  g894(.A(new_n1133), .B1(new_n1319), .B2(new_n1126), .ZN(new_n1320));
  NOR2_X1   g895(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g896(.A1(new_n1308), .A2(new_n1321), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g897(.A1(new_n1099), .A2(new_n1110), .ZN(new_n1324));
  OAI21_X1  g898(.A(G319), .B1(new_n700), .B2(new_n701), .ZN(new_n1325));
  NOR2_X1   g899(.A1(new_n1325), .A2(G227), .ZN(new_n1326));
  NAND3_X1  g900(.A1(new_n1022), .A2(new_n746), .A3(new_n1326), .ZN(new_n1327));
  NOR2_X1   g901(.A1(new_n1324), .A2(new_n1327), .ZN(G308));
  AND2_X1   g902(.A1(new_n746), .A2(new_n1326), .ZN(new_n1329));
  OAI211_X1 g903(.A(new_n1329), .B(new_n1022), .C1(new_n1110), .C2(new_n1099), .ZN(G225));
endmodule


