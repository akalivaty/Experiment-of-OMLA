//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 0 1 1 0 0 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 1 0 1 0 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:19 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375, new_n1376;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT64), .Z(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n202), .A2(new_n203), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n213), .A2(G50), .ZN(new_n214));
  INV_X1    g0014(.A(new_n214), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n220));
  INV_X1    g0020(.A(G77), .ZN(new_n221));
  INV_X1    g0021(.A(G244), .ZN(new_n222));
  INV_X1    g0022(.A(G87), .ZN(new_n223));
  INV_X1    g0023(.A(G250), .ZN(new_n224));
  OAI221_X1 g0024(.A(new_n220), .B1(new_n221), .B2(new_n222), .C1(new_n223), .C2(new_n224), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n226));
  INV_X1    g0026(.A(G226), .ZN(new_n227));
  INV_X1    g0027(.A(G97), .ZN(new_n228));
  INV_X1    g0028(.A(G257), .ZN(new_n229));
  OAI221_X1 g0029(.A(new_n226), .B1(new_n201), .B2(new_n227), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n209), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n212), .B(new_n219), .C1(KEYINPUT1), .C2(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n231), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G68), .B(G77), .Z(new_n247));
  XOR2_X1   g0047(.A(G50), .B(G58), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g0049(.A(new_n246), .B(new_n249), .Z(G351));
  INV_X1    g0050(.A(G41), .ZN(new_n251));
  INV_X1    g0051(.A(G45), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT67), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G1), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n253), .A2(new_n255), .A3(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT68), .ZN(new_n259));
  INV_X1    g0059(.A(new_n216), .ZN(new_n260));
  NAND2_X1  g0060(.A1(G33), .A2(G41), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND3_X1   g0062(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n259), .B1(new_n258), .B2(new_n262), .ZN(new_n264));
  OAI21_X1  g0064(.A(KEYINPUT73), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n262), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(KEYINPUT68), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT73), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n258), .A2(new_n259), .A3(new_n262), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n265), .A2(new_n270), .A3(G238), .ZN(new_n271));
  INV_X1    g0071(.A(G274), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n272), .B1(new_n260), .B2(new_n261), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n251), .B2(new_n252), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(KEYINPUT3), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G226), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT72), .B1(new_n281), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  INV_X1    g0085(.A(KEYINPUT72), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n285), .A2(new_n286), .A3(G226), .A4(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(G33), .A2(G97), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(G232), .A3(G1698), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n284), .A2(new_n287), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(new_n262), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n276), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n271), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n293), .A2(KEYINPUT13), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n271), .A2(new_n295), .A3(new_n292), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT77), .ZN(new_n300));
  AND3_X1   g0100(.A1(new_n271), .A2(new_n295), .A3(new_n292), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n295), .B1(new_n271), .B2(new_n292), .ZN(new_n302));
  OAI21_X1  g0102(.A(G169), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n300), .B1(new_n303), .B2(KEYINPUT14), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT14), .ZN(new_n305));
  NAND4_X1  g0105(.A1(new_n297), .A2(KEYINPUT77), .A3(new_n305), .A4(G169), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n299), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(G169), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n294), .B2(new_n296), .ZN(new_n309));
  OAI21_X1  g0109(.A(KEYINPUT76), .B1(new_n309), .B2(new_n305), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT76), .ZN(new_n311));
  NAND3_X1  g0111(.A1(new_n303), .A2(new_n311), .A3(KEYINPUT14), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND4_X1  g0114(.A1(new_n255), .A2(new_n257), .A3(G13), .A4(G20), .ZN(new_n315));
  NAND3_X1  g0115(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n216), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n315), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT67), .B(G1), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G20), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT70), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n315), .A2(new_n318), .A3(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n320), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(G68), .ZN(new_n326));
  INV_X1    g0126(.A(new_n315), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n203), .ZN(new_n328));
  XNOR2_X1  g0128(.A(new_n328), .B(KEYINPUT12), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(KEYINPUT75), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G20), .A2(G33), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G50), .ZN(new_n334));
  XOR2_X1   g0134(.A(new_n334), .B(KEYINPUT74), .Z(new_n335));
  NOR2_X1   g0135(.A1(new_n277), .A2(G20), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(G77), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n217), .B2(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n317), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n339), .B(KEYINPUT11), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n331), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n314), .A2(new_n341), .ZN(new_n342));
  AND3_X1   g0142(.A1(new_n331), .A2(new_n332), .A3(new_n340), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n294), .A2(G190), .A3(new_n296), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n297), .A2(G200), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n342), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT81), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT79), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n349), .B1(new_n277), .B2(KEYINPUT3), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n279), .A2(KEYINPUT79), .A3(G33), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT78), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n353), .B1(new_n279), .B2(G33), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n277), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(G223), .A2(G1698), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n227), .B2(G1698), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n352), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(G33), .A2(G87), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n291), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n258), .A2(G232), .A3(new_n262), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(new_n275), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n308), .B1(new_n362), .B2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n262), .B1(new_n359), .B2(new_n360), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n367), .A2(new_n364), .A3(new_n298), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n348), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  AOI22_X1  g0169(.A1(new_n350), .A2(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n370));
  AOI22_X1  g0170(.A1(new_n370), .A2(new_n358), .B1(G33), .B2(G87), .ZN(new_n371));
  OAI211_X1 g0171(.A(new_n365), .B(G179), .C1(new_n371), .C2(new_n262), .ZN(new_n372));
  OAI21_X1  g0172(.A(G169), .B1(new_n367), .B2(new_n364), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n372), .A2(new_n373), .A3(KEYINPUT81), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(G58), .A2(G68), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n213), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(G20), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT80), .ZN(new_n379));
  INV_X1    g0179(.A(G159), .ZN(new_n380));
  INV_X1    g0180(.A(new_n333), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n380), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n217), .B1(new_n213), .B2(new_n376), .ZN(new_n384));
  OAI21_X1  g0184(.A(KEYINPUT80), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(G20), .B1(new_n352), .B2(new_n356), .ZN(new_n387));
  INV_X1    g0187(.A(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n370), .A2(KEYINPUT7), .A3(G20), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n386), .B(KEYINPUT16), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT16), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n388), .B1(new_n285), .B2(G20), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n281), .A2(KEYINPUT7), .A3(new_n217), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n203), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n392), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n391), .A2(new_n317), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n322), .A2(new_n318), .ZN(new_n399));
  NOR3_X1   g0199(.A1(new_n202), .A2(KEYINPUT69), .A3(KEYINPUT8), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT8), .B(G58), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n400), .B1(new_n401), .B2(KEYINPUT69), .ZN(new_n402));
  MUX2_X1   g0202(.A(new_n315), .B(new_n399), .S(new_n402), .Z(new_n403));
  NAND2_X1  g0203(.A1(new_n398), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n375), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n375), .A2(new_n404), .A3(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(KEYINPUT82), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g0209(.A(KEYINPUT18), .B1(new_n375), .B2(new_n404), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT82), .ZN(new_n411));
  INV_X1    g0211(.A(G200), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(new_n362), .B2(new_n365), .ZN(new_n413));
  INV_X1    g0213(.A(G190), .ZN(new_n414));
  NOR3_X1   g0214(.A1(new_n367), .A2(new_n414), .A3(new_n364), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n398), .A2(new_n416), .A3(new_n403), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT17), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT17), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n398), .A2(new_n416), .A3(new_n419), .A4(new_n403), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n410), .A2(new_n411), .B1(new_n418), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n409), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n267), .A2(new_n269), .ZN(new_n423));
  XOR2_X1   g0223(.A(KEYINPUT66), .B(G226), .Z(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n282), .A2(G222), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G223), .A2(G1698), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n285), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n262), .B1(new_n281), .B2(new_n221), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n276), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n431), .A2(new_n414), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(G200), .B2(new_n431), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n402), .A2(new_n336), .ZN(new_n434));
  AOI22_X1  g0234(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n333), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n318), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n327), .A2(new_n201), .ZN(new_n437));
  OAI21_X1  g0237(.A(new_n437), .B1(new_n399), .B2(new_n201), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g0239(.A(new_n439), .B(KEYINPUT9), .Z(new_n440));
  INV_X1    g0240(.A(KEYINPUT10), .ZN(new_n441));
  AND3_X1   g0241(.A1(new_n433), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n433), .B2(new_n440), .ZN(new_n443));
  OR2_X1    g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n431), .A2(new_n308), .ZN(new_n445));
  INV_X1    g0245(.A(new_n439), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n425), .A2(new_n430), .A3(new_n298), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n445), .A2(new_n446), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT71), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n423), .A2(G244), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G238), .A2(G1698), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n285), .B(new_n452), .C1(new_n237), .C2(G1698), .ZN(new_n453));
  INV_X1    g0253(.A(G107), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n262), .B1(new_n281), .B2(new_n454), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n276), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n451), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G200), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n325), .A2(G77), .ZN(new_n460));
  XNOR2_X1  g0260(.A(KEYINPUT15), .B(G87), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI22_X1  g0262(.A1(new_n462), .A2(new_n336), .B1(G20), .B2(G77), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n463), .B1(new_n381), .B2(new_n401), .ZN(new_n464));
  AOI22_X1  g0264(.A1(new_n464), .A2(new_n317), .B1(new_n221), .B2(new_n327), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n460), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n450), .B1(new_n459), .B2(new_n466), .ZN(new_n467));
  NAND4_X1  g0267(.A1(new_n458), .A2(KEYINPUT71), .A3(new_n460), .A4(new_n465), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n467), .B(new_n468), .C1(new_n414), .C2(new_n457), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n457), .A2(new_n308), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n451), .A2(new_n456), .A3(new_n298), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n466), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n469), .A2(new_n472), .ZN(new_n473));
  NOR4_X1   g0273(.A1(new_n347), .A2(new_n422), .A3(new_n449), .A4(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(G33), .A2(G283), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n282), .A2(KEYINPUT4), .A3(G244), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n285), .A2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT4), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n479), .B1(new_n285), .B2(G250), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n475), .B(new_n478), .C1(new_n480), .C2(new_n282), .ZN(new_n481));
  AOI21_X1  g0281(.A(KEYINPUT4), .B1(new_n370), .B2(G244), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n291), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT5), .B(G41), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n255), .A2(new_n257), .A3(G45), .ZN(new_n486));
  OAI211_X1 g0286(.A(G257), .B(new_n262), .C1(new_n485), .C2(new_n486), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n273), .A2(G45), .A3(new_n321), .A4(new_n484), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n483), .A2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  NOR3_X1   g0292(.A1(new_n492), .A2(new_n228), .A3(G107), .ZN(new_n493));
  XNOR2_X1  g0293(.A(G97), .B(G107), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n493), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n495), .A2(new_n217), .B1(new_n221), .B2(new_n381), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n454), .B1(new_n393), .B2(new_n394), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n317), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n315), .A2(G97), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n319), .B1(G33), .B2(new_n321), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G97), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n491), .A2(new_n308), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT83), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n278), .A2(new_n280), .A3(G250), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n282), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n475), .B1(new_n281), .B2(new_n476), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n352), .A2(new_n356), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n479), .B1(new_n508), .B2(new_n222), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n489), .B1(new_n510), .B2(new_n291), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n503), .B1(new_n511), .B2(new_n298), .ZN(new_n512));
  AND4_X1   g0312(.A1(new_n503), .A2(new_n483), .A3(new_n298), .A4(new_n490), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n502), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT84), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(KEYINPUT85), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n502), .B(KEYINPUT84), .C1(new_n512), .C2(new_n513), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n511), .A2(G190), .ZN(new_n519));
  AND2_X1   g0319(.A1(new_n501), .A2(new_n498), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n519), .B(new_n520), .C1(new_n412), .C2(new_n511), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n516), .A2(new_n517), .A3(new_n518), .A4(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(KEYINPUT85), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n255), .A2(new_n257), .A3(G33), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n525), .A2(G116), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n320), .A2(new_n324), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n315), .A2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n316), .A2(new_n216), .B1(G20), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n475), .B(new_n217), .C1(G33), .C2(new_n228), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n528), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G303), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n285), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n229), .A2(G1698), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n540), .B1(new_n370), .B2(new_n541), .ZN(new_n542));
  AND2_X1   g0342(.A1(G264), .A2(G1698), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n352), .A2(new_n356), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT87), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n370), .A2(KEYINPUT87), .A3(new_n543), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n291), .ZN(new_n549));
  OAI211_X1 g0349(.A(G270), .B(new_n262), .C1(new_n485), .C2(new_n486), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n488), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n538), .B1(new_n553), .B2(G200), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n551), .B1(new_n548), .B2(new_n291), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(G190), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT24), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n217), .A2(G87), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT22), .B1(new_n285), .B2(new_n560), .ZN(new_n561));
  AND3_X1   g0361(.A1(new_n454), .A2(KEYINPUT23), .A3(G20), .ZN(new_n562));
  AOI21_X1  g0362(.A(KEYINPUT23), .B1(new_n454), .B2(G20), .ZN(new_n563));
  NAND2_X1  g0363(.A1(G33), .A2(G116), .ZN(new_n564));
  OAI22_X1  g0364(.A1(new_n562), .A2(new_n563), .B1(G20), .B2(new_n564), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n561), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n559), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n352), .A2(new_n356), .A3(new_n568), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n558), .B1(new_n566), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n567), .B1(new_n281), .B2(new_n559), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n564), .A2(G20), .ZN(new_n572));
  INV_X1    g0372(.A(new_n563), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n454), .A2(KEYINPUT23), .A3(G20), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n572), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n558), .A2(new_n569), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n317), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  OR3_X1    g0377(.A1(new_n315), .A2(KEYINPUT25), .A3(G107), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n315), .A2(new_n318), .A3(new_n525), .A4(G107), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT25), .B1(new_n315), .B2(G107), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(G264), .B(new_n262), .C1(new_n485), .C2(new_n486), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(new_n488), .ZN(new_n584));
  INV_X1    g0384(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g0385(.A1(G250), .A2(G1698), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n586), .B1(new_n229), .B2(G1698), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n352), .A2(new_n356), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(G33), .A2(G294), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n262), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n585), .A2(new_n591), .A3(G190), .ZN(new_n592));
  OAI21_X1  g0392(.A(G200), .B1(new_n584), .B2(new_n590), .ZN(new_n593));
  NAND4_X1  g0393(.A1(new_n577), .A2(new_n582), .A3(new_n592), .A4(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n557), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g0395(.A1(new_n584), .A2(new_n590), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n298), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n569), .A2(new_n575), .A3(new_n571), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(KEYINPUT24), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n566), .A2(new_n558), .A3(new_n569), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n318), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI221_X1 g0401(.A(new_n597), .B1(G169), .B2(new_n596), .C1(new_n601), .C2(new_n581), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n298), .B1(new_n528), .B2(new_n537), .ZN(new_n603));
  AND3_X1   g0403(.A1(new_n603), .A2(new_n549), .A3(new_n552), .ZN(new_n604));
  INV_X1    g0404(.A(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT21), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n308), .B1(new_n528), .B2(new_n537), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n606), .B1(new_n553), .B2(new_n607), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n315), .A2(new_n323), .A3(new_n318), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n323), .B1(new_n315), .B2(new_n318), .ZN(new_n610));
  NOR3_X1   g0410(.A1(new_n609), .A2(new_n610), .A3(new_n526), .ZN(new_n611));
  AND3_X1   g0411(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n532), .ZN(new_n612));
  AOI21_X1  g0412(.A(KEYINPUT20), .B1(new_n531), .B2(new_n532), .ZN(new_n613));
  OAI22_X1  g0413(.A1(new_n612), .A2(new_n613), .B1(G116), .B2(new_n315), .ZN(new_n614));
  OAI21_X1  g0414(.A(G169), .B1(new_n611), .B2(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n555), .A2(new_n615), .A3(KEYINPUT21), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n602), .B(new_n605), .C1(new_n608), .C2(new_n616), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n462), .A2(new_n315), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n462), .A2(new_n315), .A3(new_n318), .A4(new_n525), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n352), .A2(new_n356), .A3(new_n217), .A4(G68), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT19), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n622), .B1(new_n288), .B2(new_n217), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n223), .A2(new_n228), .A3(new_n454), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n217), .A2(G33), .A3(G97), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n623), .A2(new_n624), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n621), .A2(new_n626), .ZN(new_n627));
  OAI211_X1 g0427(.A(new_n619), .B(new_n620), .C1(new_n627), .C2(new_n318), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n486), .A2(new_n224), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n321), .A2(G45), .A3(new_n272), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n262), .ZN(new_n631));
  NOR2_X1   g0431(.A1(G238), .A2(G1698), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n632), .B1(new_n222), .B2(G1698), .ZN(new_n633));
  AOI22_X1  g0433(.A1(new_n370), .A2(new_n633), .B1(G33), .B2(G116), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n298), .B(new_n631), .C1(new_n634), .C2(new_n262), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n352), .A2(new_n356), .A3(new_n633), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n262), .B1(new_n636), .B2(new_n564), .ZN(new_n637));
  AND3_X1   g0437(.A1(new_n629), .A2(new_n630), .A3(new_n262), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n308), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n628), .A2(new_n635), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n318), .B1(new_n621), .B2(new_n626), .ZN(new_n641));
  AND4_X1   g0441(.A1(G87), .A2(new_n315), .A3(new_n318), .A4(new_n525), .ZN(new_n642));
  NOR3_X1   g0442(.A1(new_n641), .A2(new_n618), .A3(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(G200), .B1(new_n637), .B2(new_n638), .ZN(new_n644));
  OAI211_X1 g0444(.A(G190), .B(new_n631), .C1(new_n634), .C2(new_n262), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT86), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n640), .A2(new_n646), .A3(KEYINPUT86), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n595), .A2(new_n617), .A3(new_n651), .ZN(new_n652));
  AND4_X1   g0452(.A1(new_n474), .A2(new_n522), .A3(new_n524), .A4(new_n652), .ZN(G372));
  INV_X1    g0453(.A(new_n448), .ZN(new_n654));
  INV_X1    g0454(.A(new_n472), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n346), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n342), .A2(new_n656), .A3(KEYINPUT89), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT89), .ZN(new_n658));
  INV_X1    g0458(.A(new_n656), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n343), .B1(new_n307), .B2(new_n313), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n418), .A2(new_n420), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n657), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n372), .A2(new_n373), .ZN(new_n664));
  AND3_X1   g0464(.A1(new_n404), .A2(new_n406), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n406), .B1(new_n404), .B2(new_n664), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n654), .B1(new_n668), .B2(new_n444), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n644), .A2(KEYINPUT88), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT88), .ZN(new_n671));
  OAI211_X1 g0471(.A(new_n671), .B(G200), .C1(new_n637), .C2(new_n638), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n670), .A2(new_n645), .A3(new_n643), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n673), .A2(new_n640), .ZN(new_n674));
  OR3_X1    g0474(.A1(new_n514), .A2(new_n674), .A3(KEYINPUT26), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n651), .B1(new_n516), .B2(new_n518), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT26), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n673), .A2(new_n594), .A3(new_n640), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n617), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n640), .B1(new_n523), .B2(new_n681), .ZN(new_n682));
  OR2_X1    g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n474), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n669), .A2(new_n684), .ZN(G369));
  INV_X1    g0485(.A(new_n602), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n217), .A2(G13), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n321), .A2(new_n687), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n601), .A2(new_n581), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n594), .B1(new_n696), .B2(new_n694), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(new_n602), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n553), .A2(new_n606), .A3(new_n607), .ZN(new_n701));
  OAI21_X1  g0501(.A(KEYINPUT21), .B1(new_n555), .B2(new_n615), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n604), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n693), .A2(new_n538), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n703), .A2(new_n704), .ZN(new_n706));
  OAI211_X1 g0506(.A(G330), .B(new_n557), .C1(new_n705), .C2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT90), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n708), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n700), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n703), .A2(new_n693), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n700), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n713), .A2(new_n695), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n711), .A2(new_n715), .ZN(G399));
  INV_X1    g0516(.A(new_n650), .ZN(new_n717));
  AOI21_X1  g0517(.A(KEYINPUT86), .B1(new_n640), .B2(new_n646), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n518), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n483), .A2(new_n298), .A3(new_n490), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(KEYINPUT83), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n511), .A2(new_n503), .A3(new_n298), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(KEYINPUT84), .B1(new_n724), .B2(new_n502), .ZN(new_n725));
  OAI211_X1 g0525(.A(new_n719), .B(new_n677), .C1(new_n720), .C2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT26), .B1(new_n514), .B2(new_n674), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n694), .B1(new_n728), .B2(new_n682), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n729), .A2(KEYINPUT91), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT91), .ZN(new_n731));
  OAI211_X1 g0531(.A(new_n731), .B(new_n694), .C1(new_n728), .C2(new_n682), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT29), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n683), .A2(new_n694), .ZN(new_n735));
  INV_X1    g0535(.A(KEYINPUT29), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT92), .ZN(new_n739));
  INV_X1    g0539(.A(G330), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n524), .A2(new_n652), .A3(new_n522), .A4(new_n694), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n511), .A2(new_n549), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n637), .A2(new_n638), .ZN(new_n743));
  NAND4_X1  g0543(.A1(new_n596), .A2(new_n743), .A3(G179), .A4(new_n550), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n742), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n596), .A2(new_n743), .A3(G179), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n747), .A2(new_n491), .A3(new_n553), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n745), .B1(new_n742), .B2(new_n744), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n746), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  AND3_X1   g0550(.A1(new_n750), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n751));
  AOI21_X1  g0551(.A(KEYINPUT31), .B1(new_n750), .B2(new_n693), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n740), .B1(new_n741), .B2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n738), .A2(new_n739), .A3(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g0557(.A(new_n739), .B1(new_n738), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n254), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n624), .A2(G116), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n210), .A2(new_n251), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n761), .A2(new_n762), .A3(G1), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(new_n214), .B2(new_n762), .ZN(new_n764));
  XNOR2_X1  g0564(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n760), .A2(new_n765), .ZN(G364));
  NOR2_X1   g0566(.A1(new_n705), .A2(new_n706), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n556), .B2(new_n554), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(G13), .A2(G33), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(G20), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n216), .B1(G20), .B2(new_n308), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n217), .A2(G179), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G190), .A2(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n777), .A2(new_n380), .ZN(new_n778));
  XNOR2_X1  g0578(.A(new_n778), .B(KEYINPUT32), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n217), .A2(new_n298), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n780), .A2(G190), .A3(new_n412), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n281), .B1(new_n782), .B2(G58), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n780), .A2(new_n776), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n779), .B(new_n783), .C1(new_n221), .C2(new_n784), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n775), .A2(new_n414), .A3(G200), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n786), .B(KEYINPUT94), .Z(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n788), .A2(new_n454), .ZN(new_n789));
  NOR3_X1   g0589(.A1(new_n414), .A2(G179), .A3(G200), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n217), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n775), .A2(G190), .A3(G200), .ZN(new_n792));
  OAI22_X1  g0592(.A1(new_n791), .A2(new_n228), .B1(new_n792), .B2(new_n223), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n780), .A2(G200), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(G190), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n794), .A2(new_n414), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n796), .A2(new_n203), .B1(new_n798), .B2(new_n201), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n785), .A2(new_n789), .A3(new_n793), .A4(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G322), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n781), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G311), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n281), .B1(new_n784), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(new_n777), .ZN(new_n805));
  AOI211_X1 g0605(.A(new_n802), .B(new_n804), .C1(G329), .C2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(new_n791), .ZN(new_n807));
  INV_X1    g0607(.A(new_n792), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n807), .A2(G294), .B1(new_n808), .B2(G303), .ZN(new_n809));
  XNOR2_X1  g0609(.A(KEYINPUT95), .B(G326), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  XNOR2_X1  g0611(.A(KEYINPUT33), .B(G317), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n797), .A2(new_n811), .B1(new_n795), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n806), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(G283), .B2(new_n787), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n774), .B1(new_n800), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n687), .A2(G45), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n762), .A2(new_n817), .A3(G1), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n772), .A2(new_n774), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n508), .A2(new_n210), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n249), .A2(G45), .ZN(new_n822));
  XNOR2_X1  g0622(.A(new_n822), .B(KEYINPUT93), .ZN(new_n823));
  AOI211_X1 g0623(.A(new_n821), .B(new_n823), .C1(new_n252), .C2(new_n215), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n285), .A2(new_n210), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n207), .A2(new_n825), .B1(G116), .B2(new_n210), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n820), .B1(new_n824), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n773), .A2(new_n816), .A3(new_n819), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n709), .A2(new_n710), .ZN(new_n829));
  OAI211_X1 g0629(.A(new_n829), .B(new_n818), .C1(G330), .C2(new_n768), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n828), .A2(new_n830), .ZN(G396));
  NAND2_X1  g0631(.A1(new_n466), .A2(new_n693), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n469), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(new_n472), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n472), .A2(new_n693), .ZN(new_n835));
  INV_X1    g0635(.A(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n735), .A2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n835), .B1(new_n833), .B2(new_n472), .ZN(new_n839));
  OAI211_X1 g0639(.A(new_n839), .B(new_n694), .C1(new_n678), .C2(new_n682), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n819), .B1(new_n841), .B2(new_n755), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n842), .B1(new_n755), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n774), .A2(new_n770), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n818), .B1(new_n221), .B2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n774), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n788), .A2(new_n223), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n807), .A2(G97), .B1(new_n808), .B2(G107), .ZN(new_n848));
  INV_X1    g0648(.A(G283), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n796), .C1(new_n539), .C2(new_n798), .ZN(new_n850));
  INV_X1    g0650(.A(new_n784), .ZN(new_n851));
  AOI22_X1  g0651(.A1(G116), .A2(new_n851), .B1(new_n805), .B2(G311), .ZN(new_n852));
  INV_X1    g0652(.A(G294), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n852), .B(new_n281), .C1(new_n853), .C2(new_n781), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n847), .A2(new_n850), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(new_n782), .A2(G143), .B1(new_n851), .B2(G159), .ZN(new_n856));
  INV_X1    g0656(.A(G137), .ZN(new_n857));
  INV_X1    g0657(.A(G150), .ZN(new_n858));
  OAI221_X1 g0658(.A(new_n856), .B1(new_n798), .B2(new_n857), .C1(new_n858), .C2(new_n796), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT34), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n788), .A2(new_n203), .ZN(new_n862));
  INV_X1    g0662(.A(G132), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n370), .B1(new_n863), .B2(new_n777), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n791), .A2(new_n202), .B1(new_n792), .B2(new_n201), .ZN(new_n865));
  NOR4_X1   g0665(.A1(new_n861), .A2(new_n862), .A3(new_n864), .A4(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n859), .A2(new_n860), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n855), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  OAI221_X1 g0668(.A(new_n845), .B1(new_n846), .B2(new_n868), .C1(new_n839), .C2(new_n771), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n843), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(G384));
  INV_X1    g0671(.A(new_n495), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n872), .A2(KEYINPUT35), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n872), .A2(KEYINPUT35), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n873), .A2(G116), .A3(new_n218), .A4(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT36), .Z(new_n876));
  NAND2_X1  g0676(.A1(new_n376), .A2(G77), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n214), .A2(new_n877), .B1(G50), .B2(new_n203), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n321), .A2(G13), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n691), .B1(new_n665), .B2(new_n666), .ZN(new_n881));
  INV_X1    g0681(.A(KEYINPUT38), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n391), .A2(new_n317), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n387), .A2(new_n388), .ZN(new_n884));
  OAI21_X1  g0684(.A(KEYINPUT7), .B1(new_n370), .B2(G20), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n884), .A2(new_n885), .A3(G68), .ZN(new_n886));
  AOI21_X1  g0686(.A(KEYINPUT16), .B1(new_n886), .B2(new_n386), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n403), .B1(new_n883), .B2(new_n887), .ZN(new_n888));
  INV_X1    g0688(.A(new_n691), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n409), .B2(new_n421), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n888), .A2(new_n664), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n892), .A2(new_n890), .A3(new_n417), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n404), .A2(new_n889), .ZN(new_n894));
  AND2_X1   g0694(.A1(new_n894), .A2(new_n417), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT37), .B1(new_n375), .B2(new_n404), .ZN(new_n896));
  AOI22_X1  g0696(.A1(KEYINPUT37), .A2(new_n893), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n882), .B1(new_n891), .B2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n890), .ZN(new_n899));
  AND3_X1   g0699(.A1(new_n375), .A2(KEYINPUT18), .A3(new_n404), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n900), .A2(new_n410), .A3(new_n411), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n405), .A2(new_n411), .A3(new_n406), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n662), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n899), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n895), .A2(new_n896), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(KEYINPUT38), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n341), .A2(new_n693), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g0712(.A(KEYINPUT97), .B1(new_n314), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT97), .ZN(new_n914));
  AOI211_X1 g0714(.A(new_n914), .B(new_n911), .C1(new_n307), .C2(new_n313), .ZN(new_n915));
  OAI22_X1  g0715(.A1(new_n347), .A2(new_n912), .B1(new_n913), .B2(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n835), .B(KEYINPUT96), .Z(new_n917));
  NAND2_X1  g0717(.A1(new_n840), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT39), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n894), .B1(new_n667), .B2(new_n662), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n404), .A2(new_n664), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(new_n894), .A3(new_n417), .ZN(new_n923));
  AOI22_X1  g0723(.A1(new_n895), .A2(new_n896), .B1(new_n923), .B2(KEYINPUT37), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n882), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n908), .A2(new_n920), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n926), .A2(KEYINPUT99), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n909), .A2(KEYINPUT39), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT99), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n908), .A2(new_n925), .A3(new_n929), .A4(new_n920), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n928), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n931), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n314), .A2(new_n341), .A3(new_n694), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT98), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n660), .A2(KEYINPUT98), .A3(new_n694), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  OAI221_X1 g0738(.A(new_n881), .B1(new_n910), .B2(new_n919), .C1(new_n932), .C2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n734), .A2(new_n474), .A3(new_n737), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n669), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n939), .B(new_n941), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n837), .B1(new_n741), .B2(new_n753), .ZN(new_n943));
  AND2_X1   g0743(.A1(new_n916), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n945), .B1(new_n908), .B2(new_n925), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n913), .A2(new_n915), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n660), .A2(new_n948), .A3(new_n912), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n909), .B(new_n943), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n944), .A2(new_n946), .B1(new_n950), .B2(new_n945), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n741), .A2(new_n753), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n474), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(G330), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n955), .B1(new_n954), .B2(new_n952), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n942), .A2(new_n956), .B1(new_n321), .B2(new_n687), .ZN(new_n957));
  AND2_X1   g0757(.A1(new_n942), .A2(new_n956), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n880), .B1(new_n957), .B2(new_n958), .ZN(G367));
  NOR2_X1   g0759(.A1(new_n694), .A2(new_n643), .ZN(new_n960));
  MUX2_X1   g0760(.A(new_n674), .B(new_n640), .S(new_n960), .Z(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT100), .Z(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(new_n772), .ZN(new_n963));
  INV_X1    g0763(.A(new_n241), .ZN(new_n964));
  OAI221_X1 g0764(.A(new_n820), .B1(new_n210), .B2(new_n461), .C1(new_n964), .C2(new_n821), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n965), .A2(new_n819), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n796), .A2(new_n853), .B1(new_n454), .B2(new_n791), .ZN(new_n967));
  INV_X1    g0767(.A(new_n786), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n967), .B1(G97), .B2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(G317), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n781), .A2(new_n539), .B1(new_n777), .B2(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G283), .B2(new_n851), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n370), .B1(new_n797), .B2(G311), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n808), .A2(G116), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n969), .A2(new_n972), .A3(new_n973), .A4(new_n975), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n781), .A2(new_n858), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n791), .A2(new_n203), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n977), .B(new_n978), .C1(G143), .C2(new_n797), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT106), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n784), .A2(new_n201), .B1(new_n777), .B2(new_n857), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G159), .B2(new_n795), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n285), .B1(new_n786), .B2(new_n221), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT107), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n808), .A2(G58), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n982), .A2(new_n985), .A3(new_n986), .A4(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n976), .B1(new_n980), .B2(new_n988), .ZN(new_n989));
  XNOR2_X1  g0789(.A(new_n989), .B(KEYINPUT47), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n966), .B1(new_n990), .B2(new_n774), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n963), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n516), .A2(new_n518), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n724), .A2(new_n502), .A3(new_n693), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(KEYINPUT101), .Z(new_n996));
  OR2_X1    g0796(.A1(new_n520), .A2(new_n694), .ZN(new_n997));
  NAND4_X1  g0797(.A1(new_n516), .A2(new_n518), .A3(new_n521), .A4(new_n997), .ZN(new_n998));
  AND2_X1   g0798(.A1(new_n996), .A2(new_n998), .ZN(new_n999));
  OAI211_X1 g0799(.A(KEYINPUT102), .B(new_n994), .C1(new_n999), .C2(new_n602), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT102), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n602), .B1(new_n996), .B2(new_n998), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1001), .B1(new_n1002), .B2(new_n993), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n694), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT42), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1005), .B1(new_n999), .B2(new_n713), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n996), .A2(new_n998), .ZN(new_n1007));
  NAND4_X1  g0807(.A1(new_n1007), .A2(KEYINPUT42), .A3(new_n700), .A4(new_n712), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1004), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT103), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT43), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n962), .B1(new_n1004), .B2(new_n1009), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1010), .A2(KEYINPUT103), .A3(KEYINPUT43), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n962), .ZN(new_n1018));
  AOI21_X1  g0818(.A(KEYINPUT43), .B1(new_n1010), .B2(KEYINPUT103), .ZN(new_n1019));
  INV_X1    g0819(.A(KEYINPUT103), .ZN(new_n1020));
  AOI211_X1 g0820(.A(new_n1020), .B(new_n1012), .C1(new_n1004), .C2(new_n1009), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1018), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n711), .A2(new_n999), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n1024), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1017), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n817), .A2(G1), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n1030));
  OR3_X1    g0830(.A1(new_n999), .A2(new_n714), .A3(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n1030), .B1(new_n999), .B2(new_n714), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT105), .B(KEYINPUT44), .Z(new_n1033));
  NAND3_X1  g0833(.A1(new_n999), .A2(new_n714), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1033), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n715), .B2(new_n1007), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .A4(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n711), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1037), .B(new_n1038), .ZN(new_n1039));
  NOR3_X1   g0839(.A1(new_n709), .A2(new_n710), .A3(new_n700), .ZN(new_n1040));
  INV_X1    g0840(.A(new_n1040), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1041), .A2(new_n711), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n712), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1039), .A2(new_n1044), .B1(new_n757), .B2(new_n758), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n762), .B(KEYINPUT41), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n1046), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1029), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n992), .B1(new_n1028), .B2(new_n1048), .ZN(G387));
  NAND2_X1  g0849(.A1(new_n238), .A2(G45), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT109), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n401), .A2(G50), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n761), .ZN(new_n1054));
  AOI211_X1 g0854(.A(G45), .B(new_n1054), .C1(G68), .C2(G77), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n821), .B(new_n1051), .C1(new_n1053), .C2(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n825), .A2(new_n761), .B1(G107), .B2(new_n210), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n820), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G68), .A2(new_n851), .B1(new_n805), .B2(G150), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n201), .B2(new_n781), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1060), .B1(new_n402), .B2(new_n795), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n791), .A2(new_n461), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n370), .B1(new_n221), .B2(new_n792), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G159), .C2(new_n797), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n1061), .B(new_n1064), .C1(new_n228), .C2(new_n788), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n370), .B1(new_n805), .B2(new_n811), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n791), .A2(new_n849), .B1(new_n792), .B2(new_n853), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n782), .A2(G317), .B1(new_n851), .B2(G303), .ZN(new_n1068));
  OAI221_X1 g0868(.A(new_n1068), .B1(new_n798), .B2(new_n801), .C1(new_n803), .C2(new_n796), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT48), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1067), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1071), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1066), .B1(new_n530), .B2(new_n786), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1065), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n818), .B1(new_n1076), .B2(new_n774), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1058), .A2(new_n1077), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n699), .B2(new_n772), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1029), .ZN(new_n1080));
  OR3_X1    g0880(.A1(new_n1044), .A2(KEYINPUT108), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g0881(.A(KEYINPUT108), .B1(new_n1044), .B2(new_n1080), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1079), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n738), .A2(new_n755), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT92), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1085), .A2(new_n1044), .A3(KEYINPUT110), .A4(new_n756), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n762), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n1087), .C1(new_n759), .C2(new_n1044), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT110), .B1(new_n759), .B2(new_n1044), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1083), .B1(new_n1088), .B2(new_n1089), .ZN(G393));
  INV_X1    g0890(.A(new_n1039), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n1029), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n798), .A2(new_n858), .B1(new_n380), .B2(new_n781), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT51), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n847), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n784), .A2(new_n401), .ZN(new_n1096));
  AOI211_X1 g0896(.A(new_n508), .B(new_n1096), .C1(G143), .C2(new_n805), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n796), .A2(new_n201), .B1(new_n792), .B2(new_n203), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n1098), .B1(G77), .B2(new_n807), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1094), .A2(new_n1095), .A3(new_n1097), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n281), .B1(new_n777), .B2(new_n801), .ZN(new_n1101));
  AOI211_X1 g0901(.A(new_n1101), .B(new_n789), .C1(G283), .C2(new_n808), .ZN(new_n1102));
  XNOR2_X1  g0902(.A(new_n1102), .B(KEYINPUT112), .ZN(new_n1103));
  AOI22_X1  g0903(.A1(new_n795), .A2(G303), .B1(new_n851), .B2(G294), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1103), .B(new_n1104), .C1(new_n530), .C2(new_n791), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n798), .A2(new_n970), .B1(new_n803), .B2(new_n781), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(new_n1106), .B(KEYINPUT111), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT52), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1100), .B1(new_n1105), .B2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1109), .A2(new_n774), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n999), .A2(new_n772), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n820), .B1(new_n228), .B2(new_n210), .C1(new_n246), .C2(new_n821), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n819), .A4(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1092), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1044), .B1(new_n1085), .B2(new_n756), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n762), .B1(new_n1115), .B2(new_n1091), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1039), .B1(new_n759), .B2(new_n1044), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1114), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(G390));
  OAI211_X1 g0919(.A(new_n754), .B(new_n839), .C1(new_n947), .C2(new_n949), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n908), .A2(new_n925), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n938), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n732), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n679), .B1(new_n703), .B2(new_n602), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1125), .A2(new_n516), .A3(new_n518), .A4(new_n521), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1126), .A2(new_n640), .A3(new_n727), .A4(new_n726), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n731), .B1(new_n1127), .B2(new_n694), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n839), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1129), .A2(new_n917), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1123), .B1(new_n1130), .B2(new_n916), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n937), .B1(new_n916), .B2(new_n918), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n931), .A2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1121), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n937), .B1(new_n908), .B2(new_n925), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n917), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n733), .B2(new_n839), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n314), .A2(new_n912), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1138), .A2(new_n914), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n314), .A2(KEYINPUT97), .A3(new_n912), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n948), .B1(new_n314), .B2(new_n341), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1139), .A2(new_n1140), .B1(new_n1141), .B2(new_n911), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1135), .B1(new_n1137), .B2(new_n1142), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n840), .A2(new_n917), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n938), .B1(new_n1144), .B2(new_n1142), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(KEYINPUT99), .A2(new_n926), .B1(new_n909), .B2(KEYINPUT39), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1145), .A2(new_n930), .A3(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1147), .A3(new_n1120), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n474), .A2(new_n754), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n669), .A2(new_n940), .A3(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n754), .A2(new_n839), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1151), .A2(new_n1142), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n1120), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1153), .A2(new_n918), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1137), .A2(new_n1120), .A3(new_n1152), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND4_X1  g0956(.A1(new_n1134), .A2(new_n1148), .A3(new_n1150), .A4(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n1087), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT113), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1157), .A2(KEYINPUT113), .A3(new_n1087), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1134), .A2(new_n1148), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  NAND3_X1  g0964(.A1(new_n1160), .A2(new_n1161), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n932), .A2(new_n770), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n844), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n819), .B1(new_n402), .B2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n781), .A2(new_n863), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(KEYINPUT54), .B(G143), .ZN(new_n1170));
  OAI21_X1  g0970(.A(new_n285), .B1(new_n784), .B2(new_n1170), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(G125), .C2(new_n805), .ZN(new_n1172));
  NOR2_X1   g0972(.A1(new_n792), .A2(new_n858), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT53), .ZN(new_n1174));
  AOI22_X1  g0974(.A1(new_n795), .A2(G137), .B1(new_n968), .B2(G50), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G159), .A2(new_n807), .B1(new_n797), .B2(G128), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1172), .A2(new_n1174), .A3(new_n1175), .A4(new_n1176), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n862), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n781), .A2(new_n530), .B1(new_n777), .B2(new_n853), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n1179), .B1(G97), .B2(new_n851), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n797), .A2(G283), .ZN(new_n1181));
  AOI22_X1  g0981(.A1(G77), .A2(new_n807), .B1(new_n795), .B2(G107), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1178), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n281), .B1(new_n792), .B2(new_n223), .ZN(new_n1184));
  XNOR2_X1  g0984(.A(new_n1184), .B(KEYINPUT114), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1177), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1168), .B1(new_n1186), .B2(new_n774), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1166), .A2(new_n1187), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1188), .B1(new_n1162), .B2(new_n1080), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1165), .A2(new_n1190), .ZN(G378));
  NAND2_X1  g0991(.A1(new_n1157), .A2(new_n1150), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n950), .A2(new_n945), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n916), .A2(new_n943), .A3(new_n946), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(G330), .A3(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT115), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n449), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n439), .A2(new_n691), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n449), .A2(new_n1197), .ZN(new_n1202));
  OR3_X1    g1002(.A1(new_n1199), .A2(new_n1201), .A3(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1201), .B1(new_n1199), .B2(new_n1202), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1195), .A2(new_n1196), .A3(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(KEYINPUT115), .B1(new_n951), .B2(G330), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1193), .A2(KEYINPUT115), .A3(G330), .A4(new_n1194), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1205), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  OAI211_X1 g1010(.A(new_n939), .B(new_n1206), .C1(new_n1207), .C2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n1208), .A3(new_n1209), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n939), .B1(new_n1214), .B2(new_n1206), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1192), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT57), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(KEYINPUT57), .B(new_n1192), .C1(new_n1212), .C2(new_n1215), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1218), .A2(new_n1087), .A3(new_n1219), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1029), .B1(new_n1212), .B2(new_n1215), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n818), .B1(new_n201), .B2(new_n844), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G150), .A2(new_n807), .B1(new_n797), .B2(G125), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1223), .B1(new_n863), .B2(new_n796), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n792), .A2(new_n1170), .ZN(new_n1225));
  INV_X1    g1025(.A(G128), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n781), .A2(new_n1226), .B1(new_n784), .B2(new_n857), .ZN(new_n1227));
  NOR3_X1   g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1227), .ZN(new_n1228));
  INV_X1    g1028(.A(KEYINPUT59), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n968), .A2(G159), .ZN(new_n1232));
  AOI211_X1 g1032(.A(G33), .B(G41), .C1(new_n805), .C2(G124), .ZN(new_n1233));
  NAND4_X1  g1033(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .A4(new_n1233), .ZN(new_n1234));
  AOI22_X1  g1034(.A1(new_n782), .A2(G107), .B1(new_n851), .B2(new_n462), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1235), .B1(new_n849), .B2(new_n777), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n978), .B(new_n1236), .C1(G77), .C2(new_n808), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n796), .A2(new_n228), .B1(new_n798), .B2(new_n530), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1238), .B1(G58), .B2(new_n968), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1237), .A2(new_n251), .A3(new_n508), .A4(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT58), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G50), .B1(new_n277), .B2(new_n251), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1243), .B1(new_n370), .B2(G41), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1240), .A2(new_n1241), .ZN(new_n1245));
  AND4_X1   g1045(.A1(new_n1234), .A2(new_n1242), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI221_X1 g1046(.A(new_n1222), .B1(new_n846), .B2(new_n1246), .C1(new_n1205), .C2(new_n771), .ZN(new_n1247));
  AND2_X1   g1047(.A1(new_n1221), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1220), .A2(new_n1248), .ZN(G375));
  AOI21_X1  g1049(.A(new_n1144), .B1(new_n1152), .B2(new_n1120), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1152), .A2(new_n1120), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1250), .B1(new_n1137), .B2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n669), .A2(new_n940), .A3(new_n1149), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1163), .A3(new_n1047), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(new_n916), .A2(new_n771), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1256), .B(KEYINPUT116), .ZN(new_n1257));
  OAI22_X1  g1057(.A1(new_n792), .A2(new_n380), .B1(new_n777), .B2(new_n1226), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT120), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n508), .B1(G150), .B2(new_n851), .ZN(new_n1260));
  AOI22_X1  g1060(.A1(new_n807), .A2(G50), .B1(new_n968), .B2(G58), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  XOR2_X1   g1062(.A(new_n1262), .B(KEYINPUT121), .Z(new_n1263));
  OAI22_X1  g1063(.A1(new_n796), .A2(new_n1170), .B1(new_n857), .B2(new_n781), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT119), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n798), .B2(new_n863), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n797), .A2(KEYINPUT119), .A3(G132), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1264), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n797), .A2(G294), .B1(new_n851), .B2(G107), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1269), .B1(new_n530), .B2(new_n796), .ZN(new_n1270));
  XNOR2_X1  g1070(.A(new_n1270), .B(KEYINPUT117), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n788), .A2(new_n221), .ZN(new_n1272));
  OAI22_X1  g1072(.A1(new_n792), .A2(new_n228), .B1(new_n777), .B2(new_n539), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(new_n1273), .B(KEYINPUT118), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n281), .B1(new_n781), .B2(new_n849), .ZN(new_n1275));
  NOR4_X1   g1075(.A1(new_n1272), .A2(new_n1062), .A3(new_n1274), .A4(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1263), .A2(new_n1268), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n819), .B1(G68), .B2(new_n1167), .C1(new_n1277), .C2(new_n846), .ZN(new_n1278));
  OAI22_X1  g1078(.A1(new_n1252), .A2(new_n1080), .B1(new_n1257), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1255), .A2(new_n1280), .ZN(new_n1281));
  XOR2_X1   g1081(.A(new_n1281), .B(KEYINPUT122), .Z(new_n1282));
  INV_X1    g1082(.A(new_n1282), .ZN(G381));
  INV_X1    g1083(.A(G375), .ZN(new_n1284));
  AOI22_X1  g1084(.A1(new_n1158), .A2(new_n1159), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n1189), .B1(new_n1285), .B2(new_n1161), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1118), .A2(new_n870), .ZN(new_n1287));
  INV_X1    g1087(.A(G396), .ZN(new_n1288));
  OAI211_X1 g1088(.A(new_n1083), .B(new_n1288), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1287), .A2(G387), .A3(new_n1289), .ZN(new_n1290));
  NAND4_X1  g1090(.A1(new_n1284), .A2(new_n1286), .A3(new_n1282), .A4(new_n1290), .ZN(G407));
  NAND2_X1  g1091(.A1(new_n692), .A2(G213), .ZN(new_n1292));
  XOR2_X1   g1092(.A(new_n1292), .B(KEYINPUT123), .Z(new_n1293));
  NAND3_X1  g1093(.A1(new_n1284), .A2(new_n1286), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G407), .A2(G213), .A3(new_n1294), .ZN(G409));
  NAND2_X1  g1095(.A1(new_n1293), .A2(G2897), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(KEYINPUT60), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1299));
  OAI21_X1  g1099(.A(KEYINPUT124), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT60), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1301), .B1(new_n1150), .B2(new_n1156), .ZN(new_n1302));
  INV_X1    g1102(.A(KEYINPUT124), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1302), .A2(new_n1303), .A3(new_n1163), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1300), .A2(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1253), .A2(KEYINPUT60), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT125), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1252), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1253), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1308), .A2(new_n1087), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1305), .A2(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(G384), .B1(new_n1311), .B2(new_n1280), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n870), .B(new_n1279), .C1(new_n1305), .C2(new_n1310), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1297), .B1(new_n1312), .B2(new_n1313), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1308), .A2(new_n1087), .A3(new_n1309), .ZN(new_n1315));
  AOI21_X1  g1115(.A(new_n1315), .B1(new_n1304), .B2(new_n1300), .ZN(new_n1316));
  OAI21_X1  g1116(.A(new_n870), .B1(new_n1316), .B2(new_n1279), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1311), .A2(G384), .A3(new_n1280), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1317), .A2(new_n1318), .A3(new_n1296), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1314), .A2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(new_n1320), .ZN(new_n1321));
  OAI21_X1  g1121(.A(new_n1206), .B1(new_n1207), .B2(new_n1210), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n939), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  AOI22_X1  g1124(.A1(new_n1324), .A2(new_n1211), .B1(new_n1150), .B2(new_n1157), .ZN(new_n1325));
  OAI21_X1  g1125(.A(new_n1087), .B1(new_n1325), .B2(KEYINPUT57), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1219), .ZN(new_n1327));
  OAI211_X1 g1127(.A(G378), .B(new_n1248), .C1(new_n1326), .C2(new_n1327), .ZN(new_n1328));
  OAI211_X1 g1128(.A(new_n1221), .B(new_n1247), .C1(new_n1216), .C2(new_n1046), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(new_n1286), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1328), .A2(new_n1330), .ZN(new_n1331));
  INV_X1    g1131(.A(new_n1293), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT61), .B1(new_n1321), .B2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(KEYINPUT63), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1312), .A2(new_n1313), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1333), .B2(new_n1337), .ZN(new_n1338));
  INV_X1    g1138(.A(KEYINPUT126), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(G393), .A2(G396), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1340), .A2(new_n1289), .ZN(new_n1341));
  INV_X1    g1141(.A(new_n992), .ZN(new_n1342));
  AND3_X1   g1142(.A1(new_n1017), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1026), .B1(new_n1017), .B2(new_n1022), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1080), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n1342), .B1(new_n1345), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1348), .A2(G390), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(G387), .A2(new_n1118), .ZN(new_n1350));
  AND4_X1   g1150(.A1(new_n1339), .A2(new_n1341), .A3(new_n1349), .A4(new_n1350), .ZN(new_n1351));
  OAI21_X1  g1151(.A(KEYINPUT126), .B1(new_n1348), .B2(G390), .ZN(new_n1352));
  AOI22_X1  g1152(.A1(new_n1352), .A2(new_n1341), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1353));
  NOR2_X1   g1153(.A1(new_n1351), .A2(new_n1353), .ZN(new_n1354));
  INV_X1    g1154(.A(new_n1354), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1293), .B1(new_n1328), .B2(new_n1330), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1356), .A2(KEYINPUT63), .A3(new_n1336), .ZN(new_n1357));
  NAND4_X1  g1157(.A1(new_n1334), .A2(new_n1338), .A3(new_n1355), .A4(new_n1357), .ZN(new_n1358));
  INV_X1    g1158(.A(KEYINPUT62), .ZN(new_n1359));
  AND3_X1   g1159(.A1(new_n1356), .A2(new_n1359), .A3(new_n1336), .ZN(new_n1360));
  INV_X1    g1160(.A(KEYINPUT61), .ZN(new_n1361));
  OAI21_X1  g1161(.A(new_n1361), .B1(new_n1356), .B2(new_n1320), .ZN(new_n1362));
  AOI21_X1  g1162(.A(new_n1359), .B1(new_n1356), .B2(new_n1336), .ZN(new_n1363));
  NOR3_X1   g1163(.A1(new_n1360), .A2(new_n1362), .A3(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1358), .B1(new_n1364), .B2(new_n1355), .ZN(G405));
  AOI21_X1  g1165(.A(G378), .B1(new_n1220), .B2(new_n1248), .ZN(new_n1366));
  INV_X1    g1166(.A(new_n1366), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1367), .A2(new_n1328), .A3(new_n1337), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1328), .ZN(new_n1369));
  OAI21_X1  g1169(.A(new_n1336), .B1(new_n1369), .B2(new_n1366), .ZN(new_n1370));
  NAND3_X1  g1170(.A1(new_n1354), .A2(new_n1368), .A3(new_n1370), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1371), .A2(KEYINPUT127), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT127), .ZN(new_n1373));
  NAND4_X1  g1173(.A1(new_n1354), .A2(new_n1368), .A3(new_n1370), .A4(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1368), .A2(new_n1370), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1375), .A2(new_n1355), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1372), .A2(new_n1374), .A3(new_n1376), .ZN(G402));
endmodule


