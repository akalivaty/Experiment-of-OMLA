

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n566), .A2(n523), .ZN(n797) );
  XNOR2_X2 U551 ( .A(n593), .B(n592), .ZN(n705) );
  BUF_X1 U552 ( .A(n892), .Z(n516) );
  BUF_X1 U553 ( .A(n892), .Z(n517) );
  NOR2_X1 U554 ( .A1(n678), .A2(n677), .ZN(n692) );
  INV_X1 U555 ( .A(n662), .ZN(n518) );
  OR2_X1 U556 ( .A1(n692), .A2(n681), .ZN(n688) );
  NOR2_X1 U557 ( .A1(n635), .A2(n945), .ZN(n629) );
  NOR2_X1 U558 ( .A1(n660), .A2(n659), .ZN(n661) );
  AND2_X1 U559 ( .A1(n696), .A2(n699), .ZN(n702) );
  INV_X1 U560 ( .A(KEYINPUT13), .ZN(n612) );
  XOR2_X1 U561 ( .A(KEYINPUT65), .B(n524), .Z(n801) );
  XNOR2_X1 U562 ( .A(n613), .B(n612), .ZN(n614) );
  NOR2_X1 U563 ( .A1(G651), .A2(n566), .ZN(n800) );
  INV_X1 U564 ( .A(G651), .ZN(n523) );
  NOR2_X1 U565 ( .A1(G543), .A2(n523), .ZN(n519) );
  XOR2_X1 U566 ( .A(KEYINPUT1), .B(n519), .Z(n796) );
  NAND2_X1 U567 ( .A1(G65), .A2(n796), .ZN(n521) );
  XOR2_X1 U568 ( .A(G543), .B(KEYINPUT0), .Z(n566) );
  NAND2_X1 U569 ( .A1(G53), .A2(n800), .ZN(n520) );
  NAND2_X1 U570 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U571 ( .A(KEYINPUT69), .B(n522), .ZN(n528) );
  NAND2_X1 U572 ( .A1(G78), .A2(n797), .ZN(n526) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n524) );
  NAND2_X1 U574 ( .A1(G91), .A2(n801), .ZN(n525) );
  AND2_X1 U575 ( .A1(n526), .A2(n525), .ZN(n527) );
  NAND2_X1 U576 ( .A1(n528), .A2(n527), .ZN(G299) );
  INV_X1 U577 ( .A(G2105), .ZN(n532) );
  AND2_X1 U578 ( .A1(n532), .A2(G2104), .ZN(n898) );
  NAND2_X1 U579 ( .A1(G102), .A2(n898), .ZN(n531) );
  NOR2_X1 U580 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  XOR2_X2 U581 ( .A(KEYINPUT17), .B(n529), .Z(n896) );
  NAND2_X1 U582 ( .A1(G138), .A2(n896), .ZN(n530) );
  NAND2_X1 U583 ( .A1(n531), .A2(n530), .ZN(n536) );
  AND2_X1 U584 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U585 ( .A1(G114), .A2(n891), .ZN(n534) );
  NOR2_X1 U586 ( .A1(G2104), .A2(n532), .ZN(n892) );
  NAND2_X1 U587 ( .A1(G126), .A2(n517), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n536), .A2(n535), .ZN(G164) );
  NAND2_X1 U590 ( .A1(G77), .A2(n797), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G90), .A2(n801), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U593 ( .A(KEYINPUT9), .B(n539), .ZN(n543) );
  NAND2_X1 U594 ( .A1(G64), .A2(n796), .ZN(n541) );
  NAND2_X1 U595 ( .A1(G52), .A2(n800), .ZN(n540) );
  AND2_X1 U596 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U597 ( .A1(n543), .A2(n542), .ZN(G301) );
  INV_X1 U598 ( .A(G301), .ZN(G171) );
  NAND2_X1 U599 ( .A1(G63), .A2(n796), .ZN(n545) );
  NAND2_X1 U600 ( .A1(G51), .A2(n800), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U602 ( .A(n546), .B(KEYINPUT75), .ZN(n547) );
  XNOR2_X1 U603 ( .A(n547), .B(KEYINPUT6), .ZN(n554) );
  XNOR2_X1 U604 ( .A(KEYINPUT74), .B(KEYINPUT5), .ZN(n552) );
  NAND2_X1 U605 ( .A1(n801), .A2(G89), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT4), .ZN(n550) );
  NAND2_X1 U607 ( .A1(G76), .A2(n797), .ZN(n549) );
  NAND2_X1 U608 ( .A1(n550), .A2(n549), .ZN(n551) );
  XNOR2_X1 U609 ( .A(n552), .B(n551), .ZN(n553) );
  NAND2_X1 U610 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U611 ( .A(KEYINPUT7), .B(n555), .ZN(G168) );
  XOR2_X1 U612 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U613 ( .A1(G62), .A2(n796), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G75), .A2(n797), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n560) );
  NAND2_X1 U616 ( .A1(n801), .A2(G88), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT80), .B(n558), .Z(n559) );
  NOR2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n800), .A2(G50), .ZN(n561) );
  NAND2_X1 U620 ( .A1(n562), .A2(n561), .ZN(G303) );
  NAND2_X1 U621 ( .A1(G49), .A2(n800), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U624 ( .A1(n796), .A2(n565), .ZN(n568) );
  NAND2_X1 U625 ( .A1(n566), .A2(G87), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n568), .A2(n567), .ZN(G288) );
  NAND2_X1 U627 ( .A1(G73), .A2(n797), .ZN(n569) );
  XNOR2_X1 U628 ( .A(n569), .B(KEYINPUT2), .ZN(n576) );
  NAND2_X1 U629 ( .A1(G61), .A2(n796), .ZN(n571) );
  NAND2_X1 U630 ( .A1(G86), .A2(n801), .ZN(n570) );
  NAND2_X1 U631 ( .A1(n571), .A2(n570), .ZN(n574) );
  NAND2_X1 U632 ( .A1(G48), .A2(n800), .ZN(n572) );
  XNOR2_X1 U633 ( .A(KEYINPUT79), .B(n572), .ZN(n573) );
  NOR2_X1 U634 ( .A1(n574), .A2(n573), .ZN(n575) );
  NAND2_X1 U635 ( .A1(n576), .A2(n575), .ZN(G305) );
  NAND2_X1 U636 ( .A1(n796), .A2(G60), .ZN(n577) );
  XNOR2_X1 U637 ( .A(n577), .B(KEYINPUT66), .ZN(n579) );
  NAND2_X1 U638 ( .A1(G47), .A2(n800), .ZN(n578) );
  NAND2_X1 U639 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U640 ( .A(KEYINPUT67), .B(n580), .ZN(n584) );
  NAND2_X1 U641 ( .A1(G72), .A2(n797), .ZN(n582) );
  NAND2_X1 U642 ( .A1(G85), .A2(n801), .ZN(n581) );
  AND2_X1 U643 ( .A1(n582), .A2(n581), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n584), .A2(n583), .ZN(G290) );
  INV_X1 U645 ( .A(KEYINPUT94), .ZN(n594) );
  NOR2_X1 U646 ( .A1(G164), .A2(G1384), .ZN(n706) );
  NAND2_X1 U647 ( .A1(n896), .A2(G137), .ZN(n587) );
  NAND2_X1 U648 ( .A1(G101), .A2(n898), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT23), .B(n585), .Z(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(n779) );
  INV_X1 U651 ( .A(G40), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G113), .A2(n891), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G125), .A2(n516), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n778) );
  OR2_X1 U655 ( .A1(n590), .A2(n778), .ZN(n591) );
  OR2_X1 U656 ( .A1(n779), .A2(n591), .ZN(n593) );
  INV_X1 U657 ( .A(KEYINPUT86), .ZN(n592) );
  NAND2_X2 U658 ( .A1(n706), .A2(n705), .ZN(n662) );
  NAND2_X1 U659 ( .A1(n594), .A2(n662), .ZN(n596) );
  NAND2_X1 U660 ( .A1(KEYINPUT94), .A2(n518), .ZN(n595) );
  NAND2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G2072), .A2(n598), .ZN(n597) );
  XOR2_X1 U663 ( .A(KEYINPUT27), .B(n597), .Z(n601) );
  BUF_X1 U664 ( .A(n598), .Z(n599) );
  INV_X1 U665 ( .A(n599), .ZN(n630) );
  NAND2_X1 U666 ( .A1(n630), .A2(G1956), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n640) );
  NOR2_X1 U668 ( .A1(G299), .A2(n640), .ZN(n602) );
  XOR2_X1 U669 ( .A(n602), .B(KEYINPUT96), .Z(n639) );
  XOR2_X1 U670 ( .A(KEYINPUT64), .B(KEYINPUT26), .Z(n604) );
  NAND2_X1 U671 ( .A1(n518), .A2(G1996), .ZN(n603) );
  XNOR2_X1 U672 ( .A(n604), .B(n603), .ZN(n618) );
  XOR2_X1 U673 ( .A(KEYINPUT14), .B(KEYINPUT70), .Z(n606) );
  NAND2_X1 U674 ( .A1(G56), .A2(n796), .ZN(n605) );
  XNOR2_X1 U675 ( .A(n606), .B(n605), .ZN(n615) );
  NAND2_X1 U676 ( .A1(n797), .A2(G68), .ZN(n607) );
  XNOR2_X1 U677 ( .A(KEYINPUT72), .B(n607), .ZN(n611) );
  XOR2_X1 U678 ( .A(KEYINPUT12), .B(KEYINPUT71), .Z(n609) );
  NAND2_X1 U679 ( .A1(G81), .A2(n801), .ZN(n608) );
  XNOR2_X1 U680 ( .A(n609), .B(n608), .ZN(n610) );
  NAND2_X1 U681 ( .A1(n611), .A2(n610), .ZN(n613) );
  NOR2_X1 U682 ( .A1(n615), .A2(n614), .ZN(n617) );
  NAND2_X1 U683 ( .A1(n800), .A2(G43), .ZN(n616) );
  NAND2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n952) );
  NOR2_X1 U685 ( .A1(n618), .A2(n952), .ZN(n620) );
  NAND2_X1 U686 ( .A1(G1341), .A2(n662), .ZN(n619) );
  NAND2_X1 U687 ( .A1(n620), .A2(n619), .ZN(n635) );
  NAND2_X1 U688 ( .A1(n800), .A2(G54), .ZN(n627) );
  NAND2_X1 U689 ( .A1(G79), .A2(n797), .ZN(n622) );
  NAND2_X1 U690 ( .A1(G92), .A2(n801), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n622), .A2(n621), .ZN(n625) );
  NAND2_X1 U692 ( .A1(G66), .A2(n796), .ZN(n623) );
  XNOR2_X1 U693 ( .A(KEYINPUT73), .B(n623), .ZN(n624) );
  NOR2_X1 U694 ( .A1(n625), .A2(n624), .ZN(n626) );
  NAND2_X1 U695 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U696 ( .A(KEYINPUT15), .B(n628), .Z(n945) );
  XNOR2_X1 U697 ( .A(n629), .B(KEYINPUT95), .ZN(n634) );
  NAND2_X1 U698 ( .A1(G1348), .A2(n662), .ZN(n632) );
  NAND2_X1 U699 ( .A1(G2067), .A2(n599), .ZN(n631) );
  NAND2_X1 U700 ( .A1(n632), .A2(n631), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n634), .A2(n633), .ZN(n637) );
  NAND2_X1 U702 ( .A1(n945), .A2(n635), .ZN(n636) );
  NAND2_X1 U703 ( .A1(n637), .A2(n636), .ZN(n638) );
  NAND2_X1 U704 ( .A1(n639), .A2(n638), .ZN(n643) );
  NAND2_X1 U705 ( .A1(G299), .A2(n640), .ZN(n641) );
  XNOR2_X1 U706 ( .A(n641), .B(KEYINPUT28), .ZN(n642) );
  NAND2_X1 U707 ( .A1(n643), .A2(n642), .ZN(n645) );
  XOR2_X1 U708 ( .A(KEYINPUT29), .B(KEYINPUT97), .Z(n644) );
  XNOR2_X1 U709 ( .A(n645), .B(n644), .ZN(n649) );
  XNOR2_X1 U710 ( .A(KEYINPUT25), .B(G2078), .ZN(n981) );
  NAND2_X1 U711 ( .A1(n599), .A2(n981), .ZN(n647) );
  INV_X1 U712 ( .A(G1961), .ZN(n918) );
  NAND2_X1 U713 ( .A1(n918), .A2(n662), .ZN(n646) );
  NAND2_X1 U714 ( .A1(n647), .A2(n646), .ZN(n655) );
  AND2_X1 U715 ( .A1(n655), .A2(G171), .ZN(n648) );
  NOR2_X1 U716 ( .A1(n649), .A2(n648), .ZN(n650) );
  XNOR2_X1 U717 ( .A(n650), .B(KEYINPUT98), .ZN(n660) );
  NAND2_X1 U718 ( .A1(G8), .A2(n662), .ZN(n699) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n699), .ZN(n676) );
  NOR2_X1 U720 ( .A1(G2084), .A2(n662), .ZN(n651) );
  XNOR2_X1 U721 ( .A(KEYINPUT93), .B(n651), .ZN(n671) );
  NAND2_X1 U722 ( .A1(G8), .A2(n671), .ZN(n652) );
  NOR2_X1 U723 ( .A1(n676), .A2(n652), .ZN(n653) );
  XOR2_X1 U724 ( .A(KEYINPUT30), .B(n653), .Z(n654) );
  NOR2_X1 U725 ( .A1(G168), .A2(n654), .ZN(n657) );
  NOR2_X1 U726 ( .A1(G171), .A2(n655), .ZN(n656) );
  NOR2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U728 ( .A(KEYINPUT31), .B(n658), .ZN(n659) );
  XNOR2_X1 U729 ( .A(n661), .B(KEYINPUT99), .ZN(n674) );
  NAND2_X1 U730 ( .A1(n674), .A2(G286), .ZN(n669) );
  INV_X1 U731 ( .A(G8), .ZN(n667) );
  NOR2_X1 U732 ( .A1(G1971), .A2(n699), .ZN(n664) );
  NOR2_X1 U733 ( .A1(G2090), .A2(n662), .ZN(n663) );
  NOR2_X1 U734 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U735 ( .A1(n665), .A2(G303), .ZN(n666) );
  OR2_X1 U736 ( .A1(n667), .A2(n666), .ZN(n668) );
  AND2_X1 U737 ( .A1(n669), .A2(n668), .ZN(n670) );
  XOR2_X1 U738 ( .A(n670), .B(KEYINPUT32), .Z(n678) );
  INV_X1 U739 ( .A(n671), .ZN(n672) );
  NAND2_X1 U740 ( .A1(G8), .A2(n672), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U742 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U743 ( .A1(G1971), .A2(G303), .ZN(n947) );
  XOR2_X1 U744 ( .A(n947), .B(KEYINPUT100), .Z(n680) );
  NOR2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n957) );
  INV_X1 U746 ( .A(n957), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  INV_X1 U748 ( .A(n699), .ZN(n682) );
  NAND2_X1 U749 ( .A1(G1976), .A2(G288), .ZN(n948) );
  AND2_X1 U750 ( .A1(n682), .A2(n948), .ZN(n686) );
  NAND2_X1 U751 ( .A1(n957), .A2(KEYINPUT33), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n683), .A2(n699), .ZN(n685) );
  XOR2_X1 U753 ( .A(G1981), .B(G305), .Z(n964) );
  INV_X1 U754 ( .A(n964), .ZN(n684) );
  NOR2_X1 U755 ( .A1(n685), .A2(n684), .ZN(n689) );
  AND2_X1 U756 ( .A1(n686), .A2(n689), .ZN(n687) );
  NAND2_X1 U757 ( .A1(n688), .A2(n687), .ZN(n691) );
  NAND2_X1 U758 ( .A1(n689), .A2(KEYINPUT33), .ZN(n690) );
  AND2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n704) );
  INV_X1 U760 ( .A(n692), .ZN(n695) );
  NOR2_X1 U761 ( .A1(G2090), .A2(G303), .ZN(n693) );
  NAND2_X1 U762 ( .A1(G8), .A2(n693), .ZN(n694) );
  NAND2_X1 U763 ( .A1(n695), .A2(n694), .ZN(n696) );
  NOR2_X1 U764 ( .A1(G1981), .A2(G305), .ZN(n697) );
  XOR2_X1 U765 ( .A(n697), .B(KEYINPUT24), .Z(n698) );
  NOR2_X1 U766 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U767 ( .A(n700), .B(KEYINPUT92), .ZN(n701) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n741) );
  INV_X1 U770 ( .A(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n707), .A2(n706), .ZN(n752) );
  XNOR2_X1 U772 ( .A(G2067), .B(KEYINPUT37), .ZN(n749) );
  NAND2_X1 U773 ( .A1(G104), .A2(n898), .ZN(n709) );
  NAND2_X1 U774 ( .A1(G140), .A2(n896), .ZN(n708) );
  NAND2_X1 U775 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U776 ( .A(KEYINPUT34), .B(n710), .ZN(n716) );
  NAND2_X1 U777 ( .A1(G116), .A2(n891), .ZN(n712) );
  NAND2_X1 U778 ( .A1(G128), .A2(n517), .ZN(n711) );
  NAND2_X1 U779 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U780 ( .A(KEYINPUT35), .B(n713), .ZN(n714) );
  XNOR2_X1 U781 ( .A(KEYINPUT87), .B(n714), .ZN(n715) );
  NOR2_X1 U782 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U783 ( .A(KEYINPUT36), .B(n717), .ZN(n906) );
  NOR2_X1 U784 ( .A1(n749), .A2(n906), .ZN(n718) );
  XNOR2_X1 U785 ( .A(n718), .B(KEYINPUT88), .ZN(n1022) );
  NAND2_X1 U786 ( .A1(n752), .A2(n1022), .ZN(n747) );
  NAND2_X1 U787 ( .A1(G107), .A2(n891), .ZN(n720) );
  NAND2_X1 U788 ( .A1(G119), .A2(n517), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n725) );
  NAND2_X1 U790 ( .A1(G95), .A2(n898), .ZN(n722) );
  NAND2_X1 U791 ( .A1(G131), .A2(n896), .ZN(n721) );
  NAND2_X1 U792 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U793 ( .A(KEYINPUT89), .B(n723), .Z(n724) );
  NOR2_X1 U794 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U795 ( .A(KEYINPUT90), .B(n726), .Z(n907) );
  NAND2_X1 U796 ( .A1(G1991), .A2(n907), .ZN(n735) );
  NAND2_X1 U797 ( .A1(G141), .A2(n896), .ZN(n728) );
  NAND2_X1 U798 ( .A1(G129), .A2(n517), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n731) );
  NAND2_X1 U800 ( .A1(n898), .A2(G105), .ZN(n729) );
  XOR2_X1 U801 ( .A(KEYINPUT38), .B(n729), .Z(n730) );
  NOR2_X1 U802 ( .A1(n731), .A2(n730), .ZN(n733) );
  NAND2_X1 U803 ( .A1(n891), .A2(G117), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n886) );
  NAND2_X1 U805 ( .A1(G1996), .A2(n886), .ZN(n734) );
  NAND2_X1 U806 ( .A1(n735), .A2(n734), .ZN(n1008) );
  NAND2_X1 U807 ( .A1(n752), .A2(n1008), .ZN(n736) );
  XNOR2_X1 U808 ( .A(KEYINPUT91), .B(n736), .ZN(n744) );
  INV_X1 U809 ( .A(n744), .ZN(n737) );
  NAND2_X1 U810 ( .A1(n747), .A2(n737), .ZN(n739) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n963) );
  AND2_X1 U812 ( .A1(n963), .A2(n752), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n755) );
  NOR2_X1 U815 ( .A1(G1996), .A2(n886), .ZN(n1001) );
  NOR2_X1 U816 ( .A1(G1986), .A2(G290), .ZN(n742) );
  NOR2_X1 U817 ( .A1(G1991), .A2(n907), .ZN(n1014) );
  NOR2_X1 U818 ( .A1(n742), .A2(n1014), .ZN(n743) );
  NOR2_X1 U819 ( .A1(n744), .A2(n743), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n1001), .A2(n745), .ZN(n746) );
  XNOR2_X1 U821 ( .A(KEYINPUT39), .B(n746), .ZN(n748) );
  NAND2_X1 U822 ( .A1(n748), .A2(n747), .ZN(n751) );
  AND2_X1 U823 ( .A1(n749), .A2(n906), .ZN(n750) );
  XNOR2_X1 U824 ( .A(n750), .B(KEYINPUT101), .ZN(n1019) );
  NAND2_X1 U825 ( .A1(n751), .A2(n1019), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U827 ( .A1(n755), .A2(n754), .ZN(n756) );
  XNOR2_X1 U828 ( .A(n756), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U829 ( .A(G2443), .B(G2435), .ZN(n766) );
  XOR2_X1 U830 ( .A(G2427), .B(KEYINPUT103), .Z(n758) );
  XNOR2_X1 U831 ( .A(G2454), .B(G2430), .ZN(n757) );
  XNOR2_X1 U832 ( .A(n758), .B(n757), .ZN(n762) );
  XOR2_X1 U833 ( .A(KEYINPUT102), .B(G2446), .Z(n760) );
  XNOR2_X1 U834 ( .A(G1348), .B(G1341), .ZN(n759) );
  XNOR2_X1 U835 ( .A(n760), .B(n759), .ZN(n761) );
  XOR2_X1 U836 ( .A(n762), .B(n761), .Z(n764) );
  XNOR2_X1 U837 ( .A(G2451), .B(G2438), .ZN(n763) );
  XNOR2_X1 U838 ( .A(n764), .B(n763), .ZN(n765) );
  XNOR2_X1 U839 ( .A(n766), .B(n765), .ZN(n767) );
  AND2_X1 U840 ( .A1(n767), .A2(G14), .ZN(G401) );
  NAND2_X1 U841 ( .A1(G123), .A2(n517), .ZN(n768) );
  XNOR2_X1 U842 ( .A(n768), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U843 ( .A1(n898), .A2(G99), .ZN(n769) );
  XNOR2_X1 U844 ( .A(n769), .B(KEYINPUT78), .ZN(n771) );
  NAND2_X1 U845 ( .A1(G135), .A2(n896), .ZN(n770) );
  NAND2_X1 U846 ( .A1(n771), .A2(n770), .ZN(n774) );
  NAND2_X1 U847 ( .A1(G111), .A2(n891), .ZN(n772) );
  XNOR2_X1 U848 ( .A(KEYINPUT77), .B(n772), .ZN(n773) );
  NOR2_X1 U849 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U850 ( .A1(n776), .A2(n775), .ZN(n1012) );
  XNOR2_X1 U851 ( .A(G2096), .B(n1012), .ZN(n777) );
  OR2_X1 U852 ( .A1(G2100), .A2(n777), .ZN(G156) );
  INV_X1 U853 ( .A(G108), .ZN(G238) );
  INV_X1 U854 ( .A(G120), .ZN(G236) );
  INV_X1 U855 ( .A(G69), .ZN(G235) );
  INV_X1 U856 ( .A(G132), .ZN(G219) );
  INV_X1 U857 ( .A(G82), .ZN(G220) );
  NOR2_X1 U858 ( .A1(n779), .A2(n778), .ZN(G160) );
  NAND2_X1 U859 ( .A1(G94), .A2(G452), .ZN(n780) );
  XOR2_X1 U860 ( .A(KEYINPUT68), .B(n780), .Z(G173) );
  NAND2_X1 U861 ( .A1(G7), .A2(G661), .ZN(n781) );
  XNOR2_X1 U862 ( .A(n781), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U863 ( .A(G223), .ZN(n836) );
  NAND2_X1 U864 ( .A1(n836), .A2(G567), .ZN(n782) );
  XOR2_X1 U865 ( .A(KEYINPUT11), .B(n782), .Z(G234) );
  INV_X1 U866 ( .A(G860), .ZN(n787) );
  OR2_X1 U867 ( .A1(n952), .A2(n787), .ZN(G153) );
  NAND2_X1 U868 ( .A1(G868), .A2(G301), .ZN(n784) );
  INV_X1 U869 ( .A(G868), .ZN(n816) );
  NAND2_X1 U870 ( .A1(n945), .A2(n816), .ZN(n783) );
  NAND2_X1 U871 ( .A1(n784), .A2(n783), .ZN(G284) );
  NOR2_X1 U872 ( .A1(G286), .A2(n816), .ZN(n786) );
  NOR2_X1 U873 ( .A1(G868), .A2(G299), .ZN(n785) );
  NOR2_X1 U874 ( .A1(n786), .A2(n785), .ZN(G297) );
  NAND2_X1 U875 ( .A1(n787), .A2(G559), .ZN(n788) );
  INV_X1 U876 ( .A(n945), .ZN(n794) );
  NAND2_X1 U877 ( .A1(n788), .A2(n794), .ZN(n789) );
  XNOR2_X1 U878 ( .A(n789), .B(KEYINPUT76), .ZN(n790) );
  XNOR2_X1 U879 ( .A(KEYINPUT16), .B(n790), .ZN(G148) );
  NOR2_X1 U880 ( .A1(G868), .A2(n952), .ZN(n793) );
  NAND2_X1 U881 ( .A1(G868), .A2(n794), .ZN(n791) );
  NOR2_X1 U882 ( .A1(G559), .A2(n791), .ZN(n792) );
  NOR2_X1 U883 ( .A1(n793), .A2(n792), .ZN(G282) );
  NAND2_X1 U884 ( .A1(n794), .A2(G559), .ZN(n814) );
  XNOR2_X1 U885 ( .A(n952), .B(n814), .ZN(n795) );
  NOR2_X1 U886 ( .A1(n795), .A2(G860), .ZN(n806) );
  NAND2_X1 U887 ( .A1(G67), .A2(n796), .ZN(n799) );
  NAND2_X1 U888 ( .A1(G80), .A2(n797), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G55), .A2(n800), .ZN(n803) );
  NAND2_X1 U891 ( .A1(G93), .A2(n801), .ZN(n802) );
  NAND2_X1 U892 ( .A1(n803), .A2(n802), .ZN(n804) );
  OR2_X1 U893 ( .A1(n805), .A2(n804), .ZN(n817) );
  XOR2_X1 U894 ( .A(n806), .B(n817), .Z(G145) );
  XNOR2_X1 U895 ( .A(G290), .B(n952), .ZN(n813) );
  XOR2_X1 U896 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n807) );
  XNOR2_X1 U897 ( .A(G288), .B(n807), .ZN(n810) );
  XOR2_X1 U898 ( .A(n817), .B(G299), .Z(n808) );
  XNOR2_X1 U899 ( .A(n808), .B(G303), .ZN(n809) );
  XNOR2_X1 U900 ( .A(n810), .B(n809), .ZN(n811) );
  XNOR2_X1 U901 ( .A(n811), .B(G305), .ZN(n812) );
  XNOR2_X1 U902 ( .A(n813), .B(n812), .ZN(n844) );
  XNOR2_X1 U903 ( .A(n814), .B(n844), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n815), .A2(G868), .ZN(n819) );
  NAND2_X1 U905 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U906 ( .A1(n819), .A2(n818), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2084), .A2(G2078), .ZN(n821) );
  XOR2_X1 U908 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n820) );
  XNOR2_X1 U909 ( .A(n821), .B(n820), .ZN(n822) );
  NAND2_X1 U910 ( .A1(n822), .A2(G2090), .ZN(n823) );
  XOR2_X1 U911 ( .A(KEYINPUT21), .B(n823), .Z(n824) );
  XNOR2_X1 U912 ( .A(KEYINPUT83), .B(n824), .ZN(n825) );
  NAND2_X1 U913 ( .A1(n825), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U915 ( .A1(G220), .A2(G219), .ZN(n826) );
  XOR2_X1 U916 ( .A(KEYINPUT22), .B(n826), .Z(n827) );
  NOR2_X1 U917 ( .A1(G218), .A2(n827), .ZN(n828) );
  NAND2_X1 U918 ( .A1(G96), .A2(n828), .ZN(n842) );
  NAND2_X1 U919 ( .A1(n842), .A2(G2106), .ZN(n834) );
  NOR2_X1 U920 ( .A1(G235), .A2(G236), .ZN(n829) );
  XNOR2_X1 U921 ( .A(KEYINPUT84), .B(n829), .ZN(n830) );
  NAND2_X1 U922 ( .A1(n830), .A2(G57), .ZN(n831) );
  NOR2_X1 U923 ( .A1(n831), .A2(G238), .ZN(n832) );
  XNOR2_X1 U924 ( .A(n832), .B(KEYINPUT85), .ZN(n843) );
  NAND2_X1 U925 ( .A1(n843), .A2(G567), .ZN(n833) );
  NAND2_X1 U926 ( .A1(n834), .A2(n833), .ZN(n917) );
  NAND2_X1 U927 ( .A1(G483), .A2(G661), .ZN(n835) );
  NOR2_X1 U928 ( .A1(n917), .A2(n835), .ZN(n839) );
  NAND2_X1 U929 ( .A1(n839), .A2(G36), .ZN(G176) );
  INV_X1 U930 ( .A(G303), .ZN(G166) );
  NAND2_X1 U931 ( .A1(G2106), .A2(n836), .ZN(G217) );
  NAND2_X1 U932 ( .A1(G15), .A2(G2), .ZN(n837) );
  XOR2_X1 U933 ( .A(KEYINPUT104), .B(n837), .Z(n838) );
  NAND2_X1 U934 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n840) );
  NAND2_X1 U936 ( .A1(n840), .A2(n839), .ZN(n841) );
  XOR2_X1 U937 ( .A(KEYINPUT105), .B(n841), .Z(G188) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  INV_X1 U940 ( .A(G57), .ZN(G237) );
  NOR2_X1 U941 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  XNOR2_X1 U943 ( .A(G286), .B(n945), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n845), .B(n844), .ZN(n846) );
  XNOR2_X1 U945 ( .A(n846), .B(G171), .ZN(n847) );
  NOR2_X1 U946 ( .A1(G37), .A2(n847), .ZN(G397) );
  XNOR2_X1 U947 ( .A(G1996), .B(KEYINPUT41), .ZN(n857) );
  XOR2_X1 U948 ( .A(G1971), .B(G1956), .Z(n849) );
  XNOR2_X1 U949 ( .A(G1991), .B(G1961), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U951 ( .A(G1966), .B(G1976), .Z(n851) );
  XNOR2_X1 U952 ( .A(G1986), .B(G1981), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n852) );
  XOR2_X1 U954 ( .A(n853), .B(n852), .Z(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT108), .B(G2474), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U957 ( .A(n857), .B(n856), .ZN(G229) );
  XOR2_X1 U958 ( .A(KEYINPUT43), .B(G2678), .Z(n859) );
  XNOR2_X1 U959 ( .A(KEYINPUT106), .B(KEYINPUT107), .ZN(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n863) );
  XOR2_X1 U961 ( .A(KEYINPUT42), .B(G2090), .Z(n861) );
  XNOR2_X1 U962 ( .A(G2067), .B(G2072), .ZN(n860) );
  XNOR2_X1 U963 ( .A(n861), .B(n860), .ZN(n862) );
  XOR2_X1 U964 ( .A(n863), .B(n862), .Z(n865) );
  XNOR2_X1 U965 ( .A(G2096), .B(G2100), .ZN(n864) );
  XNOR2_X1 U966 ( .A(n865), .B(n864), .ZN(n867) );
  XOR2_X1 U967 ( .A(G2084), .B(G2078), .Z(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(G227) );
  NAND2_X1 U969 ( .A1(G124), .A2(n517), .ZN(n868) );
  XOR2_X1 U970 ( .A(KEYINPUT109), .B(n868), .Z(n869) );
  XNOR2_X1 U971 ( .A(n869), .B(KEYINPUT44), .ZN(n871) );
  NAND2_X1 U972 ( .A1(G100), .A2(n898), .ZN(n870) );
  NAND2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n875) );
  NAND2_X1 U974 ( .A1(G136), .A2(n896), .ZN(n873) );
  NAND2_X1 U975 ( .A1(G112), .A2(n891), .ZN(n872) );
  NAND2_X1 U976 ( .A1(n873), .A2(n872), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(G162) );
  XOR2_X1 U978 ( .A(KEYINPUT48), .B(KEYINPUT112), .Z(n877) );
  XNOR2_X1 U979 ( .A(G164), .B(KEYINPUT46), .ZN(n876) );
  XNOR2_X1 U980 ( .A(n877), .B(n876), .ZN(n878) );
  XNOR2_X1 U981 ( .A(G162), .B(n878), .ZN(n888) );
  NAND2_X1 U982 ( .A1(G103), .A2(n898), .ZN(n880) );
  NAND2_X1 U983 ( .A1(G139), .A2(n896), .ZN(n879) );
  NAND2_X1 U984 ( .A1(n880), .A2(n879), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G115), .A2(n891), .ZN(n882) );
  NAND2_X1 U986 ( .A1(G127), .A2(n517), .ZN(n881) );
  NAND2_X1 U987 ( .A1(n882), .A2(n881), .ZN(n883) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n883), .Z(n884) );
  NOR2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n1003) );
  XNOR2_X1 U990 ( .A(n886), .B(n1003), .ZN(n887) );
  XNOR2_X1 U991 ( .A(n888), .B(n887), .ZN(n889) );
  XOR2_X1 U992 ( .A(G160), .B(n889), .Z(n890) );
  XNOR2_X1 U993 ( .A(n1012), .B(n890), .ZN(n905) );
  NAND2_X1 U994 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U995 ( .A1(G130), .A2(n517), .ZN(n893) );
  NAND2_X1 U996 ( .A1(n894), .A2(n893), .ZN(n895) );
  XNOR2_X1 U997 ( .A(KEYINPUT110), .B(n895), .ZN(n903) );
  NAND2_X1 U998 ( .A1(n896), .A2(G142), .ZN(n897) );
  XOR2_X1 U999 ( .A(KEYINPUT111), .B(n897), .Z(n900) );
  NAND2_X1 U1000 ( .A1(n898), .A2(G106), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1002 ( .A(n901), .B(KEYINPUT45), .Z(n902) );
  NOR2_X1 U1003 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1004 ( .A(n905), .B(n904), .Z(n909) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n910), .ZN(G395) );
  NOR2_X1 U1008 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1009 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1010 ( .A1(G397), .A2(n912), .ZN(n916) );
  NOR2_X1 U1011 ( .A1(G401), .A2(n917), .ZN(n913) );
  XNOR2_X1 U1012 ( .A(KEYINPUT113), .B(n913), .ZN(n914) );
  NOR2_X1 U1013 ( .A1(G395), .A2(n914), .ZN(n915) );
  NAND2_X1 U1014 ( .A1(n916), .A2(n915), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(n917), .ZN(G319) );
  XOR2_X1 U1017 ( .A(G1966), .B(G21), .Z(n920) );
  XNOR2_X1 U1018 ( .A(n918), .B(G5), .ZN(n919) );
  NAND2_X1 U1019 ( .A1(n920), .A2(n919), .ZN(n941) );
  XNOR2_X1 U1020 ( .A(G1348), .B(KEYINPUT59), .ZN(n921) );
  XNOR2_X1 U1021 ( .A(n921), .B(G4), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G1981), .B(G6), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G1341), .B(G19), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1026 ( .A(KEYINPUT121), .B(G1956), .Z(n926) );
  XNOR2_X1 U1027 ( .A(G20), .B(n926), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1029 ( .A(KEYINPUT122), .B(n929), .ZN(n930) );
  XNOR2_X1 U1030 ( .A(n930), .B(KEYINPUT60), .ZN(n939) );
  XOR2_X1 U1031 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n937) );
  XNOR2_X1 U1032 ( .A(G1986), .B(G24), .ZN(n932) );
  XNOR2_X1 U1033 ( .A(G22), .B(G1971), .ZN(n931) );
  NOR2_X1 U1034 ( .A1(n932), .A2(n931), .ZN(n935) );
  XNOR2_X1 U1035 ( .A(G1976), .B(KEYINPUT123), .ZN(n933) );
  XNOR2_X1 U1036 ( .A(n933), .B(G23), .ZN(n934) );
  NAND2_X1 U1037 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1038 ( .A(n937), .B(n936), .ZN(n938) );
  NAND2_X1 U1039 ( .A1(n939), .A2(n938), .ZN(n940) );
  NOR2_X1 U1040 ( .A1(n941), .A2(n940), .ZN(n942) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n942), .Z(n943) );
  NOR2_X1 U1042 ( .A1(G16), .A2(n943), .ZN(n944) );
  XOR2_X1 U1043 ( .A(KEYINPUT125), .B(n944), .Z(n998) );
  XNOR2_X1 U1044 ( .A(G1348), .B(n945), .ZN(n946) );
  NOR2_X1 U1045 ( .A1(n947), .A2(n946), .ZN(n949) );
  NAND2_X1 U1046 ( .A1(n949), .A2(n948), .ZN(n951) );
  XNOR2_X1 U1047 ( .A(G1961), .B(G301), .ZN(n950) );
  NOR2_X1 U1048 ( .A1(n951), .A2(n950), .ZN(n961) );
  XNOR2_X1 U1049 ( .A(n952), .B(G1341), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(G299), .B(G1956), .ZN(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n956) );
  NAND2_X1 U1052 ( .A1(G1971), .A2(G303), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(KEYINPUT120), .B(n957), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  NOR2_X1 U1057 ( .A1(n963), .A2(n962), .ZN(n968) );
  XNOR2_X1 U1058 ( .A(G1966), .B(G168), .ZN(n965) );
  NAND2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT57), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n971) );
  XOR2_X1 U1062 ( .A(G16), .B(KEYINPUT56), .Z(n969) );
  XNOR2_X1 U1063 ( .A(KEYINPUT119), .B(n969), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n996) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n972) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n972), .ZN(n988) );
  XNOR2_X1 U1067 ( .A(G2090), .B(G35), .ZN(n986) );
  XNOR2_X1 U1068 ( .A(G1991), .B(G25), .ZN(n974) );
  XNOR2_X1 U1069 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1070 ( .A1(n974), .A2(n973), .ZN(n980) );
  XOR2_X1 U1071 ( .A(G2067), .B(G26), .Z(n975) );
  NAND2_X1 U1072 ( .A1(n975), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(KEYINPUT116), .B(G1996), .ZN(n976) );
  XNOR2_X1 U1074 ( .A(G32), .B(n976), .ZN(n977) );
  NOR2_X1 U1075 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n983) );
  XOR2_X1 U1077 ( .A(G27), .B(n981), .Z(n982) );
  NOR2_X1 U1078 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1079 ( .A(KEYINPUT53), .B(n984), .ZN(n985) );
  NOR2_X1 U1080 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n989), .B(KEYINPUT117), .ZN(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT55), .B(n990), .ZN(n992) );
  INV_X1 U1084 ( .A(G29), .ZN(n991) );
  NAND2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1086 ( .A1(n993), .A2(G11), .ZN(n994) );
  XOR2_X1 U1087 ( .A(KEYINPUT118), .B(n994), .Z(n995) );
  NAND2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1089 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1090 ( .A(KEYINPUT126), .B(n999), .ZN(n1028) );
  XOR2_X1 U1091 ( .A(G2090), .B(G162), .Z(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XOR2_X1 U1093 ( .A(KEYINPUT51), .B(n1002), .Z(n1011) );
  XNOR2_X1 U1094 ( .A(G164), .B(G2078), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(G2072), .B(n1003), .Z(n1004) );
  XNOR2_X1 U1096 ( .A(KEYINPUT115), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(n1007), .B(KEYINPUT50), .ZN(n1009) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G160), .B(G2084), .ZN(n1013) );
  NAND2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XOR2_X1 U1104 ( .A(KEYINPUT114), .B(n1016), .Z(n1017) );
  NOR2_X1 U1105 ( .A1(n1018), .A2(n1017), .ZN(n1020) );
  NAND2_X1 U1106 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1107 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1108 ( .A(KEYINPUT52), .B(n1023), .ZN(n1025) );
  INV_X1 U1109 ( .A(KEYINPUT55), .ZN(n1024) );
  NAND2_X1 U1110 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(G29), .ZN(n1027) );
  NAND2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1029), .B(KEYINPUT62), .ZN(n1030) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1030), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

