//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 1 1 0 1 1 0 0 0 1 1 1 1 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:57 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT3), .B1(new_n188), .B2(G107), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n190));
  INV_X1    g004(.A(G107), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G104), .ZN(new_n192));
  INV_X1    g006(.A(G101), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n188), .A2(G107), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n189), .A2(new_n192), .A3(new_n193), .A4(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT76), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n191), .A2(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(new_n194), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n196), .B1(new_n198), .B2(G101), .ZN(new_n199));
  AOI211_X1 g013(.A(KEYINPUT76), .B(new_n193), .C1(new_n197), .C2(new_n194), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n195), .B1(new_n199), .B2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  OAI21_X1  g016(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n203));
  NOR2_X1   g017(.A1(new_n202), .A2(G146), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  OAI211_X1 g020(.A(G128), .B(new_n203), .C1(new_n204), .C2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n205), .A2(G143), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n202), .A2(G146), .ZN(new_n209));
  INV_X1    g023(.A(G128), .ZN(new_n210));
  OAI211_X1 g024(.A(new_n208), .B(new_n209), .C1(KEYINPUT1), .C2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n187), .B1(new_n201), .B2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT10), .ZN(new_n214));
  AND2_X1   g028(.A1(new_n207), .A2(new_n211), .ZN(new_n215));
  XNOR2_X1  g029(.A(G104), .B(G107), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT76), .B1(new_n216), .B2(new_n193), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n198), .A2(new_n196), .A3(G101), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n215), .A2(new_n219), .A3(KEYINPUT77), .A4(new_n195), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n213), .A2(new_n214), .A3(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n189), .A2(new_n192), .A3(new_n194), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(KEYINPUT4), .A3(new_n195), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n208), .A2(new_n209), .A3(KEYINPUT0), .A4(G128), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n204), .A2(new_n206), .ZN(new_n226));
  XNOR2_X1  g040(.A(KEYINPUT0), .B(G128), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT4), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n222), .A2(new_n230), .A3(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n224), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n215), .A2(new_n219), .A3(KEYINPUT10), .A4(new_n195), .ZN(new_n233));
  AND2_X1   g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  OR2_X1    g048(.A1(KEYINPUT65), .A2(G137), .ZN(new_n235));
  NAND2_X1  g049(.A1(KEYINPUT65), .A2(G137), .ZN(new_n236));
  AND2_X1   g050(.A1(KEYINPUT11), .A2(G134), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G137), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT11), .B1(new_n239), .B2(G134), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G134), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G137), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G131), .ZN(new_n245));
  AOI21_X1  g059(.A(G131), .B1(new_n242), .B2(G137), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n238), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n245), .A2(KEYINPUT78), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(KEYINPUT78), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n221), .A2(new_n234), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n201), .A2(new_n212), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n213), .A2(new_n220), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g067(.A1(KEYINPUT65), .A2(G137), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT65), .A2(G137), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n240), .B1(new_n256), .B2(new_n237), .ZN(new_n257));
  AOI22_X1  g071(.A1(G131), .A2(new_n244), .B1(new_n257), .B2(new_n246), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AND3_X1   g073(.A1(new_n253), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(KEYINPUT12), .B1(new_n253), .B2(new_n259), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n251), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(G110), .B(G140), .ZN(new_n263));
  INV_X1    g077(.A(G227), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n263), .B(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n251), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n258), .B1(new_n221), .B2(new_n234), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n262), .A2(new_n266), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI21_X1  g085(.A(G469), .B1(new_n271), .B2(G902), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT79), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT79), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n274), .B(G469), .C1(new_n271), .C2(G902), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n221), .A2(new_n234), .A3(new_n250), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n266), .B1(new_n276), .B2(new_n269), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT80), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT80), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n279), .B(new_n266), .C1(new_n276), .C2(new_n269), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n253), .A2(new_n259), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT12), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n253), .A2(KEYINPUT12), .A3(new_n259), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n268), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n280), .A3(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(G469), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n273), .A2(new_n275), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  INV_X1    g106(.A(G119), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(G116), .ZN(new_n294));
  INV_X1    g108(.A(G116), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G119), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g111(.A(KEYINPUT2), .B(G113), .ZN(new_n298));
  OAI21_X1  g112(.A(new_n292), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  XNOR2_X1  g113(.A(G116), .B(G119), .ZN(new_n300));
  INV_X1    g114(.A(G113), .ZN(new_n301));
  AND2_X1   g115(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(KEYINPUT2), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n300), .B(KEYINPUT67), .C1(new_n302), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT66), .B1(new_n294), .B2(new_n296), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n300), .A2(KEYINPUT66), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n307), .A2(new_n308), .A3(new_n298), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n305), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(new_n224), .A3(new_n231), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n294), .A2(new_n296), .A3(KEYINPUT66), .ZN(new_n312));
  OAI21_X1  g126(.A(KEYINPUT5), .B1(new_n312), .B2(new_n306), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT81), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n314), .B1(new_n294), .B2(KEYINPUT5), .ZN(new_n315));
  INV_X1    g129(.A(KEYINPUT5), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n316), .A2(new_n293), .A3(KEYINPUT81), .A4(G116), .ZN(new_n317));
  AND3_X1   g131(.A1(new_n315), .A2(G113), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  AND3_X1   g133(.A1(new_n189), .A2(new_n192), .A3(new_n194), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n217), .A2(new_n218), .B1(new_n320), .B2(new_n193), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n321), .A3(new_n305), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n311), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT82), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT6), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n311), .A2(new_n322), .A3(KEYINPUT82), .ZN(new_n327));
  XNOR2_X1  g141(.A(G110), .B(G122), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n325), .A2(new_n326), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n225), .B(G125), .C1(new_n226), .C2(new_n227), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n331), .B1(new_n212), .B2(G125), .ZN(new_n332));
  INV_X1    g146(.A(G224), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G953), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n332), .B(new_n334), .Z(new_n335));
  AND3_X1   g149(.A1(new_n311), .A2(new_n322), .A3(KEYINPUT82), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT82), .B1(new_n311), .B2(new_n322), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n336), .A2(new_n337), .A3(new_n328), .ZN(new_n338));
  OAI21_X1  g152(.A(KEYINPUT6), .B1(new_n323), .B2(new_n329), .ZN(new_n339));
  OAI211_X1 g153(.A(new_n330), .B(new_n335), .C1(new_n338), .C2(new_n339), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n311), .A2(new_n322), .A3(new_n328), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n294), .A2(new_n296), .A3(KEYINPUT5), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n315), .A2(new_n342), .A3(G113), .A4(new_n317), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n305), .A2(new_n219), .A3(new_n195), .A4(new_n343), .ZN(new_n344));
  AOI22_X1  g158(.A1(new_n313), .A2(new_n318), .B1(new_n299), .B2(new_n304), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(new_n321), .ZN(new_n346));
  XOR2_X1   g160(.A(new_n328), .B(KEYINPUT8), .Z(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT7), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n332), .B1(new_n349), .B2(new_n334), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n334), .A2(new_n349), .ZN(new_n351));
  OAI211_X1 g165(.A(new_n331), .B(new_n351), .C1(new_n212), .C2(G125), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n346), .A2(new_n348), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT83), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n341), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n319), .A2(new_n305), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n356), .A2(new_n201), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n347), .B1(new_n357), .B2(new_n344), .ZN(new_n358));
  AND2_X1   g172(.A1(new_n350), .A2(new_n352), .ZN(new_n359));
  OAI21_X1  g173(.A(KEYINPUT83), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(G902), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n340), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(G210), .B1(G237), .B2(G902), .ZN(new_n363));
  XOR2_X1   g177(.A(new_n363), .B(KEYINPUT84), .Z(new_n364));
  NAND2_X1  g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n340), .A2(new_n361), .A3(new_n363), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G221), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT9), .B(G234), .ZN(new_n369));
  XNOR2_X1  g183(.A(new_n369), .B(KEYINPUT75), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n368), .B1(new_n370), .B2(new_n289), .ZN(new_n371));
  OAI21_X1  g185(.A(G214), .B1(G237), .B2(G902), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g188(.A1(new_n291), .A2(new_n367), .A3(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(G113), .B(G122), .ZN(new_n376));
  XNOR2_X1  g190(.A(new_n376), .B(new_n188), .ZN(new_n377));
  INV_X1    g191(.A(G140), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G125), .ZN(new_n379));
  INV_X1    g193(.A(G125), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G140), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n382), .B(new_n205), .ZN(new_n383));
  INV_X1    g197(.A(G237), .ZN(new_n384));
  INV_X1    g198(.A(G953), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G214), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n202), .ZN(new_n387));
  NOR2_X1   g201(.A1(G237), .A2(G953), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(G143), .A3(G214), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT18), .A3(G131), .ZN(new_n391));
  NAND2_X1  g205(.A1(KEYINPUT18), .A2(G131), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(new_n389), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n383), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT87), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT17), .ZN(new_n396));
  AND4_X1   g210(.A1(G143), .A2(new_n384), .A3(new_n385), .A4(G214), .ZN(new_n397));
  AOI21_X1  g211(.A(G143), .B1(new_n388), .B2(G214), .ZN(new_n398));
  OAI21_X1  g212(.A(G131), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT85), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT85), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n401), .A3(G131), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n396), .B1(new_n400), .B2(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT16), .ZN(new_n404));
  OR3_X1    g218(.A1(new_n380), .A2(KEYINPUT16), .A3(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n205), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n404), .A2(new_n405), .A3(G146), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n395), .B1(new_n403), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n401), .B1(new_n390), .B2(G131), .ZN(new_n411));
  INV_X1    g225(.A(G131), .ZN(new_n412));
  AOI211_X1 g226(.A(KEYINPUT85), .B(new_n412), .C1(new_n387), .C2(new_n389), .ZN(new_n413));
  OAI21_X1  g227(.A(KEYINPUT17), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n409), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(KEYINPUT87), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n411), .A2(new_n413), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT88), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n387), .A2(new_n412), .A3(new_n389), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n418), .A2(new_n419), .A3(new_n396), .A4(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n400), .A2(new_n402), .A3(new_n396), .A4(new_n420), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT88), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n421), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n377), .B(new_n394), .C1(new_n417), .C2(new_n424), .ZN(new_n425));
  AND3_X1   g239(.A1(new_n400), .A2(new_n402), .A3(new_n420), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT73), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n408), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n404), .A2(new_n405), .A3(KEYINPUT73), .A4(G146), .ZN(new_n429));
  AND3_X1   g243(.A1(new_n379), .A2(new_n381), .A3(KEYINPUT19), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT19), .B1(new_n379), .B2(new_n381), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n428), .B(new_n429), .C1(G146), .C2(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n394), .B1(new_n426), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(KEYINPUT86), .ZN(new_n435));
  INV_X1    g249(.A(new_n377), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT86), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n437), .B(new_n394), .C1(new_n426), .C2(new_n433), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  NOR2_X1   g255(.A1(G475), .A2(G902), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(KEYINPUT89), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT89), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n425), .A2(new_n439), .A3(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n445), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n444), .B1(new_n448), .B2(KEYINPUT20), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n394), .B1(new_n417), .B2(new_n424), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n436), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(new_n425), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n289), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n453), .A2(G475), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n385), .A2(G952), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(G234), .B2(G237), .ZN(new_n456));
  NAND2_X1  g270(.A1(G234), .A2(G237), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n457), .A2(G902), .A3(G953), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(KEYINPUT21), .B(G898), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(G122), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(G116), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n295), .A2(G122), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G107), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n191), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT90), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n210), .A2(G143), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT13), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n242), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g287(.A(G128), .B(G143), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n473), .B(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n466), .A2(new_n467), .A3(KEYINPUT90), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n470), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n295), .A2(KEYINPUT14), .A3(G122), .ZN(new_n478));
  OAI211_X1 g292(.A(G107), .B(new_n478), .C1(new_n465), .C2(KEYINPUT14), .ZN(new_n479));
  OR2_X1    g293(.A1(new_n474), .A2(G134), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n474), .A2(G134), .ZN(new_n481));
  NAND4_X1  g295(.A1(new_n479), .A2(new_n480), .A3(new_n467), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n370), .A2(G217), .A3(new_n385), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n484), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n486), .A2(new_n477), .A3(new_n482), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n485), .A2(KEYINPUT91), .A3(new_n487), .ZN(new_n488));
  OR3_X1    g302(.A1(new_n483), .A2(KEYINPUT91), .A3(new_n484), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(new_n489), .A3(new_n289), .ZN(new_n490));
  INV_X1    g304(.A(G478), .ZN(new_n491));
  NOR2_X1   g305(.A1(new_n491), .A2(KEYINPUT15), .ZN(new_n492));
  OR2_X1    g306(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n490), .A2(new_n492), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR4_X1   g309(.A1(new_n449), .A2(new_n454), .A3(new_n461), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n375), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT25), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n293), .A2(G128), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n210), .A2(KEYINPUT23), .A3(G119), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n293), .A2(G128), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n499), .B(new_n500), .C1(new_n501), .C2(KEYINPUT23), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  XNOR2_X1  g317(.A(G119), .B(G128), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n502), .A2(G110), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n409), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT72), .B(G110), .ZN(new_n507));
  OAI22_X1  g321(.A1(new_n502), .A2(new_n507), .B1(new_n503), .B2(new_n504), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n382), .A2(new_n205), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n428), .A2(new_n508), .A3(new_n429), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  AND3_X1   g326(.A1(new_n385), .A2(G221), .A3(G234), .ZN(new_n513));
  XOR2_X1   g327(.A(new_n512), .B(new_n513), .Z(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n506), .A2(new_n510), .A3(new_n514), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n498), .B1(new_n518), .B2(G902), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n516), .A2(KEYINPUT25), .A3(new_n289), .A4(new_n517), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n519), .A2(KEYINPUT74), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(G217), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(G234), .B2(new_n289), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n519), .B2(KEYINPUT74), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  NOR3_X1   g339(.A1(new_n518), .A2(G902), .A3(new_n523), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(G472), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n312), .A2(new_n306), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n530), .A2(new_n298), .B1(new_n299), .B2(new_n304), .ZN(new_n531));
  AOI21_X1  g345(.A(G134), .B1(new_n235), .B2(new_n236), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n239), .A2(G134), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G131), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n535), .A2(new_n247), .A3(new_n211), .A4(new_n207), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n258), .B2(new_n228), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n531), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT68), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT30), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n238), .A2(new_n241), .A3(new_n246), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n242), .B1(new_n254), .B2(new_n255), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n412), .B1(new_n543), .B2(new_n533), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n541), .B1(new_n545), .B2(new_n215), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n412), .B1(new_n257), .B2(new_n243), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n229), .B1(new_n547), .B2(new_n542), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n540), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(KEYINPUT65), .B(G137), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n534), .B1(new_n550), .B2(new_n242), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n247), .B1(new_n551), .B2(new_n412), .ZN(new_n552));
  OAI21_X1  g366(.A(KEYINPUT30), .B1(new_n552), .B2(new_n212), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n228), .B1(new_n245), .B2(new_n247), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT68), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n539), .B1(new_n549), .B2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT31), .ZN(new_n557));
  INV_X1    g371(.A(new_n536), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n558), .A2(new_n554), .A3(new_n310), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n388), .A2(G210), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT27), .ZN(new_n561));
  XNOR2_X1  g375(.A(KEYINPUT26), .B(G101), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n559), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n556), .A2(new_n557), .A3(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT28), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n310), .B1(new_n558), .B2(new_n554), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n531), .B(new_n536), .C1(new_n258), .C2(new_n228), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n569), .A2(new_n567), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n564), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n557), .B1(new_n556), .B2(new_n565), .ZN(new_n574));
  OAI211_X1 g388(.A(new_n529), .B(new_n289), .C1(new_n573), .C2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT32), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g391(.A1(new_n576), .A2(G472), .A3(G902), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n578), .B1(new_n573), .B2(new_n574), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  OAI211_X1 g395(.A(KEYINPUT71), .B(new_n578), .C1(new_n573), .C2(new_n574), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(KEYINPUT70), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n563), .A2(KEYINPUT29), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n570), .A2(new_n571), .A3(new_n585), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n584), .B1(new_n586), .B2(G902), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n531), .B1(new_n548), .B2(new_n536), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT28), .B1(new_n559), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n569), .A2(new_n567), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  OAI211_X1 g405(.A(KEYINPUT70), .B(new_n289), .C1(new_n591), .C2(new_n585), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n589), .A2(new_n563), .A3(new_n590), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT29), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n546), .A2(new_n540), .A3(new_n548), .ZN(new_n595));
  OAI21_X1  g409(.A(KEYINPUT68), .B1(new_n553), .B2(new_n554), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n559), .B1(new_n597), .B2(new_n539), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n593), .B(new_n594), .C1(new_n563), .C2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT69), .ZN(new_n600));
  OAI211_X1 g414(.A(new_n587), .B(new_n592), .C1(new_n599), .C2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n570), .A2(new_n571), .ZN(new_n602));
  AOI21_X1  g416(.A(KEYINPUT29), .B1(new_n602), .B2(new_n563), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n556), .A2(new_n569), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n604), .A2(new_n564), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT69), .B1(new_n603), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(G472), .B1(new_n601), .B2(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n528), .B1(new_n583), .B2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n497), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n193), .ZN(G3));
  AOI22_X1  g425(.A1(new_n277), .A2(KEYINPUT80), .B1(new_n285), .B2(new_n268), .ZN(new_n612));
  AOI21_X1  g426(.A(G902), .B1(new_n612), .B2(new_n280), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n288), .A2(new_n613), .B1(new_n272), .B2(KEYINPUT79), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n371), .B1(new_n614), .B2(new_n275), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n556), .A2(new_n565), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT31), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n617), .A2(new_n566), .A3(new_n572), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n289), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n619), .A2(G472), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n575), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n528), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n449), .A2(new_n454), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT94), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n487), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n485), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n483), .A2(new_n625), .A3(new_n484), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(KEYINPUT33), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(KEYINPUT95), .ZN(new_n630));
  INV_X1    g444(.A(KEYINPUT95), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n627), .A2(new_n631), .A3(KEYINPUT33), .A4(new_n628), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT92), .B(KEYINPUT33), .Z(new_n634));
  NAND3_X1  g448(.A1(new_n488), .A2(new_n489), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT93), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n488), .A2(new_n489), .A3(KEYINPUT93), .A4(new_n634), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n491), .A2(G902), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n633), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n490), .A2(new_n491), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n642), .A2(KEYINPUT96), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n490), .A2(new_n644), .A3(new_n491), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n641), .A2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  INV_X1    g462(.A(new_n461), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n340), .A2(new_n361), .A3(new_n363), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n363), .B1(new_n340), .B2(new_n361), .ZN(new_n651));
  OAI211_X1 g465(.A(new_n649), .B(new_n372), .C1(new_n650), .C2(new_n651), .ZN(new_n652));
  NOR3_X1   g466(.A1(new_n624), .A2(new_n648), .A3(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n623), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  NAND2_X1  g470(.A1(new_n453), .A2(G475), .ZN(new_n657));
  AND3_X1   g471(.A1(new_n425), .A2(new_n446), .A3(new_n439), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n446), .B1(new_n425), .B2(new_n439), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n441), .B1(new_n660), .B2(new_n442), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n657), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n461), .B(KEYINPUT97), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n665), .B1(new_n493), .B2(new_n494), .ZN(new_n666));
  OAI211_X1 g480(.A(new_n666), .B(new_n372), .C1(new_n650), .C2(new_n651), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n663), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n623), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g483(.A(KEYINPUT35), .B(G107), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n669), .B(new_n670), .ZN(G9));
  NOR2_X1   g485(.A1(new_n515), .A2(KEYINPUT36), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n511), .B(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n523), .A2(G902), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n521), .B2(new_n524), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n620), .A2(new_n575), .A3(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n497), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(KEYINPUT37), .B(G110), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  NOR2_X1   g494(.A1(new_n650), .A2(new_n651), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n291), .A2(new_n374), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n660), .A2(new_n441), .A3(new_n442), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n456), .B(KEYINPUT98), .Z(new_n687));
  INV_X1    g501(.A(new_n687), .ZN(new_n688));
  INV_X1    g502(.A(G900), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n688), .B1(new_n689), .B2(new_n459), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n657), .A2(new_n686), .A3(new_n495), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n676), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n693), .B1(new_n583), .B2(new_n607), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n683), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G128), .ZN(G30));
  NAND3_X1  g510(.A1(new_n577), .A2(new_n581), .A3(new_n582), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT101), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n564), .B1(new_n559), .B2(new_n588), .ZN(new_n699));
  OR2_X1    g513(.A1(new_n699), .A2(KEYINPUT100), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(KEYINPUT100), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n700), .A2(G472), .A3(new_n616), .A4(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(G472), .A2(G902), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n698), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  AND3_X1   g518(.A1(new_n702), .A2(new_n698), .A3(new_n703), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n697), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n367), .B(new_n707), .Z(new_n708));
  XOR2_X1   g522(.A(new_n690), .B(KEYINPUT39), .Z(new_n709));
  NAND2_X1  g523(.A1(new_n615), .A2(new_n709), .ZN(new_n710));
  AOI211_X1 g524(.A(new_n706), .B(new_n708), .C1(new_n710), .C2(KEYINPUT40), .ZN(new_n711));
  OAI211_X1 g525(.A(new_n495), .B(new_n372), .C1(new_n449), .C2(new_n454), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n676), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT102), .ZN(new_n714));
  OAI211_X1 g528(.A(new_n711), .B(new_n714), .C1(KEYINPUT40), .C2(new_n710), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  OAI211_X1 g530(.A(new_n647), .B(new_n691), .C1(new_n449), .C2(new_n454), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n683), .A2(new_n694), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT103), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n601), .ZN(new_n722));
  INV_X1    g536(.A(new_n606), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n529), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n676), .B1(new_n724), .B2(new_n697), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n291), .A2(new_n374), .A3(new_n682), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(KEYINPUT103), .A3(new_n718), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n721), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G146), .ZN(G48));
  INV_X1    g544(.A(new_n582), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT71), .B1(new_n618), .B2(new_n578), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n607), .A3(new_n577), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n288), .B1(new_n287), .B2(new_n289), .ZN(new_n736));
  NOR3_X1   g550(.A1(new_n735), .A2(new_n736), .A3(new_n371), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n734), .A2(new_n527), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n685), .A2(new_n443), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n657), .ZN(new_n740));
  INV_X1    g554(.A(new_n652), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n647), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT104), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n653), .A2(new_n608), .A3(new_n744), .A4(new_n737), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT41), .B(G113), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n746), .B(new_n747), .ZN(G15));
  NAND3_X1  g562(.A1(new_n608), .A2(new_n668), .A3(new_n737), .ZN(new_n749));
  XNOR2_X1  g563(.A(KEYINPUT105), .B(G116), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n749), .B(new_n750), .ZN(G18));
  NAND2_X1  g565(.A1(new_n287), .A2(new_n289), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(G469), .ZN(new_n753));
  INV_X1    g567(.A(new_n371), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n753), .A2(new_n754), .A3(new_n290), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n372), .B1(new_n650), .B2(new_n651), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n694), .A2(new_n757), .A3(new_n496), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  NOR3_X1   g573(.A1(new_n621), .A2(new_n528), .A3(new_n665), .ZN(new_n760));
  AOI22_X1  g574(.A1(new_n739), .A2(new_n657), .B1(new_n494), .B2(new_n493), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n757), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G122), .ZN(G24));
  NOR2_X1   g577(.A1(new_n717), .A2(new_n677), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n757), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT106), .B(G125), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G27));
  NAND3_X1  g581(.A1(new_n365), .A2(new_n366), .A3(new_n372), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT108), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n365), .A2(KEYINPUT108), .A3(new_n366), .A4(new_n372), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(new_n754), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT107), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n290), .A2(new_n773), .A3(new_n272), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n773), .B1(new_n290), .B2(new_n272), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n577), .A2(new_n579), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n528), .B1(new_n780), .B2(new_n607), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n718), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT42), .B1(new_n778), .B2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n770), .A2(new_n754), .A3(new_n771), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n290), .A2(new_n272), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n785), .A2(KEYINPUT107), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n786), .A2(new_n774), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n784), .A2(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n717), .A2(KEYINPUT42), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n608), .A3(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n783), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(new_n412), .ZN(G33));
  NAND4_X1  g606(.A1(new_n772), .A2(new_n608), .A3(new_n692), .A4(new_n777), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G134), .ZN(G36));
  NOR2_X1   g608(.A1(new_n271), .A2(KEYINPUT45), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n795), .A2(new_n288), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n271), .A2(KEYINPUT45), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(G469), .A2(G902), .ZN(new_n799));
  AOI21_X1  g613(.A(KEYINPUT46), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n735), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n798), .A2(KEYINPUT46), .A3(new_n799), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n371), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(new_n709), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n770), .A2(new_n771), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT43), .B1(new_n740), .B2(new_n648), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n624), .A2(new_n808), .A3(new_n647), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n807), .A2(new_n621), .A3(new_n676), .A4(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT44), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n811), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n804), .A2(new_n806), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  OR2_X1    g629(.A1(new_n803), .A2(KEYINPUT47), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n803), .A2(KEYINPUT47), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n805), .A2(new_n734), .A3(new_n527), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n718), .A3(new_n819), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(G140), .ZN(G42));
  INV_X1    g635(.A(KEYINPUT53), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n712), .A2(new_n681), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n371), .B1(new_n691), .B2(KEYINPUT111), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n693), .B(new_n824), .C1(KEYINPUT111), .C2(new_n691), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n705), .A2(new_n704), .ZN(new_n826));
  AOI21_X1  g640(.A(new_n825), .B1(new_n583), .B2(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n823), .A2(new_n827), .A3(new_n777), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n695), .A2(new_n828), .A3(new_n765), .ZN(new_n829));
  AND3_X1   g643(.A1(new_n729), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT52), .B1(new_n729), .B2(new_n829), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT109), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n743), .A2(new_n745), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n749), .A2(new_n758), .A3(new_n762), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT110), .ZN(new_n837));
  XNOR2_X1  g651(.A(new_n495), .B(new_n837), .ZN(new_n838));
  AND3_X1   g652(.A1(new_n770), .A2(new_n771), .A3(new_n838), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n686), .A2(new_n657), .A3(new_n691), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n694), .A3(new_n615), .A4(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n772), .A2(new_n764), .A3(new_n777), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n793), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT42), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n527), .B1(new_n724), .B2(new_n779), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n717), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n844), .B1(new_n846), .B2(new_n788), .ZN(new_n847));
  AND4_X1   g661(.A1(new_n608), .A2(new_n772), .A3(new_n789), .A4(new_n777), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n843), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n749), .A2(new_n758), .A3(new_n762), .ZN(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(KEYINPUT109), .A3(new_n746), .ZN(new_n851));
  INV_X1    g665(.A(new_n677), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n375), .B(new_n496), .C1(new_n608), .C2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n624), .A2(new_n648), .ZN(new_n854));
  INV_X1    g668(.A(new_n838), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n854), .B1(new_n624), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n375), .A2(new_n760), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n836), .A2(new_n849), .A3(new_n851), .A4(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n822), .B1(new_n832), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT113), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT103), .B1(new_n727), .B2(new_n718), .ZN(new_n864));
  NOR4_X1   g678(.A1(new_n725), .A2(new_n726), .A3(new_n720), .A4(new_n717), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n695), .A2(new_n828), .A3(new_n765), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n863), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n729), .A2(new_n829), .A3(KEYINPUT52), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n850), .A2(KEYINPUT109), .A3(new_n746), .ZN(new_n871));
  AOI21_X1  g685(.A(KEYINPUT109), .B1(new_n850), .B2(new_n746), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n791), .A2(new_n858), .A3(new_n843), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n870), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT113), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n876), .A3(new_n822), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT54), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n822), .B1(new_n868), .B2(new_n869), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n879), .A2(new_n746), .A3(new_n850), .A4(new_n874), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n862), .A2(new_n877), .A3(new_n878), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n870), .A2(new_n873), .A3(KEYINPUT53), .A4(new_n874), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n861), .A2(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT112), .B1(new_n883), .B2(KEYINPUT54), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT112), .ZN(new_n885));
  AOI211_X1 g699(.A(new_n885), .B(new_n878), .C1(new_n861), .C2(new_n882), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n881), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(KEYINPUT114), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT114), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n889), .B(new_n881), .C1(new_n884), .C2(new_n886), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n807), .A2(new_n688), .A3(new_n809), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT115), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n891), .A2(new_n892), .ZN(new_n894));
  AOI211_X1 g708(.A(new_n755), .B(new_n805), .C1(new_n893), .C2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n805), .A2(new_n755), .ZN(new_n896));
  AND4_X1   g710(.A1(new_n527), .A2(new_n896), .A3(new_n456), .A4(new_n706), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n740), .A2(new_n647), .ZN(new_n898));
  AOI22_X1  g712(.A1(new_n895), .A2(new_n852), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n622), .ZN(new_n900));
  AOI21_X1  g714(.A(new_n900), .B1(new_n893), .B2(new_n894), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n708), .A2(new_n373), .A3(new_n737), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT50), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT50), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n899), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(KEYINPUT51), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n901), .A2(new_n806), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n753), .A2(new_n371), .A3(new_n290), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n816), .A2(new_n817), .A3(new_n910), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n909), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(KEYINPUT117), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n905), .A2(new_n906), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT117), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n915), .A2(new_n916), .A3(new_n899), .A4(new_n912), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n901), .A2(new_n757), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT118), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n455), .B1(new_n897), .B2(new_n854), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n919), .A2(new_n920), .A3(new_n921), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n920), .B1(new_n919), .B2(new_n921), .ZN(new_n923));
  XOR2_X1   g737(.A(KEYINPUT119), .B(KEYINPUT48), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n895), .A2(new_n781), .A3(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n925), .B1(new_n895), .B2(new_n781), .ZN(new_n927));
  OAI22_X1  g741(.A1(new_n922), .A2(new_n923), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n816), .A2(KEYINPUT116), .A3(new_n817), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(new_n910), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT116), .B1(new_n816), .B2(new_n817), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n909), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OAI211_X1 g746(.A(new_n932), .B(new_n899), .C1(new_n906), .C2(new_n905), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n933), .B2(new_n908), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n918), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n888), .A2(new_n890), .A3(new_n935), .ZN(new_n936));
  OR2_X1    g750(.A1(G952), .A2(G953), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  AND4_X1   g752(.A1(new_n527), .A2(new_n706), .A3(new_n624), .A4(new_n647), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n708), .A2(new_n374), .ZN(new_n940));
  OAI21_X1  g754(.A(KEYINPUT49), .B1(new_n735), .B2(new_n736), .ZN(new_n941));
  OR3_X1    g755(.A1(new_n735), .A2(new_n736), .A3(KEYINPUT49), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n938), .A2(new_n943), .ZN(G75));
  OAI21_X1  g758(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n335), .ZN(new_n946));
  XOR2_X1   g760(.A(KEYINPUT120), .B(KEYINPUT55), .Z(new_n947));
  XNOR2_X1  g761(.A(new_n946), .B(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n862), .A2(new_n877), .A3(new_n880), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n949), .A2(G902), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(G210), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT56), .ZN(new_n952));
  AOI21_X1  g766(.A(new_n948), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n948), .A2(new_n952), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n954), .B1(new_n950), .B2(new_n364), .ZN(new_n955));
  NOR2_X1   g769(.A1(new_n385), .A2(G952), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n953), .A2(new_n955), .A3(new_n956), .ZN(G51));
  INV_X1    g771(.A(new_n798), .ZN(new_n958));
  AOI21_X1  g772(.A(KEYINPUT121), .B1(new_n950), .B2(new_n958), .ZN(new_n959));
  AND4_X1   g773(.A1(KEYINPUT121), .A2(new_n949), .A3(G902), .A4(new_n958), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n799), .B(KEYINPUT57), .Z(new_n962));
  AND2_X1   g776(.A1(new_n949), .A2(KEYINPUT54), .ZN(new_n963));
  INV_X1    g777(.A(new_n881), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(new_n287), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n956), .B1(new_n961), .B2(new_n966), .ZN(G54));
  NAND3_X1  g781(.A1(new_n950), .A2(KEYINPUT58), .A3(G475), .ZN(new_n968));
  INV_X1    g782(.A(new_n660), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n956), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n968), .A2(new_n969), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G60));
  AND2_X1   g788(.A1(new_n633), .A2(new_n639), .ZN(new_n975));
  NAND2_X1  g789(.A1(G478), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT59), .Z(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI211_X1 g792(.A(new_n975), .B(new_n978), .C1(new_n963), .C2(new_n964), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n971), .ZN(new_n980));
  INV_X1    g794(.A(new_n890), .ZN(new_n981));
  INV_X1    g795(.A(new_n860), .ZN(new_n982));
  AOI22_X1  g796(.A1(new_n875), .A2(new_n822), .B1(new_n982), .B2(new_n879), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n885), .B1(new_n983), .B2(new_n878), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n883), .A2(KEYINPUT112), .A3(KEYINPUT54), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n889), .B1(new_n986), .B2(new_n881), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n978), .B1(new_n981), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n975), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n980), .B1(new_n988), .B2(new_n989), .ZN(G63));
  NAND2_X1  g804(.A1(G217), .A2(G902), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(KEYINPUT122), .ZN(new_n992));
  XNOR2_X1  g806(.A(new_n992), .B(KEYINPUT60), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n949), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n994), .A2(new_n518), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n949), .A2(new_n673), .A3(new_n993), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n995), .A2(new_n971), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT61), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(G66));
  OAI21_X1  g813(.A(G953), .B1(new_n460), .B2(new_n333), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n873), .A2(new_n859), .ZN(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n1000), .B1(new_n1002), .B2(G953), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n945), .B1(G898), .B2(new_n385), .ZN(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(KEYINPUT124), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  XNOR2_X1  g820(.A(new_n1003), .B(new_n1006), .ZN(G69));
  NAND2_X1  g821(.A1(new_n537), .A2(new_n538), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n597), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1009), .B(new_n432), .ZN(new_n1010));
  OR4_X1    g824(.A1(new_n609), .A2(new_n856), .A3(new_n710), .A4(new_n805), .ZN(new_n1011));
  NAND3_X1  g825(.A1(new_n820), .A2(new_n814), .A3(new_n1011), .ZN(new_n1012));
  AND3_X1   g826(.A1(new_n729), .A2(new_n695), .A3(new_n765), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1013), .A2(new_n715), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1012), .B1(KEYINPUT62), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1015), .B1(KEYINPUT62), .B2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1010), .B1(new_n1016), .B2(new_n385), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n804), .A2(new_n781), .A3(new_n823), .ZN(new_n1018));
  AND4_X1   g832(.A1(new_n783), .A2(new_n1018), .A3(new_n790), .A4(new_n793), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n1019), .A2(new_n814), .A3(new_n820), .A4(new_n1013), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n1020), .A2(G953), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1010), .B1(new_n689), .B2(new_n385), .ZN(new_n1022));
  OAI21_X1  g836(.A(KEYINPUT125), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1017), .A2(new_n1023), .ZN(new_n1024));
  OAI21_X1  g838(.A(G953), .B1(new_n264), .B2(new_n689), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(G72));
  XNOR2_X1  g840(.A(new_n703), .B(KEYINPUT63), .ZN(new_n1027));
  INV_X1    g841(.A(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n1020), .B2(new_n1001), .ZN(new_n1029));
  INV_X1    g843(.A(KEYINPUT126), .ZN(new_n1030));
  AOI211_X1 g844(.A(new_n563), .B(new_n604), .C1(new_n1029), .C2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g845(.A(new_n1031), .B1(new_n1030), .B2(new_n1029), .ZN(new_n1032));
  OAI21_X1  g846(.A(new_n1028), .B1(new_n1016), .B2(new_n1001), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1033), .A2(new_n563), .A3(new_n604), .ZN(new_n1034));
  AOI21_X1  g848(.A(new_n1027), .B1(new_n605), .B2(new_n616), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n956), .B1(new_n883), .B2(new_n1035), .ZN(new_n1036));
  AND3_X1   g850(.A1(new_n1032), .A2(new_n1034), .A3(new_n1036), .ZN(G57));
endmodule


