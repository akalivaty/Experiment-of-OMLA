//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 0 1 0 1 0 1 1 0 0 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 1 1 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n202, new_n203, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286, new_n1287,
    new_n1288, new_n1289, new_n1290;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  INV_X1    g0001(.A(G97), .ZN(new_n202));
  INV_X1    g0002(.A(G107), .ZN(new_n203));
  NAND2_X1  g0003(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n204), .A2(G87), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G355));
  INV_X1    g0006(.A(G77), .ZN(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  INV_X1    g0010(.A(G68), .ZN(new_n211));
  INV_X1    g0011(.A(G238), .ZN(new_n212));
  INV_X1    g0012(.A(G264), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n203), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n209), .B(new_n214), .C1(G116), .C2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G20), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  XOR2_X1   g0022(.A(new_n222), .B(KEYINPUT1), .Z(new_n223));
  NOR2_X1   g0023(.A1(new_n221), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND3_X1  g0026(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n227));
  OAI21_X1  g0027(.A(G50), .B1(G58), .B2(G68), .ZN(new_n228));
  XOR2_X1   g0028(.A(new_n228), .B(KEYINPUT65), .Z(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n223), .B(new_n226), .C1(new_n227), .C2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT68), .ZN(new_n234));
  XOR2_X1   g0034(.A(G226), .B(G232), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(G250), .B(G257), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(new_n213), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n238), .B(new_n241), .ZN(G358));
  XOR2_X1   g0042(.A(G50), .B(G58), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT69), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G68), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G87), .B(G97), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n247), .B(KEYINPUT70), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n246), .B(new_n250), .Z(G351));
  INV_X1    g0051(.A(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT3), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1698), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G222), .ZN(new_n259));
  INV_X1    g0059(.A(G223), .ZN(new_n260));
  OAI211_X1 g0060(.A(new_n257), .B(new_n259), .C1(new_n260), .C2(new_n258), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G41), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n262), .A2(G1), .A3(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n261), .B(new_n264), .C1(G77), .C2(new_n257), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n263), .A2(new_n267), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n265), .B(new_n270), .C1(new_n217), .C2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G169), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n274), .B1(G179), .B2(new_n272), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n276), .A2(G50), .ZN(new_n277));
  NAND3_X1  g0077(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(G1), .A2(G13), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  XNOR2_X1  g0081(.A(KEYINPUT8), .B(G58), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(KEYINPUT71), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT71), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n284), .A2(new_n218), .A3(KEYINPUT8), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n252), .A2(G20), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G20), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G58), .A2(G68), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n289), .B1(new_n290), .B2(new_n216), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n291), .B1(G150), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n281), .B1(new_n288), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n266), .A2(G20), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n281), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  AOI211_X1 g0097(.A(new_n277), .B(new_n294), .C1(G50), .C2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n275), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n272), .A2(G200), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(KEYINPUT74), .ZN(new_n302));
  INV_X1    g0102(.A(G190), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n272), .A2(new_n303), .ZN(new_n304));
  OAI211_X1 g0104(.A(new_n301), .B(new_n304), .C1(new_n298), .C2(KEYINPUT9), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n294), .A2(new_n277), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n216), .B2(new_n296), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT9), .ZN(new_n308));
  NOR2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n302), .B1(new_n305), .B2(new_n309), .ZN(new_n310));
  AOI22_X1  g0110(.A1(new_n307), .A2(new_n308), .B1(G200), .B2(new_n272), .ZN(new_n311));
  INV_X1    g0111(.A(new_n302), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n298), .A2(KEYINPUT9), .ZN(new_n313));
  NAND4_X1  g0113(.A1(new_n311), .A2(new_n312), .A3(new_n313), .A4(new_n304), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n299), .B1(new_n310), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n217), .A2(new_n258), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n219), .A2(G1698), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n253), .A2(new_n316), .A3(new_n255), .A4(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G33), .A2(G97), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n318), .A2(KEYINPUT75), .A3(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(KEYINPUT75), .B1(new_n318), .B2(new_n319), .ZN(new_n322));
  NOR3_X1   g0122(.A1(new_n321), .A2(new_n322), .A3(new_n263), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT76), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n271), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n263), .A2(KEYINPUT76), .A3(new_n267), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(G238), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(new_n270), .ZN(new_n328));
  OAI21_X1  g0128(.A(KEYINPUT13), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(new_n328), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT13), .ZN(new_n331));
  INV_X1    g0131(.A(new_n322), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n332), .A2(new_n264), .A3(new_n320), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT77), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n330), .A2(new_n333), .A3(KEYINPUT77), .A4(new_n331), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(G169), .A3(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT14), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n336), .A2(new_n340), .A3(G169), .A4(new_n337), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n329), .A2(new_n334), .A3(G179), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n339), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n287), .A2(G77), .ZN(new_n344));
  INV_X1    g0144(.A(new_n292), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n344), .B1(new_n289), .B2(G68), .C1(new_n216), .C2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(new_n280), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT11), .ZN(new_n348));
  OAI21_X1  g0148(.A(KEYINPUT12), .B1(new_n276), .B2(G68), .ZN(new_n349));
  OR3_X1    g0149(.A1(new_n276), .A2(KEYINPUT12), .A3(G68), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n297), .A2(G68), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  AND2_X1   g0151(.A1(new_n348), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n336), .A2(G200), .A3(new_n337), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n329), .A2(new_n334), .A3(G190), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n355), .A2(new_n352), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(KEYINPUT78), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT78), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n355), .A2(new_n359), .A3(new_n352), .A4(new_n356), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n358), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(G238), .A2(G1698), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n257), .B(new_n362), .C1(new_n219), .C2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n363), .B(new_n264), .C1(G107), .C2(new_n257), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n271), .A2(new_n208), .ZN(new_n365));
  OR3_X1    g0165(.A1(new_n365), .A2(KEYINPUT72), .A3(new_n269), .ZN(new_n366));
  OAI21_X1  g0166(.A(KEYINPUT72), .B1(new_n365), .B2(new_n269), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n364), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OR2_X1    g0168(.A1(new_n368), .A2(G179), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n297), .A2(G77), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n282), .A2(new_n345), .B1(new_n289), .B2(new_n207), .ZN(new_n371));
  XOR2_X1   g0171(.A(KEYINPUT15), .B(G87), .Z(new_n372));
  AOI21_X1  g0172(.A(new_n371), .B1(new_n287), .B2(new_n372), .ZN(new_n373));
  OAI221_X1 g0173(.A(new_n370), .B1(G77), .B2(new_n276), .C1(new_n373), .C2(new_n281), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n368), .A2(new_n273), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(new_n374), .A3(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n315), .A2(new_n354), .A3(new_n361), .A4(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n253), .ZN(new_n378));
  XNOR2_X1  g0178(.A(KEYINPUT79), .B(KEYINPUT3), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(G33), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n260), .A2(new_n258), .ZN(new_n381));
  OAI211_X1 g0181(.A(new_n380), .B(new_n381), .C1(G226), .C2(new_n258), .ZN(new_n382));
  NAND2_X1  g0182(.A1(G33), .A2(G87), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n263), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n270), .B1(new_n271), .B2(new_n219), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n273), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(G179), .ZN(new_n389));
  NOR3_X1   g0189(.A1(new_n384), .A2(new_n389), .A3(new_n386), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n388), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n218), .A2(new_n211), .ZN(new_n392));
  OAI21_X1  g0192(.A(G20), .B1(new_n392), .B2(new_n290), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n292), .A2(G159), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AND2_X1   g0196(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n397));
  NOR2_X1   g0197(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n398));
  OAI21_X1  g0198(.A(G33), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(G20), .B1(new_n399), .B2(new_n253), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  OAI21_X1  g0201(.A(G68), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR3_X1   g0202(.A1(new_n380), .A2(KEYINPUT7), .A3(G20), .ZN(new_n403));
  OAI211_X1 g0203(.A(KEYINPUT16), .B(new_n396), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT79), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n254), .ZN(new_n406));
  NAND2_X1  g0206(.A1(KEYINPUT79), .A2(KEYINPUT3), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n252), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(new_n255), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n409), .A2(KEYINPUT7), .A3(new_n289), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT7), .B1(new_n256), .B2(new_n289), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n395), .B1(new_n413), .B2(G68), .ZN(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n415));
  OAI211_X1 g0215(.A(new_n404), .B(new_n280), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n286), .A2(new_n276), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n417), .B1(new_n297), .B2(new_n286), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n416), .A2(KEYINPUT81), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT81), .B1(new_n416), .B2(new_n418), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n391), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  OAI211_X1 g0224(.A(KEYINPUT18), .B(new_n391), .C1(new_n420), .C2(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n385), .A2(G190), .A3(new_n387), .ZN(new_n427));
  OAI21_X1  g0227(.A(G200), .B1(new_n384), .B2(new_n386), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n416), .A2(new_n427), .A3(new_n428), .A4(new_n418), .ZN(new_n429));
  XNOR2_X1  g0229(.A(new_n429), .B(KEYINPUT17), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n368), .A2(G200), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n374), .A2(KEYINPUT73), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n374), .A2(KEYINPUT73), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n431), .B1(new_n303), .B2(new_n368), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n426), .A2(new_n430), .A3(new_n434), .ZN(new_n435));
  OR2_X1    g0235(.A1(new_n377), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(G257), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n438), .A2(new_n258), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n213), .A2(G1698), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n399), .A2(new_n253), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n256), .A2(G303), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(new_n264), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT90), .ZN(new_n445));
  INV_X1    g0245(.A(G45), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(G1), .ZN(new_n447));
  NOR2_X1   g0247(.A1(KEYINPUT5), .A2(G41), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT5), .A2(G41), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n447), .B(G274), .C1(new_n448), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n447), .B1(new_n449), .B2(new_n448), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n452), .A2(new_n263), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n451), .B1(new_n454), .B2(G270), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT90), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n443), .A2(new_n456), .A3(new_n264), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n445), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  AOI21_X1  g0258(.A(G20), .B1(G33), .B2(G283), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n459), .B1(G33), .B2(new_n202), .ZN(new_n460));
  XOR2_X1   g0260(.A(KEYINPUT88), .B(G116), .Z(new_n461));
  OAI211_X1 g0261(.A(new_n280), .B(new_n460), .C1(new_n461), .C2(new_n289), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT20), .ZN(new_n463));
  XNOR2_X1  g0263(.A(new_n462), .B(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n461), .A2(new_n276), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n276), .ZN(new_n467));
  AOI211_X1 g0267(.A(new_n280), .B(new_n467), .C1(new_n266), .C2(G33), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n468), .A2(G116), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n464), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n458), .A2(new_n470), .A3(G169), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(KEYINPUT21), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT21), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n458), .A2(new_n470), .A3(new_n473), .A4(G169), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n470), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n445), .A2(G179), .A3(new_n455), .A4(new_n457), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT91), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n458), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT91), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n479), .A2(new_n470), .A3(new_n480), .A4(G179), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n458), .A2(G200), .ZN(new_n483));
  OAI211_X1 g0283(.A(new_n483), .B(new_n476), .C1(new_n303), .C2(new_n458), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n475), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT22), .ZN(new_n486));
  INV_X1    g0286(.A(G87), .ZN(new_n487));
  NOR3_X1   g0287(.A1(new_n486), .A2(new_n487), .A3(G20), .ZN(new_n488));
  NAND4_X1  g0288(.A1(new_n253), .A2(new_n255), .A3(new_n289), .A4(G87), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n380), .A2(new_n488), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n461), .A2(new_n287), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n289), .A2(G107), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT23), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n490), .A2(KEYINPUT24), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n399), .A2(new_n253), .A3(new_n488), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n489), .A2(new_n486), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n493), .A2(new_n495), .A3(new_n496), .A4(new_n491), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT24), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n494), .A2(new_n499), .A3(new_n280), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n468), .A2(G107), .ZN(new_n501));
  OR3_X1    g0301(.A1(new_n276), .A2(KEYINPUT92), .A3(G107), .ZN(new_n502));
  OAI21_X1  g0302(.A(KEYINPUT92), .B1(new_n276), .B2(G107), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n504), .B(KEYINPUT25), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n500), .A2(new_n501), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(G250), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n258), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n438), .A2(G1698), .ZN(new_n509));
  NAND4_X1  g0309(.A1(new_n399), .A2(new_n253), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(G33), .A2(G294), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n263), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n453), .A2(new_n213), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(new_n450), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n303), .ZN(new_n516));
  INV_X1    g0316(.A(G200), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n514), .B2(new_n450), .ZN(new_n518));
  OR3_X1    g0318(.A1(new_n506), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NOR4_X1   g0319(.A1(new_n512), .A2(new_n513), .A3(G179), .A4(new_n451), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n520), .B1(new_n515), .B2(new_n273), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT93), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n521), .A2(new_n506), .A3(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n522), .B1(new_n521), .B2(new_n506), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n519), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n485), .A2(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n372), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n467), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n212), .A2(new_n258), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n208), .A2(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n399), .A2(new_n253), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n461), .A2(G33), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n264), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n266), .A2(new_n268), .A3(G45), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n263), .B(new_n535), .C1(G250), .C2(new_n447), .ZN(new_n536));
  XNOR2_X1  g0336(.A(new_n536), .B(KEYINPUT87), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G200), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT19), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n287), .A2(new_n540), .A3(G97), .ZN(new_n541));
  NOR2_X1   g0341(.A1(G97), .A2(G107), .ZN(new_n542));
  AOI22_X1  g0342(.A1(new_n542), .A2(new_n487), .B1(new_n319), .B2(new_n289), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n543), .B2(new_n540), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n399), .A2(new_n289), .A3(G68), .A4(new_n253), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT89), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n544), .A2(new_n545), .A3(KEYINPUT89), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n548), .A2(new_n280), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n468), .A2(G87), .ZN(new_n551));
  AND4_X1   g0351(.A1(new_n528), .A2(new_n539), .A3(new_n550), .A4(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(new_n538), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(G190), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n468), .ZN(new_n556));
  OAI211_X1 g0356(.A(new_n550), .B(new_n528), .C1(new_n527), .C2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n273), .B1(new_n534), .B2(new_n537), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n534), .A2(new_n537), .A3(G179), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n557), .B1(new_n558), .B2(new_n560), .ZN(new_n561));
  AND2_X1   g0361(.A1(new_n555), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT85), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n563), .B1(new_n467), .B2(new_n202), .ZN(new_n564));
  NOR3_X1   g0364(.A1(new_n276), .A2(KEYINPUT85), .A3(G97), .ZN(new_n565));
  OAI22_X1  g0365(.A1(new_n556), .A2(new_n202), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(G97), .A2(G107), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT82), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n569), .A2(KEYINPUT6), .ZN(new_n570));
  AND2_X1   g0370(.A1(KEYINPUT6), .A2(G107), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n204), .B(new_n568), .C1(new_n570), .C2(new_n571), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT83), .ZN(new_n573));
  INV_X1    g0373(.A(new_n568), .ZN(new_n574));
  OAI22_X1  g0374(.A1(new_n574), .A2(new_n542), .B1(new_n569), .B2(KEYINPUT6), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n573), .B1(new_n572), .B2(new_n575), .ZN(new_n577));
  OAI21_X1  g0377(.A(G20), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  AOI211_X1 g0378(.A(new_n401), .B(G20), .C1(new_n408), .C2(new_n255), .ZN(new_n579));
  OAI21_X1  g0379(.A(G107), .B1(new_n579), .B2(new_n411), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n292), .A2(G77), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT84), .ZN(new_n583));
  AND3_X1   g0383(.A1(new_n582), .A2(new_n583), .A3(new_n280), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n583), .B1(new_n582), .B2(new_n280), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n567), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n453), .A2(new_n438), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT4), .B1(new_n256), .B2(new_n507), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n588), .A2(G1698), .B1(G33), .B2(G283), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n399), .A2(new_n253), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n590), .B1(new_n591), .B2(new_n208), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n257), .A2(KEYINPUT4), .A3(G244), .A4(new_n258), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI211_X1 g0394(.A(new_n451), .B(new_n587), .C1(new_n594), .C2(new_n264), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G179), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n594), .A2(new_n264), .ZN(new_n597));
  INV_X1    g0397(.A(new_n587), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n597), .A2(new_n450), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(G169), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n596), .A2(new_n600), .ZN(new_n601));
  AND2_X1   g0401(.A1(new_n586), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT86), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n586), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(G20), .B1(new_n408), .B2(new_n255), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n411), .B1(new_n605), .B2(KEYINPUT7), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n581), .B1(new_n606), .B2(new_n203), .ZN(new_n607));
  INV_X1    g0407(.A(new_n577), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n609));
  AOI21_X1  g0409(.A(new_n289), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n280), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT84), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n582), .A2(new_n583), .A3(new_n280), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(KEYINPUT86), .A3(new_n567), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n604), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n599), .A2(new_n303), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n617), .B1(G200), .B2(new_n599), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n602), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND4_X1   g0419(.A1(new_n437), .A2(new_n526), .A3(new_n562), .A4(new_n619), .ZN(G372));
  AOI21_X1  g0420(.A(KEYINPUT86), .B1(new_n614), .B2(new_n567), .ZN(new_n621));
  AOI211_X1 g0421(.A(new_n603), .B(new_n566), .C1(new_n612), .C2(new_n613), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT87), .ZN(new_n624));
  XNOR2_X1  g0424(.A(new_n536), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n263), .B1(new_n531), .B2(new_n532), .ZN(new_n626));
  OAI21_X1  g0426(.A(G169), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT94), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n559), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n628), .B1(new_n627), .B2(new_n559), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n557), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND3_X1   g0432(.A1(new_n519), .A2(new_n555), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n586), .A2(new_n601), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n521), .A2(new_n506), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n475), .A2(new_n482), .A3(new_n635), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n623), .A2(new_n633), .A3(new_n634), .A4(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n621), .A2(new_n622), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  INV_X1    g0439(.A(new_n631), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n629), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n641), .A2(new_n557), .B1(new_n552), .B2(new_n554), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n638), .A2(new_n639), .A3(new_n601), .A4(new_n642), .ZN(new_n643));
  INV_X1    g0443(.A(new_n632), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n555), .A2(new_n586), .A3(new_n601), .A4(new_n561), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n644), .B1(new_n645), .B2(KEYINPUT26), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n637), .A2(new_n643), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n437), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n416), .A2(new_n418), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n388), .A2(new_n390), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n423), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n391), .A2(KEYINPUT18), .A3(new_n649), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n376), .ZN(new_n655));
  AOI22_X1  g0455(.A1(new_n343), .A2(new_n353), .B1(new_n357), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(new_n430), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n310), .A2(new_n314), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n299), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n648), .A2(new_n660), .ZN(G369));
  NAND2_X1  g0461(.A1(new_n475), .A2(new_n482), .ZN(new_n662));
  INV_X1    g0462(.A(G13), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(G20), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n266), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n476), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n662), .A2(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n673), .B1(new_n485), .B2(new_n672), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT95), .Z(new_n675));
  AND2_X1   g0475(.A1(new_n506), .A2(new_n670), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n525), .A2(new_n676), .B1(new_n635), .B2(new_n671), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n675), .A2(G330), .A3(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n525), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n670), .B1(new_n475), .B2(new_n482), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n635), .B2(new_n670), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n678), .A2(new_n683), .ZN(G399));
  NOR3_X1   g0484(.A1(new_n204), .A2(G87), .A3(G116), .ZN(new_n685));
  INV_X1    g0485(.A(G41), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n224), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n685), .A2(new_n687), .A3(G1), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n230), .B2(new_n687), .ZN(new_n689));
  XOR2_X1   g0489(.A(new_n689), .B(KEYINPUT28), .Z(new_n690));
  XNOR2_X1  g0490(.A(new_n632), .B(KEYINPUT96), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n642), .A2(new_n604), .A3(new_n601), .A4(new_n615), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n691), .B1(new_n692), .B2(KEYINPUT26), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n475), .B(new_n482), .C1(new_n524), .C2(new_n523), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n623), .A2(new_n694), .A3(new_n633), .A4(new_n634), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n562), .A2(new_n639), .A3(new_n602), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(KEYINPUT29), .A3(new_n671), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT97), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n647), .A2(new_n671), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT29), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT97), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n700), .B1(new_n698), .B2(new_n703), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n619), .A2(new_n526), .A3(new_n562), .A4(new_n671), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n595), .A2(new_n479), .A3(new_n514), .A4(new_n560), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT30), .ZN(new_n707));
  OR2_X1    g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n706), .A2(new_n707), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n553), .A2(G179), .ZN(new_n710));
  NAND4_X1  g0510(.A1(new_n710), .A2(new_n599), .A3(new_n515), .A4(new_n458), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n708), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(new_n670), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n713), .ZN(new_n714));
  OR2_X1    g0514(.A1(new_n713), .A2(KEYINPUT31), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n716), .A2(G330), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n704), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n690), .B1(new_n718), .B2(new_n266), .ZN(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT98), .ZN(G364));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(new_n289), .ZN(new_n722));
  XOR2_X1   g0522(.A(new_n722), .B(KEYINPUT102), .Z(new_n723));
  OR2_X1    g0523(.A1(new_n675), .A2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n279), .B1(G20), .B2(new_n273), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT100), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT100), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n289), .A2(new_n303), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n389), .A2(new_n517), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n216), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n517), .A2(G179), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n729), .A2(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n257), .B1(new_n734), .B2(new_n487), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT101), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n289), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n730), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G68), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT32), .ZN(new_n741));
  NOR2_X1   g0541(.A1(G179), .A2(G200), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n737), .A2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n741), .B1(new_n744), .B2(G159), .ZN(new_n745));
  INV_X1    g0545(.A(G159), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n743), .A2(KEYINPUT32), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n737), .A2(new_n733), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n203), .ZN(new_n749));
  NOR3_X1   g0549(.A1(new_n745), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n389), .A2(G200), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n729), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  AOI21_X1  g0553(.A(new_n289), .B1(new_n742), .B2(G190), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n753), .A2(G58), .B1(new_n755), .B2(G97), .ZN(new_n756));
  NAND4_X1  g0556(.A1(new_n736), .A2(new_n740), .A3(new_n750), .A4(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n737), .A2(new_n751), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI211_X1 g0559(.A(new_n732), .B(new_n757), .C1(G77), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G317), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT33), .ZN(new_n762));
  OR2_X1    g0562(.A1(new_n761), .A2(KEYINPUT33), .ZN(new_n763));
  NAND3_X1  g0563(.A1(new_n739), .A2(new_n762), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n744), .A2(G329), .ZN(new_n765));
  INV_X1    g0565(.A(G283), .ZN(new_n766));
  OAI211_X1 g0566(.A(new_n764), .B(new_n765), .C1(new_n766), .C2(new_n748), .ZN(new_n767));
  INV_X1    g0567(.A(new_n731), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n767), .B1(G326), .B2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n734), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G303), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n257), .B1(new_n753), .B2(G322), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n755), .A2(G294), .ZN(new_n773));
  NAND4_X1  g0573(.A1(new_n769), .A2(new_n771), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G311), .B2(new_n759), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n728), .B1(new_n760), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g0576(.A1(G355), .A2(new_n224), .A3(new_n257), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n246), .A2(new_n446), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n591), .A2(new_n224), .ZN(new_n779));
  XNOR2_X1  g0579(.A(new_n779), .B(KEYINPUT99), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n780), .B1(G45), .B2(new_n230), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n777), .B1(G116), .B2(new_n224), .C1(new_n778), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n722), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n728), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n664), .A2(G45), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n687), .A2(G1), .A3(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND4_X1  g0588(.A1(new_n724), .A2(new_n776), .A3(new_n785), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n675), .A2(G330), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n675), .A2(G330), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(new_n787), .ZN(new_n792));
  OAI21_X1  g0592(.A(new_n789), .B1(new_n790), .B2(new_n792), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT103), .Z(G396));
  NAND2_X1  g0594(.A1(new_n374), .A2(new_n670), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n434), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(new_n376), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n655), .A2(new_n671), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n701), .B(new_n800), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(new_n717), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(new_n787), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G143), .A2(new_n753), .B1(new_n759), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(G137), .ZN(new_n805));
  INV_X1    g0605(.A(G150), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n804), .B1(new_n805), .B2(new_n731), .C1(new_n806), .C2(new_n738), .ZN(new_n807));
  XOR2_X1   g0607(.A(new_n807), .B(KEYINPUT34), .Z(new_n808));
  AOI211_X1 g0608(.A(new_n591), .B(new_n808), .C1(G132), .C2(new_n744), .ZN(new_n809));
  INV_X1    g0609(.A(new_n748), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n810), .A2(G68), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n809), .B(new_n811), .C1(new_n216), .C2(new_n734), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(G58), .B2(new_n755), .ZN(new_n813));
  AOI22_X1  g0613(.A1(G311), .A2(new_n744), .B1(new_n755), .B2(G97), .ZN(new_n814));
  XOR2_X1   g0614(.A(KEYINPUT104), .B(G283), .Z(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n814), .B1(new_n738), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(new_n817), .B1(G303), .B2(new_n768), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n748), .A2(new_n487), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n257), .B(new_n819), .C1(new_n461), .C2(new_n759), .ZN(new_n820));
  INV_X1    g0620(.A(G294), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n818), .B(new_n820), .C1(new_n821), .C2(new_n752), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(G107), .B2(new_n770), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n728), .B1(new_n813), .B2(new_n823), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n728), .A2(new_n721), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n207), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n799), .A2(new_n721), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n788), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  AND2_X1   g0628(.A1(new_n803), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(G384));
  INV_X1    g0630(.A(KEYINPUT40), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT38), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT107), .ZN(new_n833));
  OAI21_X1  g0633(.A(KEYINPUT7), .B1(new_n380), .B2(G20), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n591), .A2(new_n401), .A3(new_n289), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n834), .A2(G68), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n415), .B1(new_n836), .B2(new_n396), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n833), .B1(new_n837), .B2(new_n281), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n252), .B1(new_n406), .B2(new_n407), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n289), .B1(new_n839), .B2(new_n378), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n211), .B1(new_n840), .B2(KEYINPUT7), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n395), .B1(new_n841), .B2(new_n835), .ZN(new_n842));
  OAI211_X1 g0642(.A(KEYINPUT107), .B(new_n280), .C1(new_n842), .C2(new_n415), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n838), .A2(new_n404), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n651), .B1(new_n844), .B2(new_n418), .ZN(new_n845));
  INV_X1    g0645(.A(new_n429), .ZN(new_n846));
  OAI21_X1  g0646(.A(KEYINPUT108), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT108), .ZN(new_n848));
  INV_X1    g0648(.A(new_n418), .ZN(new_n849));
  INV_X1    g0649(.A(new_n404), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n280), .B1(new_n842), .B2(new_n415), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n850), .B1(new_n851), .B2(new_n833), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n849), .B1(new_n852), .B2(new_n843), .ZN(new_n853));
  OAI211_X1 g0653(.A(new_n848), .B(new_n429), .C1(new_n853), .C2(new_n651), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n844), .A2(new_n418), .ZN(new_n855));
  INV_X1    g0655(.A(new_n668), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n847), .A2(new_n854), .A3(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT109), .ZN(new_n859));
  INV_X1    g0659(.A(KEYINPUT81), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n649), .A2(new_n860), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n861), .A2(new_n419), .B1(new_n651), .B2(new_n668), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT37), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n429), .A2(new_n863), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n859), .B1(new_n862), .B2(new_n864), .ZN(new_n865));
  OAI22_X1  g0665(.A1(new_n420), .A2(new_n421), .B1(new_n391), .B2(new_n856), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n866), .A2(KEYINPUT109), .A3(new_n863), .A4(new_n429), .ZN(new_n867));
  AOI22_X1  g0667(.A1(new_n858), .A2(KEYINPUT37), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n857), .B1(new_n426), .B2(new_n430), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n832), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(new_n425), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n861), .A2(new_n419), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT18), .B1(new_n872), .B2(new_n391), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n430), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n853), .A2(new_n668), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n429), .B1(new_n853), .B2(new_n651), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n875), .B1(new_n877), .B2(KEYINPUT108), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n863), .B1(new_n878), .B2(new_n854), .ZN(new_n879));
  AND2_X1   g0679(.A1(new_n867), .A2(new_n865), .ZN(new_n880));
  OAI211_X1 g0680(.A(KEYINPUT38), .B(new_n876), .C1(new_n879), .C2(new_n880), .ZN(new_n881));
  AND2_X1   g0681(.A1(new_n870), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n354), .A2(new_n361), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n352), .A2(new_n671), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OAI211_X1 g0685(.A(new_n354), .B(new_n357), .C1(new_n352), .C2(new_n671), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n799), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n887), .A2(new_n714), .A3(new_n715), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n831), .B1(new_n882), .B2(new_n888), .ZN(new_n889));
  AND4_X1   g0689(.A1(KEYINPUT40), .A2(new_n887), .A3(new_n714), .A4(new_n715), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT110), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n872), .A2(new_n856), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(new_n654), .B2(new_n430), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n867), .A2(new_n865), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n846), .B1(new_n649), .B2(new_n391), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n892), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(KEYINPUT37), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n893), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n891), .B1(new_n898), .B2(KEYINPUT38), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n865), .A2(new_n867), .B1(new_n896), .B2(KEYINPUT37), .ZN(new_n900));
  OAI211_X1 g0700(.A(KEYINPUT110), .B(new_n832), .C1(new_n900), .C2(new_n893), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n899), .A2(new_n901), .A3(new_n881), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n889), .A2(G330), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n437), .A2(new_n716), .A3(G330), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT111), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n889), .A2(new_n716), .A3(new_n903), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n907), .B1(new_n436), .B2(new_n908), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT39), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n910), .B1(new_n911), .B2(new_n902), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n354), .A2(new_n670), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n654), .A2(new_n856), .ZN(new_n915));
  INV_X1    g0715(.A(new_n882), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n885), .A2(new_n886), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n647), .A2(new_n671), .A3(new_n800), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n918), .B1(new_n798), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n915), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  AND2_X1   g0721(.A1(new_n914), .A2(new_n921), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n704), .A2(new_n436), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n923), .A2(new_n660), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  XNOR2_X1  g0725(.A(new_n909), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n926), .B1(new_n266), .B2(new_n664), .ZN(new_n927));
  NOR3_X1   g0727(.A1(new_n230), .A2(new_n207), .A3(new_n392), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n211), .A2(G50), .ZN(new_n929));
  OAI211_X1 g0729(.A(G1), .B(new_n663), .C1(new_n928), .C2(new_n929), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n576), .A2(new_n577), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n931), .B(KEYINPUT105), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT35), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n227), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI211_X1 g0734(.A(new_n934), .B(G116), .C1(new_n933), .C2(new_n932), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(KEYINPUT106), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT36), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n927), .A2(new_n930), .A3(new_n937), .ZN(G367));
  INV_X1    g0738(.A(new_n780), .ZN(new_n939));
  OAI221_X1 g0739(.A(new_n784), .B1(new_n224), .B2(new_n527), .C1(new_n939), .C2(new_n241), .ZN(new_n940));
  OAI22_X1  g0740(.A1(new_n218), .A2(new_n734), .B1(new_n752), .B2(new_n806), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n768), .A2(G143), .B1(new_n755), .B2(G68), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n942), .B1(new_n805), .B2(new_n743), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n941), .B(new_n943), .C1(G159), .C2(new_n739), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n810), .A2(G77), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n759), .A2(G50), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n944), .A2(new_n257), .A3(new_n945), .A4(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(G311), .ZN(new_n948));
  INV_X1    g0748(.A(G303), .ZN(new_n949));
  OAI22_X1  g0749(.A1(new_n731), .A2(new_n948), .B1(new_n752), .B2(new_n949), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT112), .Z(new_n951));
  INV_X1    g0751(.A(KEYINPUT46), .ZN(new_n952));
  INV_X1    g0752(.A(new_n461), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(new_n734), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n810), .A2(G97), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n770), .A2(KEYINPUT46), .A3(G116), .ZN(new_n956));
  NAND4_X1  g0756(.A1(new_n954), .A2(new_n591), .A3(new_n955), .A4(new_n956), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n951), .A2(new_n957), .ZN(new_n958));
  AOI22_X1  g0758(.A1(G294), .A2(new_n739), .B1(new_n759), .B2(new_n815), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n958), .B(new_n959), .C1(new_n761), .C2(new_n743), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n754), .A2(new_n203), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n947), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(new_n962), .B(KEYINPUT47), .Z(new_n963));
  INV_X1    g0763(.A(new_n728), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n788), .B(new_n940), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(KEYINPUT113), .Z(new_n966));
  INV_X1    g0766(.A(new_n642), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n550), .A2(new_n528), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n671), .B1(new_n968), .B2(new_n551), .ZN(new_n969));
  OR2_X1    g0769(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n644), .A2(new_n969), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n966), .B1(new_n723), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n786), .A2(G1), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n619), .B1(new_n616), .B2(new_n671), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n638), .A2(new_n601), .A3(new_n670), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n977), .A2(new_n683), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT45), .Z(new_n979));
  NOR2_X1   g0779(.A1(new_n977), .A2(new_n683), .ZN(new_n980));
  XNOR2_X1  g0780(.A(new_n980), .B(KEYINPUT44), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  XOR2_X1   g0782(.A(new_n982), .B(new_n678), .Z(new_n983));
  OAI21_X1  g0783(.A(new_n681), .B1(new_n677), .B2(new_n680), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n791), .B(new_n984), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n717), .B(new_n704), .C1(new_n983), .C2(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n687), .B(KEYINPUT41), .Z(new_n987));
  AOI21_X1  g0787(.A(new_n974), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n681), .B1(new_n975), .B2(new_n976), .ZN(new_n990));
  XOR2_X1   g0790(.A(new_n990), .B(KEYINPUT42), .Z(new_n991));
  NOR2_X1   g0791(.A1(new_n523), .A2(new_n524), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n977), .A2(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n670), .B1(new_n993), .B2(new_n634), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n989), .B1(new_n991), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n678), .B1(new_n975), .B2(new_n976), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n997), .B(new_n998), .Z(new_n999));
  OAI21_X1  g0799(.A(new_n973), .B1(new_n988), .B2(new_n999), .ZN(G387));
  OR2_X1    g0800(.A1(new_n718), .A2(new_n985), .ZN(new_n1001));
  INV_X1    g0801(.A(new_n687), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n718), .A2(new_n985), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n591), .B1(G77), .B2(new_n770), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n1005), .B(new_n955), .C1(new_n806), .C2(new_n743), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT114), .Z(new_n1007));
  AOI21_X1  g0807(.A(new_n1007), .B1(new_n286), .B2(new_n739), .ZN(new_n1008));
  OAI22_X1  g0808(.A1(new_n527), .A2(new_n754), .B1(new_n216), .B2(new_n752), .ZN(new_n1009));
  XNOR2_X1  g0809(.A(new_n1009), .B(KEYINPUT115), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n768), .A2(G159), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n759), .A2(G68), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1008), .A2(new_n1010), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AOI22_X1  g0813(.A1(G322), .A2(new_n768), .B1(new_n739), .B2(G311), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n949), .B2(new_n758), .C1(new_n761), .C2(new_n752), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1015), .B(KEYINPUT48), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n1016), .B1(new_n821), .B2(new_n734), .C1(new_n754), .C2(new_n816), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT49), .Z(new_n1018));
  INV_X1    g0818(.A(G326), .ZN(new_n1019));
  OAI221_X1 g0819(.A(new_n591), .B1(new_n1019), .B2(new_n743), .C1(new_n953), .C2(new_n748), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1013), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n728), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n282), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n216), .ZN(new_n1024));
  XNOR2_X1  g0824(.A(new_n1024), .B(KEYINPUT50), .ZN(new_n1025));
  NOR2_X1   g0825(.A1(new_n211), .A2(new_n207), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n685), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1025), .A2(G45), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n780), .B1(new_n238), .B2(new_n446), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1027), .A2(new_n224), .A3(new_n257), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1028), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n224), .A2(G107), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n784), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OR2_X1    g0833(.A1(new_n677), .A2(new_n723), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1022), .A2(new_n788), .A3(new_n1033), .A4(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g0835(.A(new_n1035), .B(KEYINPUT116), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n974), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1004), .B(new_n1036), .C1(new_n1037), .C2(new_n985), .ZN(G393));
  OAI22_X1  g0838(.A1(new_n738), .A2(new_n216), .B1(new_n754), .B2(new_n207), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n731), .A2(new_n806), .B1(new_n752), .B2(new_n746), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT51), .Z(new_n1041));
  AOI211_X1 g0841(.A(new_n1039), .B(new_n1041), .C1(G68), .C2(new_n770), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n819), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n759), .A2(new_n1023), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n591), .B1(G143), .B2(new_n744), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1042), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  NOR2_X1   g0846(.A1(new_n738), .A2(new_n949), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n731), .A2(new_n761), .B1(new_n752), .B2(new_n948), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT52), .Z(new_n1049));
  AOI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(G322), .C2(new_n744), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n755), .A2(new_n461), .ZN(new_n1051));
  NOR2_X1   g0851(.A1(new_n758), .A2(new_n821), .ZN(new_n1052));
  AOI211_X1 g0852(.A(new_n749), .B(new_n1052), .C1(new_n770), .C2(new_n815), .ZN(new_n1053));
  NAND4_X1  g0853(.A1(new_n1050), .A2(new_n256), .A3(new_n1051), .A4(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n964), .B1(new_n1046), .B2(new_n1054), .ZN(new_n1055));
  NOR2_X1   g0855(.A1(new_n224), .A2(new_n202), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n784), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n1056), .B(new_n1057), .C1(new_n250), .C2(new_n780), .ZN(new_n1058));
  NOR3_X1   g0858(.A1(new_n1055), .A2(new_n787), .A3(new_n1058), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1059), .B1(new_n977), .B2(new_n722), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n1060), .B1(new_n983), .B2(new_n1037), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n983), .A2(new_n1001), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n687), .B1(new_n983), .B2(new_n1001), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(G390));
  OAI211_X1 g0865(.A(new_n660), .B(new_n905), .C1(new_n704), .C2(new_n436), .ZN(new_n1066));
  NAND4_X1  g0866(.A1(new_n714), .A2(new_n715), .A3(G330), .A4(new_n800), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n918), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT117), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  OR2_X1    g0870(.A1(new_n1067), .A2(new_n918), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n697), .A2(new_n671), .A3(new_n797), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n798), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1067), .A2(KEYINPUT117), .A3(new_n918), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n1070), .A2(new_n1071), .A3(new_n1074), .A4(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1074), .ZN(new_n1078));
  AOI21_X1  g0878(.A(KEYINPUT117), .B1(new_n1067), .B2(new_n918), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1067), .A2(new_n918), .ZN(new_n1080));
  NOR2_X1   g0880(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT118), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1078), .A2(new_n1081), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1071), .A2(new_n1068), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n919), .A2(new_n798), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1066), .B1(new_n1084), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n913), .B1(new_n1086), .B2(new_n917), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n902), .A2(new_n911), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n870), .A2(new_n881), .A3(KEYINPUT39), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1089), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1073), .A2(new_n917), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n913), .ZN(new_n1094));
  AND3_X1   g0894(.A1(new_n1093), .A2(new_n902), .A3(new_n1094), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n1080), .B1(new_n1092), .B2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1093), .A2(new_n902), .A3(new_n1094), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1097), .B(new_n1071), .C1(new_n912), .C2(new_n1089), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1088), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n1076), .A2(KEYINPUT118), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n1082), .B1(new_n1078), .B2(new_n1081), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1087), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1066), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  AND3_X1   g0906(.A1(new_n1099), .A2(new_n1106), .A3(new_n1002), .ZN(new_n1107));
  NOR3_X1   g0907(.A1(new_n912), .A2(G13), .A3(G33), .ZN(new_n1108));
  INV_X1    g0908(.A(G128), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n731), .A2(new_n1109), .B1(new_n748), .B2(new_n216), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n770), .A2(G150), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1111), .B(KEYINPUT53), .ZN(new_n1112));
  INV_X1    g0912(.A(G132), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n257), .B1(new_n752), .B2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n746), .B2(new_n754), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1110), .B(new_n1116), .C1(G125), .C2(new_n744), .ZN(new_n1117));
  XOR2_X1   g0917(.A(KEYINPUT54), .B(G143), .Z(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  OAI221_X1 g0919(.A(new_n1117), .B1(new_n805), .B2(new_n738), .C1(new_n758), .C2(new_n1119), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n811), .B1(new_n487), .B2(new_n734), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n738), .A2(new_n203), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n256), .B1(new_n754), .B2(new_n207), .ZN(new_n1123));
  OAI22_X1  g0923(.A1(new_n731), .A2(new_n766), .B1(new_n743), .B2(new_n821), .ZN(new_n1124));
  NOR4_X1   g0924(.A1(new_n1121), .A2(new_n1122), .A3(new_n1123), .A4(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(G116), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1125), .B1(new_n202), .B2(new_n758), .C1(new_n1126), .C2(new_n752), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n964), .B1(new_n1120), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n286), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n787), .B(new_n1128), .C1(new_n1129), .C2(new_n825), .ZN(new_n1130));
  XOR2_X1   g0930(.A(new_n1130), .B(KEYINPUT119), .Z(new_n1131));
  OAI22_X1  g0931(.A1(new_n1105), .A2(new_n1037), .B1(new_n1108), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT120), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1132), .B(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1107), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G378));
  NAND2_X1  g0936(.A1(new_n914), .A2(new_n921), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n299), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n659), .A2(new_n1138), .ZN(new_n1139));
  XOR2_X1   g0939(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1140));
  NAND2_X1  g0940(.A1(new_n1139), .A2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n298), .A2(new_n668), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n315), .A2(new_n1143), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1141), .A2(new_n1142), .A3(new_n1144), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1142), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1143), .B1(new_n659), .B2(new_n1138), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n299), .B(new_n1140), .C1(new_n310), .C2(new_n314), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AND3_X1   g0949(.A1(new_n1145), .A2(new_n1149), .A3(KEYINPUT122), .ZN(new_n1150));
  AOI21_X1  g0950(.A(KEYINPUT122), .B1(new_n1145), .B2(new_n1149), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n889), .A2(G330), .A3(new_n903), .A4(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1145), .A2(new_n1149), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1153), .A2(KEYINPUT123), .B1(new_n904), .B2(new_n1154), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n1154), .ZN(new_n1156));
  OAI21_X1  g0956(.A(new_n1137), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1153), .A2(KEYINPUT123), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n904), .A2(new_n1154), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n904), .A2(KEYINPUT123), .A3(new_n1154), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1160), .A2(new_n922), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(KEYINPUT124), .B1(new_n1157), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT124), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n922), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n974), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n721), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n752), .A2(new_n1109), .B1(new_n758), .B2(new_n805), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n1119), .A2(new_n734), .B1(new_n806), .B2(new_n754), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1169), .B(new_n1170), .C1(G125), .C2(new_n768), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1171), .B1(new_n1113), .B2(new_n738), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT59), .Z(new_n1173));
  NAND2_X1  g0973(.A1(new_n744), .A2(G124), .ZN(new_n1174));
  AOI211_X1 g0974(.A(G33), .B(G41), .C1(new_n810), .C2(G159), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1173), .A2(new_n1174), .A3(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(G50), .B1(new_n252), .B2(new_n686), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n380), .B2(G41), .ZN(new_n1178));
  OAI22_X1  g0978(.A1(new_n731), .A2(new_n1126), .B1(new_n754), .B2(new_n211), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT121), .ZN(new_n1180));
  AOI22_X1  g0980(.A1(G107), .A2(new_n753), .B1(new_n759), .B2(new_n372), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n218), .B2(new_n748), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n207), .A2(new_n734), .B1(new_n738), .B2(new_n202), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n591), .B(new_n686), .C1(new_n766), .C2(new_n743), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1180), .A2(new_n1182), .A3(new_n1183), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1185), .A2(KEYINPUT58), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1176), .A2(new_n1178), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n728), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n825), .A2(new_n216), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1168), .A2(new_n788), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1167), .A2(new_n1191), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1193), .B1(new_n1077), .B2(new_n1083), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1103), .B1(new_n1194), .B2(new_n1105), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n1163), .B2(new_n1166), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT57), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1155), .A2(new_n1156), .A3(new_n1137), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n922), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1200));
  OAI211_X1 g1000(.A(KEYINPUT57), .B(new_n1195), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1201), .A2(new_n1002), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1192), .B1(new_n1198), .B2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G375));
  OAI211_X1 g1005(.A(new_n1066), .B(new_n1087), .C1(new_n1100), .C2(new_n1101), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n987), .B(KEYINPUT125), .Z(new_n1207));
  NAND3_X1  g1007(.A1(new_n1104), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n918), .A2(new_n721), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n825), .A2(new_n211), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n953), .A2(new_n738), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(G77), .A2(new_n810), .B1(new_n759), .B2(G107), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n768), .A2(G294), .B1(new_n755), .B2(new_n372), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n744), .A2(G303), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n257), .B1(new_n770), .B2(G97), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n1211), .B(new_n1216), .C1(G283), .C2(new_n753), .ZN(new_n1217));
  AOI22_X1  g1017(.A1(G132), .A2(new_n768), .B1(new_n770), .B2(G159), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1218), .B1(new_n216), .B2(new_n754), .C1(new_n806), .C2(new_n758), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n743), .A2(new_n1109), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1119), .A2(new_n738), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n380), .B1(new_n218), .B2(new_n748), .C1(new_n805), .C2(new_n752), .ZN(new_n1222));
  NOR4_X1   g1022(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .A4(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n728), .B1(new_n1217), .B2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g1024(.A1(new_n1209), .A2(new_n788), .A3(new_n1210), .A4(new_n1224), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n1225), .B1(new_n1194), .B2(new_n1037), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1208), .A2(new_n1227), .ZN(G381));
  NAND2_X1  g1028(.A1(new_n1204), .A2(new_n1135), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT126), .Z(new_n1231));
  OAI211_X1 g1031(.A(new_n1064), .B(new_n973), .C1(new_n988), .C2(new_n999), .ZN(new_n1232));
  OR4_X1    g1032(.A1(G381), .A2(new_n1229), .A3(new_n1231), .A4(new_n1232), .ZN(G407));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(G343), .C2(new_n1229), .ZN(G409));
  AND2_X1   g1034(.A1(G387), .A2(G390), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1232), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(G393), .B(G396), .ZN(new_n1237));
  OR3_X1    g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1237), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n1202), .B1(new_n1197), .B2(new_n1196), .ZN(new_n1242));
  OAI21_X1  g1042(.A(G378), .B1(new_n1242), .B2(new_n1192), .ZN(new_n1243));
  AOI21_X1  g1043(.A(KEYINPUT60), .B1(new_n1194), .B2(new_n1066), .ZN(new_n1244));
  NOR3_X1   g1044(.A1(new_n1244), .A2(new_n1088), .A3(new_n687), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT127), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT60), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1206), .B2(new_n1247), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1194), .A2(KEYINPUT127), .A3(KEYINPUT60), .A4(new_n1066), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1245), .A2(new_n1250), .ZN(new_n1251));
  AOI21_X1  g1051(.A(G384), .B1(new_n1251), .B2(new_n1227), .ZN(new_n1252));
  AOI211_X1 g1052(.A(new_n829), .B(new_n1226), .C1(new_n1245), .C2(new_n1250), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1252), .A2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n669), .A2(G213), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n974), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1256));
  OAI211_X1 g1056(.A(new_n1195), .B(new_n1207), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1135), .A2(new_n1256), .A3(new_n1191), .A4(new_n1257), .ZN(new_n1258));
  NAND4_X1  g1058(.A1(new_n1243), .A2(new_n1254), .A3(new_n1255), .A4(new_n1258), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1259), .A2(KEYINPUT62), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n669), .A2(G213), .A3(G2897), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1262), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1206), .A2(new_n1247), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1002), .A3(new_n1104), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n829), .B1(new_n1266), .B2(new_n1226), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1251), .A2(G384), .A3(new_n1227), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1267), .A2(new_n1268), .A3(new_n1261), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1263), .A2(new_n1269), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1255), .B(new_n1258), .C1(new_n1204), .C2(new_n1135), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1270), .A2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1260), .A2(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT61), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1259), .B2(KEYINPUT62), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1241), .B1(new_n1273), .B2(new_n1275), .ZN(new_n1276));
  AND2_X1   g1076(.A1(new_n1243), .A2(new_n1255), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1277), .A2(KEYINPUT63), .A3(new_n1254), .A4(new_n1258), .ZN(new_n1278));
  AOI21_X1  g1078(.A(KEYINPUT61), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT63), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1259), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1278), .B(new_n1279), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1276), .A2(new_n1283), .ZN(G405));
  NAND2_X1  g1084(.A1(new_n1229), .A2(new_n1243), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1254), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1229), .B(new_n1243), .C1(new_n1252), .C2(new_n1253), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1241), .A2(new_n1286), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1240), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1288), .A2(new_n1290), .ZN(G402));
endmodule


