//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 0 1 1 1 1 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n711, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n192), .A3(new_n195), .A4(new_n190), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT65), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  INV_X1    g015(.A(G146), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G143), .B(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n205), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n194), .A2(KEYINPUT65), .A3(new_n196), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n199), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G116), .ZN(new_n215));
  INV_X1    g029(.A(G116), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(G119), .ZN(new_n217));
  INV_X1    g031(.A(G113), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n218), .A2(KEYINPUT2), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n215), .B(new_n217), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(new_n217), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT2), .B(G113), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT64), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT64), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n222), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G128), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n209), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n200), .A2(KEYINPUT1), .A3(G146), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n231), .B(new_n232), .C1(G128), .C2(new_n209), .ZN(new_n233));
  INV_X1    g047(.A(new_n190), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n188), .A2(G137), .ZN(new_n235));
  OAI21_X1  g049(.A(G131), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n233), .A2(new_n196), .A3(new_n236), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n213), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT28), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n238), .A2(KEYINPUT67), .A3(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(KEYINPUT67), .B1(new_n238), .B2(new_n239), .ZN(new_n242));
  INV_X1    g056(.A(new_n228), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n233), .A2(new_n196), .A3(new_n236), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n194), .A2(new_n196), .B1(new_n208), .B2(new_n210), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n239), .B1(new_n238), .B2(new_n246), .ZN(new_n247));
  NOR3_X1   g061(.A1(new_n241), .A2(new_n242), .A3(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G237), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n252), .A3(G210), .ZN(new_n253));
  XNOR2_X1  g067(.A(new_n253), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n255));
  XNOR2_X1  g069(.A(new_n254), .B(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n242), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n240), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n213), .A2(new_n237), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n243), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n239), .B1(new_n260), .B2(new_n238), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n250), .B(new_n256), .C1(new_n262), .C2(new_n249), .ZN(new_n263));
  INV_X1    g077(.A(G902), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n213), .A2(KEYINPUT30), .A3(new_n237), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n266));
  OAI21_X1  g080(.A(new_n266), .B1(new_n244), .B2(new_n245), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(new_n243), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n238), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(new_n256), .ZN(new_n270));
  INV_X1    g084(.A(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n263), .B(new_n264), .C1(KEYINPUT29), .C2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G472), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n268), .A2(new_n238), .A3(new_n256), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT31), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT31), .ZN(new_n276));
  NAND4_X1  g090(.A1(new_n268), .A2(new_n276), .A3(new_n238), .A4(new_n256), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT66), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n275), .A2(KEYINPUT66), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT68), .ZN(new_n282));
  NOR3_X1   g096(.A1(new_n248), .A2(new_n282), .A3(new_n256), .ZN(new_n283));
  INV_X1    g097(.A(new_n247), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n257), .A2(new_n284), .A3(new_n240), .ZN(new_n285));
  INV_X1    g099(.A(new_n256), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT68), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n280), .B(new_n281), .C1(new_n283), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g103(.A1(G472), .A2(G902), .ZN(new_n290));
  AND3_X1   g104(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n289), .B1(new_n288), .B2(new_n290), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n273), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n273), .B(KEYINPUT69), .C1(new_n291), .C2(new_n292), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT16), .ZN(new_n297));
  INV_X1    g111(.A(G140), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n297), .A2(new_n298), .A3(G125), .ZN(new_n299));
  XOR2_X1   g113(.A(G125), .B(G140), .Z(new_n300));
  OAI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n297), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n202), .ZN(new_n302));
  OAI211_X1 g116(.A(G146), .B(new_n299), .C1(new_n300), .C2(new_n297), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n214), .A2(KEYINPUT70), .A3(G128), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n214), .A2(G128), .ZN(new_n306));
  OAI21_X1  g120(.A(KEYINPUT70), .B1(new_n214), .B2(G128), .ZN(new_n307));
  AOI21_X1  g121(.A(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  XOR2_X1   g122(.A(KEYINPUT24), .B(G110), .Z(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT23), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n311), .B1(new_n214), .B2(G128), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n229), .A2(KEYINPUT23), .A3(G119), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n306), .A3(new_n313), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(KEYINPUT71), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(G110), .A3(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n310), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n318), .B(KEYINPUT72), .ZN(new_n319));
  XOR2_X1   g133(.A(new_n303), .B(KEYINPUT73), .Z(new_n320));
  OAI22_X1  g134(.A1(new_n308), .A2(new_n309), .B1(G110), .B2(new_n314), .ZN(new_n321));
  OR2_X1    g135(.A1(new_n300), .A2(G146), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OR2_X1    g137(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT22), .B(G137), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(new_n324), .A3(new_n328), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n330), .A2(new_n264), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT25), .ZN(new_n333));
  INV_X1    g147(.A(G217), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n334), .B1(G234), .B2(new_n264), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT25), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n336), .A3(new_n264), .A4(new_n331), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n333), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  OR2_X1    g152(.A1(new_n332), .A2(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n295), .A2(new_n296), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT74), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  XOR2_X1   g158(.A(KEYINPUT9), .B(G234), .Z(new_n345));
  NAND3_X1  g159(.A1(new_n345), .A2(G217), .A3(new_n252), .ZN(new_n346));
  INV_X1    g160(.A(G122), .ZN(new_n347));
  OAI21_X1  g161(.A(KEYINPUT83), .B1(new_n347), .B2(G116), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT83), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n349), .A2(new_n216), .A3(G122), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(G116), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(G128), .B(G143), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G134), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n356), .A2(new_n188), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT84), .B1(new_n351), .B2(KEYINPUT14), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n351), .A2(KEYINPUT14), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT84), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT14), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n348), .A2(new_n350), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n362), .A2(new_n353), .A3(new_n363), .A4(new_n366), .ZN(new_n367));
  AOI211_X1 g181(.A(new_n355), .B(new_n361), .C1(new_n367), .C2(G107), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n351), .A2(new_n353), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(G107), .ZN(new_n370));
  AOI22_X1  g184(.A1(new_n370), .A2(new_n354), .B1(new_n188), .B2(new_n356), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n200), .A3(G128), .ZN(new_n373));
  OAI211_X1 g187(.A(G134), .B(new_n373), .C1(new_n357), .C2(new_n372), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n346), .B1(new_n368), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n355), .B1(new_n367), .B2(G107), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n360), .ZN(new_n379));
  INV_X1    g193(.A(new_n346), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n375), .A3(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(G902), .B1(new_n377), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT85), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT15), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(new_n385), .A3(G478), .ZN(new_n386));
  INV_X1    g200(.A(G478), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n382), .B(new_n383), .C1(KEYINPUT15), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(G234), .A2(G237), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(G952), .A3(new_n252), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  XOR2_X1   g207(.A(KEYINPUT21), .B(G898), .Z(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n391), .A2(G902), .A3(G953), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n393), .B1(new_n395), .B2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(G475), .A2(G902), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n251), .A2(new_n252), .A3(G214), .ZN(new_n402));
  NAND2_X1  g216(.A1(KEYINPUT79), .A2(G143), .ZN(new_n403));
  OR2_X1    g217(.A1(KEYINPUT79), .A2(G143), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g219(.A1(KEYINPUT79), .A2(G143), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n406), .A2(G214), .A3(new_n251), .A4(new_n252), .ZN(new_n407));
  AND2_X1   g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(KEYINPUT17), .A3(G131), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(KEYINPUT80), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n408), .A2(G131), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n405), .A2(new_n407), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(new_n195), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n412), .A2(new_n414), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n411), .B1(new_n415), .B2(KEYINPUT17), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT17), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n412), .A2(KEYINPUT81), .A3(new_n417), .A4(new_n414), .ZN(new_n418));
  INV_X1    g232(.A(new_n304), .ZN(new_n419));
  NAND4_X1  g233(.A1(new_n410), .A2(new_n416), .A3(new_n418), .A4(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(G113), .B(G122), .ZN(new_n421));
  INV_X1    g235(.A(G104), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n300), .A2(G146), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n322), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n413), .B1(new_n426), .B2(new_n195), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n425), .B(new_n427), .C1(new_n412), .C2(new_n426), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n420), .A2(new_n423), .A3(new_n428), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n300), .B(KEYINPUT19), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n415), .B1(G146), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n428), .B1(new_n431), .B2(new_n320), .ZN(new_n432));
  INV_X1    g246(.A(new_n423), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n435), .A2(KEYINPUT82), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT82), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(new_n429), .B2(new_n434), .ZN(new_n438));
  OAI211_X1 g252(.A(KEYINPUT20), .B(new_n401), .C1(new_n436), .C2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n401), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT20), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n429), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n423), .B1(new_n420), .B2(new_n428), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n264), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G475), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n439), .A2(new_n442), .A3(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n400), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(G214), .B1(G237), .B2(G902), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(KEYINPUT3), .B1(new_n422), .B2(G107), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT3), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n452), .A2(new_n352), .A3(G104), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n422), .A2(G107), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n453), .A3(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(G101), .ZN(new_n456));
  INV_X1    g270(.A(G101), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n451), .A2(new_n453), .A3(new_n457), .A4(new_n454), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(KEYINPUT4), .A3(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT4), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n455), .A2(new_n460), .A3(G101), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n459), .A2(new_n225), .A3(new_n227), .A4(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n352), .A2(G104), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n422), .A2(G107), .ZN(new_n464));
  OAI21_X1  g278(.A(G101), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g279(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT5), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(G113), .C1(KEYINPUT5), .C2(new_n215), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n466), .A2(new_n221), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n462), .A2(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(G110), .B(G122), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT77), .Z(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(new_n472), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n462), .A2(new_n469), .A3(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n473), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n462), .B2(new_n469), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT6), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(KEYINPUT78), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n211), .A2(G125), .ZN(new_n482));
  AND3_X1   g296(.A1(new_n230), .A2(new_n201), .A3(new_n203), .ZN(new_n483));
  AOI21_X1  g297(.A(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n484));
  INV_X1    g298(.A(new_n232), .ZN(new_n485));
  NOR3_X1   g299(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n482), .B1(G125), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n252), .A2(G224), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT78), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n476), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n481), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n488), .A2(KEYINPUT7), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n487), .B(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n468), .A2(new_n221), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n495), .B(new_n466), .ZN(new_n496));
  XNOR2_X1  g310(.A(new_n472), .B(KEYINPUT8), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n494), .B(new_n475), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n492), .A2(new_n264), .A3(new_n498), .ZN(new_n499));
  OAI21_X1  g313(.A(G210), .B1(G237), .B2(G902), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n490), .B1(new_n476), .B2(new_n479), .ZN(new_n503));
  AND3_X1   g317(.A1(new_n462), .A2(new_n469), .A3(new_n474), .ZN(new_n504));
  NOR2_X1   g318(.A1(new_n504), .A2(new_n477), .ZN(new_n505));
  AOI21_X1  g319(.A(KEYINPUT78), .B1(new_n505), .B2(KEYINPUT6), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(G902), .B1(new_n507), .B2(new_n489), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n500), .A3(new_n498), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n450), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n448), .A2(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n459), .A2(new_n461), .A3(new_n211), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT10), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n458), .A2(new_n465), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n486), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n233), .A2(new_n466), .A3(KEYINPUT10), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n199), .A2(new_n212), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n518), .A2(new_n519), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(KEYINPUT75), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT75), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n518), .A2(new_n523), .A3(new_n519), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n520), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  XNOR2_X1  g339(.A(G110), .B(G140), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n252), .A2(G227), .ZN(new_n527));
  XNOR2_X1  g341(.A(new_n526), .B(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT76), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n520), .ZN(new_n530));
  INV_X1    g344(.A(new_n524), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n523), .B1(new_n518), .B2(new_n519), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT76), .ZN(new_n534));
  INV_X1    g348(.A(new_n528), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n533), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n486), .B(new_n515), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(KEYINPUT12), .A3(new_n197), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n519), .A2(new_n537), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n538), .B1(new_n539), .B2(KEYINPUT12), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n520), .A2(new_n535), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n529), .A2(new_n536), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G469), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(new_n544), .A3(new_n264), .ZN(new_n545));
  NAND2_X1  g359(.A1(G469), .A2(G902), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n541), .B1(new_n531), .B2(new_n532), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n540), .A2(new_n530), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n528), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n545), .B(new_n546), .C1(new_n544), .C2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(G221), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n551), .B1(new_n345), .B2(new_n264), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g369(.A1(new_n295), .A2(KEYINPUT74), .A3(new_n296), .A4(new_n341), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n344), .A2(new_n512), .A3(new_n555), .A4(new_n556), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT86), .B(G101), .Z(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(G3));
  NAND2_X1  g373(.A1(new_n381), .A2(KEYINPUT88), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n346), .A2(KEYINPUT88), .ZN(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(KEYINPUT87), .B(new_n562), .C1(new_n368), .C2(new_n376), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n378), .A2(new_n360), .B1(new_n374), .B2(new_n371), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT87), .ZN(new_n565));
  OAI21_X1  g379(.A(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n560), .A2(new_n563), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT33), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT33), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n377), .A2(new_n569), .A3(new_n381), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(G478), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n387), .A2(new_n264), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n382), .A2(new_n387), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n571), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT89), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n571), .A2(new_n577), .A3(new_n573), .A4(new_n574), .ZN(new_n578));
  AND3_X1   g392(.A1(new_n576), .A2(new_n447), .A3(new_n578), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n450), .B(new_n398), .C1(new_n502), .C2(new_n509), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(KEYINPUT90), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n341), .A2(new_n550), .A3(new_n553), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n288), .A2(new_n290), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n282), .B1(new_n248), .B2(new_n256), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n285), .A2(KEYINPUT68), .A3(new_n286), .ZN(new_n586));
  AOI22_X1  g400(.A1(new_n585), .A2(new_n586), .B1(KEYINPUT66), .B2(new_n275), .ZN(new_n587));
  AOI21_X1  g401(.A(G902), .B1(new_n587), .B2(new_n280), .ZN(new_n588));
  INV_X1    g402(.A(G472), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n582), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(new_n592), .B(new_n422), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT91), .B(KEYINPUT34), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  OAI21_X1  g409(.A(new_n401), .B1(new_n436), .B2(new_n438), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(new_n441), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n439), .A2(new_n389), .A3(new_n446), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n580), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n599), .A2(new_n590), .A3(new_n583), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n600), .B(new_n352), .ZN(new_n601));
  XNOR2_X1  g415(.A(KEYINPUT92), .B(KEYINPUT35), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G9));
  NOR2_X1   g417(.A1(new_n329), .A2(KEYINPUT36), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT93), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n325), .B(new_n605), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n606), .B(new_n264), .C1(new_n334), .C2(G234), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n338), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n550), .A2(new_n553), .A3(new_n608), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n511), .A2(new_n590), .A3(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT37), .B(G110), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G12));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n393), .B1(new_n397), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n596), .B2(new_n441), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n295), .A2(new_n296), .A3(new_n598), .A4(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n609), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(new_n510), .ZN(new_n618));
  OR2_X1    g432(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(G128), .ZN(G30));
  XNOR2_X1  g434(.A(new_n614), .B(KEYINPUT39), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n555), .A2(new_n622), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(KEYINPUT40), .ZN(new_n624));
  OR3_X1    g438(.A1(new_n624), .A2(new_n450), .A3(new_n608), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n502), .A2(new_n509), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n626), .B(KEYINPUT38), .Z(new_n627));
  NAND2_X1  g441(.A1(new_n447), .A2(new_n389), .ZN(new_n628));
  AND2_X1   g442(.A1(new_n260), .A2(new_n238), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n264), .B1(new_n630), .B2(new_n256), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n269), .A2(new_n256), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(G472), .B1(new_n631), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n634), .B1(new_n291), .B2(new_n292), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT94), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NOR4_X1   g451(.A1(new_n625), .A2(new_n627), .A3(new_n628), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(new_n200), .ZN(G45));
  AND2_X1   g453(.A1(new_n295), .A2(new_n296), .ZN(new_n640));
  INV_X1    g454(.A(new_n614), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n579), .A2(KEYINPUT95), .A3(new_n510), .A4(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n579), .A2(new_n510), .A3(new_n641), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT95), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n554), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n640), .A2(new_n608), .A3(new_n642), .A4(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G146), .ZN(G48));
  INV_X1    g461(.A(new_n545), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n544), .B1(new_n543), .B2(new_n264), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(KEYINPUT96), .A3(new_n553), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n543), .A2(new_n264), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(G469), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n653), .A2(new_n553), .A3(new_n545), .ZN(new_n654));
  INV_X1    g468(.A(KEYINPUT96), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n651), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n295), .A2(new_n296), .A3(new_n657), .A4(new_n341), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n582), .ZN(new_n660));
  XNOR2_X1  g474(.A(KEYINPUT41), .B(G113), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n660), .B(new_n661), .ZN(G15));
  NOR2_X1   g476(.A1(new_n658), .A2(new_n599), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(new_n216), .ZN(G18));
  AOI21_X1  g478(.A(new_n500), .B1(new_n508), .B2(new_n498), .ZN(new_n665));
  AND4_X1   g479(.A1(new_n264), .A2(new_n492), .A3(new_n500), .A4(new_n498), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n449), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT97), .B1(new_n654), .B2(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(KEYINPUT97), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n650), .A2(new_n510), .A3(new_n669), .A4(new_n553), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n295), .A3(new_n296), .A4(new_n608), .ZN(new_n672));
  INV_X1    g486(.A(new_n448), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n214), .ZN(G21));
  AOI21_X1  g489(.A(new_n628), .B1(new_n651), .B2(new_n656), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n589), .B1(new_n288), .B2(new_n264), .ZN(new_n677));
  INV_X1    g491(.A(new_n278), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n286), .B1(new_n258), .B2(new_n261), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n290), .B(KEYINPUT98), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n677), .A2(new_n683), .ZN(new_n684));
  AOI21_X1  g498(.A(KEYINPUT99), .B1(new_n684), .B2(new_n341), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT99), .ZN(new_n686));
  NOR4_X1   g500(.A1(new_n677), .A2(new_n340), .A3(new_n683), .A4(new_n686), .ZN(new_n687));
  OAI211_X1 g501(.A(new_n676), .B(new_n580), .C1(new_n685), .C2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G122), .ZN(G24));
  OAI211_X1 g503(.A(new_n608), .B(new_n682), .C1(new_n588), .C2(new_n589), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n576), .A2(new_n447), .A3(new_n578), .A4(new_n641), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n671), .A2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n671), .A2(new_n692), .A3(KEYINPUT100), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(G125), .ZN(G27));
  NAND3_X1  g512(.A1(new_n502), .A2(new_n509), .A3(new_n449), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n554), .A2(new_n691), .A3(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n640), .A2(KEYINPUT101), .A3(new_n341), .A4(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n700), .A2(new_n295), .A3(new_n296), .A4(new_n341), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT101), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n702), .A3(new_n705), .ZN(new_n706));
  AND2_X1   g520(.A1(new_n293), .A2(new_n341), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(KEYINPUT42), .A3(new_n700), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G131), .ZN(G33));
  NOR3_X1   g524(.A1(new_n616), .A2(new_n583), .A3(new_n699), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(new_n188), .ZN(G36));
  XNOR2_X1  g526(.A(new_n699), .B(KEYINPUT103), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n549), .B(KEYINPUT45), .ZN(new_n714));
  OAI21_X1  g528(.A(G469), .B1(new_n714), .B2(G902), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(KEYINPUT46), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(new_n545), .A3(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n553), .A3(new_n622), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n576), .A2(new_n578), .ZN(new_n720));
  INV_X1    g534(.A(new_n447), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT43), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT43), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT102), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n724), .A2(KEYINPUT102), .A3(new_n726), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n729), .A2(new_n590), .A3(new_n608), .A4(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n719), .B1(new_n731), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n732), .A2(KEYINPUT44), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g550(.A(new_n713), .B(new_n734), .C1(new_n736), .C2(new_n733), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G137), .ZN(G39));
  NAND2_X1  g552(.A1(new_n718), .A2(new_n553), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n739), .B(KEYINPUT47), .Z(new_n740));
  INV_X1    g554(.A(new_n640), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n691), .A2(new_n341), .A3(new_n699), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G140), .ZN(G42));
  AND3_X1   g558(.A1(new_n671), .A2(KEYINPUT100), .A3(new_n692), .ZN(new_n745));
  AOI21_X1  g559(.A(KEYINPUT100), .B1(new_n671), .B2(new_n692), .ZN(new_n746));
  OAI22_X1  g560(.A1(new_n745), .A2(new_n746), .B1(new_n616), .B2(new_n618), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT107), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  OAI221_X1 g563(.A(new_n749), .B1(new_n616), .B2(new_n618), .C1(new_n745), .C2(new_n746), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n554), .A2(new_n608), .A3(new_n614), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n628), .A2(new_n667), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n751), .A2(new_n635), .A3(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT52), .ZN(new_n755));
  NOR2_X1   g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n748), .A2(new_n750), .A3(new_n646), .A4(new_n756), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n619), .A2(new_n646), .A3(new_n697), .A4(new_n753), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT108), .ZN(new_n761));
  INV_X1    g575(.A(new_n711), .ZN(new_n762));
  AND3_X1   g576(.A1(new_n295), .A2(new_n296), .A3(new_n615), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n699), .A2(new_n389), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n439), .A2(new_n446), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n763), .A2(KEYINPUT106), .A3(new_n617), .A4(new_n766), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n295), .A2(new_n617), .A3(new_n296), .A4(new_n615), .ZN(new_n769));
  INV_X1    g583(.A(new_n766), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n768), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n709), .A2(new_n762), .A3(new_n772), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n510), .A2(new_n598), .A3(new_n442), .A4(new_n399), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT105), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n580), .A2(KEYINPUT105), .A3(new_n442), .A4(new_n598), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(new_n777), .A3(new_n581), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n591), .ZN(new_n779));
  INV_X1    g593(.A(new_n610), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n779), .A2(new_n688), .A3(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n781), .A2(new_n674), .A3(new_n663), .ZN(new_n782));
  INV_X1    g596(.A(new_n690), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n700), .A2(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n782), .A2(new_n557), .A3(new_n660), .A4(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n773), .A2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT108), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n757), .A2(new_n759), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n761), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(KEYINPUT53), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n791));
  AOI221_X4 g605(.A(new_n711), .B1(new_n767), .B2(new_n771), .C1(new_n706), .C2(new_n708), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n557), .A2(new_n660), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n658), .A2(new_n599), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n640), .A2(new_n448), .A3(new_n608), .A4(new_n671), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n610), .B1(new_n778), .B2(new_n591), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n794), .A2(new_n795), .A3(new_n688), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n784), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n793), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n619), .A2(new_n646), .A3(new_n697), .A4(new_n756), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n295), .A2(new_n642), .A3(new_n296), .A4(new_n608), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n643), .A2(new_n644), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n801), .A2(new_n802), .A3(new_n554), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n747), .A2(new_n803), .A3(new_n754), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n800), .B1(new_n804), .B2(KEYINPUT52), .ZN(new_n805));
  AND4_X1   g619(.A1(new_n791), .A2(new_n792), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(KEYINPUT54), .B1(new_n790), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n786), .A2(KEYINPUT53), .A3(new_n805), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT109), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n789), .A2(new_n791), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n808), .B1(new_n814), .B2(KEYINPUT54), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n392), .B1(new_n724), .B2(new_n726), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n816), .B1(new_n685), .B2(new_n687), .ZN(new_n817));
  INV_X1    g631(.A(new_n817), .ZN(new_n818));
  INV_X1    g632(.A(new_n654), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n818), .A2(new_n450), .A3(new_n627), .A4(new_n819), .ZN(new_n820));
  NOR2_X1   g634(.A1(KEYINPUT110), .A2(KEYINPUT50), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n648), .A2(new_n649), .A3(new_n553), .ZN(new_n823));
  OR2_X1    g637(.A1(new_n740), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n713), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n654), .A2(new_n699), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n637), .A2(new_n393), .A3(new_n341), .A4(new_n828), .ZN(new_n829));
  OR3_X1    g643(.A1(new_n829), .A2(new_n447), .A3(new_n720), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n816), .A2(new_n783), .A3(new_n828), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n822), .A2(new_n827), .A3(new_n830), .A4(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT111), .B1(new_n824), .B2(new_n826), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n833), .A2(KEYINPUT51), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n832), .A2(new_n834), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n818), .A2(new_n671), .ZN(new_n837));
  XOR2_X1   g651(.A(new_n837), .B(KEYINPUT112), .Z(new_n838));
  NAND3_X1  g652(.A1(new_n816), .A2(new_n707), .A3(new_n828), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n839), .B(KEYINPUT48), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n838), .A2(G952), .A3(new_n252), .A4(new_n840), .ZN(new_n841));
  NOR3_X1   g655(.A1(new_n835), .A2(new_n836), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(new_n579), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n815), .B(new_n842), .C1(new_n843), .C2(new_n829), .ZN(new_n844));
  INV_X1    g658(.A(G952), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n845), .A2(new_n252), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT113), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n844), .A2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n627), .A2(new_n449), .A3(new_n341), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n650), .B(KEYINPUT49), .Z(new_n850));
  NOR3_X1   g664(.A1(new_n849), .A2(new_n552), .A3(new_n850), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n851), .A2(new_n637), .A3(new_n723), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n848), .A2(new_n852), .ZN(G75));
  XNOR2_X1  g667(.A(new_n507), .B(new_n489), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT114), .ZN(new_n855));
  XNOR2_X1  g669(.A(new_n855), .B(KEYINPUT55), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n806), .B1(new_n789), .B2(KEYINPUT53), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(G210), .A3(G902), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT56), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n858), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n859), .B1(new_n858), .B2(new_n860), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n856), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OR2_X1    g677(.A1(new_n862), .A2(new_n856), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n845), .A2(G953), .ZN(new_n865));
  XOR2_X1   g679(.A(new_n865), .B(KEYINPUT116), .Z(new_n866));
  XOR2_X1   g680(.A(new_n866), .B(KEYINPUT117), .Z(new_n867));
  AND3_X1   g681(.A1(new_n863), .A2(new_n864), .A3(new_n867), .ZN(G51));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n869));
  XOR2_X1   g683(.A(new_n546), .B(KEYINPUT57), .Z(new_n870));
  INV_X1    g684(.A(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  AND3_X1   g686(.A1(new_n757), .A2(new_n787), .A3(new_n759), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n787), .B1(new_n757), .B2(new_n759), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n791), .B1(new_n875), .B2(new_n786), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n872), .B1(new_n876), .B2(new_n806), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n857), .A2(KEYINPUT54), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n871), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  XNOR2_X1  g693(.A(new_n543), .B(KEYINPUT118), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n869), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AOI211_X1 g695(.A(new_n872), .B(new_n806), .C1(KEYINPUT53), .C2(new_n789), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n870), .B1(new_n882), .B2(new_n808), .ZN(new_n883));
  INV_X1    g697(.A(new_n880), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(KEYINPUT119), .A3(new_n884), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n714), .A2(G469), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n857), .A2(G902), .A3(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT120), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n887), .B(new_n888), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n881), .A2(new_n885), .A3(new_n889), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n890), .A2(new_n866), .ZN(G54));
  NAND4_X1  g705(.A1(new_n857), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n436), .A2(new_n438), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n892), .B(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n866), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(G60));
  NAND2_X1  g710(.A1(new_n568), .A2(new_n570), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n897), .B(KEYINPUT121), .ZN(new_n898));
  XNOR2_X1  g712(.A(new_n572), .B(KEYINPUT59), .ZN(new_n899));
  INV_X1    g713(.A(new_n899), .ZN(new_n900));
  OAI211_X1 g714(.A(new_n898), .B(new_n900), .C1(new_n882), .C2(new_n808), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n815), .A2(new_n899), .ZN(new_n902));
  OAI211_X1 g716(.A(new_n867), .B(new_n901), .C1(new_n902), .C2(new_n898), .ZN(new_n903));
  INV_X1    g717(.A(new_n903), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT123), .ZN(new_n906));
  XOR2_X1   g720(.A(KEYINPUT122), .B(KEYINPUT60), .Z(new_n907));
  XNOR2_X1  g721(.A(new_n906), .B(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n876), .A2(new_n806), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n606), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n330), .A2(new_n331), .ZN(new_n911));
  OAI211_X1 g725(.A(new_n910), .B(new_n867), .C1(new_n911), .C2(new_n909), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT61), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(G66));
  INV_X1    g728(.A(G224), .ZN(new_n915));
  OAI21_X1  g729(.A(G953), .B1(new_n395), .B2(new_n915), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n793), .A2(new_n797), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(G953), .ZN(new_n918));
  OAI22_X1  g732(.A1(new_n503), .A2(new_n506), .B1(G898), .B2(new_n252), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G69));
  NAND2_X1  g734(.A1(new_n737), .A2(new_n743), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n748), .A2(new_n750), .A3(new_n646), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n707), .ZN(new_n924));
  NOR4_X1   g738(.A1(new_n719), .A2(new_n924), .A3(new_n667), .A4(new_n628), .ZN(new_n925));
  AOI211_X1 g739(.A(new_n711), .B(new_n925), .C1(new_n706), .C2(new_n708), .ZN(new_n926));
  AOI21_X1  g740(.A(G953), .B1(new_n923), .B2(new_n926), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n252), .A2(G900), .ZN(new_n928));
  OR3_X1    g742(.A1(new_n927), .A2(KEYINPUT125), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n265), .A2(new_n267), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(new_n430), .Z(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(KEYINPUT125), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n929), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n344), .A2(new_n556), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n843), .B1(new_n447), .B2(new_n390), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n699), .A2(new_n621), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n935), .A2(new_n555), .A3(new_n936), .A4(new_n937), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT124), .Z(new_n939));
  INV_X1    g753(.A(new_n921), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n638), .A2(new_n922), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT62), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n941), .A2(new_n942), .ZN(new_n944));
  OAI211_X1 g758(.A(new_n939), .B(new_n940), .C1(new_n943), .C2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(new_n252), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(new_n931), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n252), .B1(G227), .B2(G900), .ZN(new_n948));
  AND3_X1   g762(.A1(new_n934), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n948), .B1(new_n934), .B2(new_n947), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(G72));
  XNOR2_X1  g765(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n589), .A2(new_n264), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n952), .B(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n917), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n954), .B1(new_n945), .B2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n895), .B1(new_n956), .B2(new_n633), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n923), .A2(new_n917), .A3(new_n926), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n954), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n270), .B(KEYINPUT127), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n814), .A2(new_n271), .A3(new_n632), .A4(new_n954), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n957), .A2(new_n961), .A3(new_n962), .ZN(G57));
endmodule


