//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n728, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966;
  INV_X1    g000(.A(KEYINPUT92), .ZN(new_n187));
  OAI21_X1  g001(.A(G210), .B1(G237), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G146), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G146), .ZN(new_n193));
  AND2_X1   g007(.A1(KEYINPUT0), .A2(G128), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n191), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(G143), .B(G146), .ZN(new_n196));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G128), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n195), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT64), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(new_n193), .ZN(new_n200));
  NOR2_X1   g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n194), .A2(new_n201), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n200), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(new_n204), .ZN(new_n205));
  AOI21_X1  g019(.A(KEYINPUT82), .B1(new_n205), .B2(G125), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n207));
  INV_X1    g021(.A(G125), .ZN(new_n208));
  AOI211_X1 g022(.A(new_n207), .B(new_n208), .C1(new_n199), .C2(new_n204), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT83), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n205), .A2(KEYINPUT82), .A3(G125), .ZN(new_n211));
  AOI21_X1  g025(.A(new_n203), .B1(KEYINPUT64), .B2(new_n198), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n207), .B1(new_n212), .B2(new_n208), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT83), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n211), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G128), .ZN(new_n216));
  OAI211_X1 g030(.A(new_n192), .B(G146), .C1(new_n216), .C2(KEYINPUT1), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n216), .A2(new_n190), .A3(G143), .ZN(new_n218));
  AND2_X1   g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT1), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n196), .A2(new_n220), .A3(G128), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n221), .A3(new_n208), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n210), .A2(new_n215), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G953), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G224), .ZN(new_n225));
  XNOR2_X1  g039(.A(new_n225), .B(KEYINPUT84), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n223), .A2(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(new_n226), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n210), .A2(new_n228), .A3(new_n215), .A4(new_n222), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(G104), .ZN(new_n231));
  OAI21_X1  g045(.A(KEYINPUT3), .B1(new_n231), .B2(G107), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT3), .ZN(new_n233));
  INV_X1    g047(.A(G107), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n233), .A2(new_n234), .A3(G104), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(G107), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n232), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(G101), .ZN(new_n238));
  INV_X1    g052(.A(G101), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n232), .A2(new_n235), .A3(new_n239), .A4(new_n236), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n238), .A2(KEYINPUT4), .A3(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G119), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G116), .ZN(new_n243));
  INV_X1    g057(.A(G116), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G119), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT2), .B(G113), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n246), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n237), .A2(new_n249), .A3(G101), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n241), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT80), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n246), .A2(new_n247), .ZN(new_n253));
  XNOR2_X1  g067(.A(G116), .B(G119), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT5), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n243), .A2(KEYINPUT5), .ZN(new_n256));
  INV_X1    g070(.A(G113), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n253), .B1(new_n255), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT75), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n260), .A2(new_n234), .A3(G104), .ZN(new_n261));
  OAI21_X1  g075(.A(KEYINPUT75), .B1(new_n234), .B2(G104), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n231), .A2(G107), .ZN(new_n263));
  OAI211_X1 g077(.A(G101), .B(new_n261), .C1(new_n262), .C2(new_n263), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(new_n240), .A3(KEYINPUT77), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT77), .B1(new_n264), .B2(new_n240), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n259), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT80), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n241), .A2(new_n248), .A3(new_n269), .A4(new_n250), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n252), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  XOR2_X1   g085(.A(G110), .B(G122), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n252), .A2(new_n274), .A3(new_n268), .A4(new_n270), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n271), .A2(new_n277), .A3(new_n272), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(KEYINPUT81), .A3(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT81), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n273), .A2(new_n280), .A3(KEYINPUT6), .A4(new_n275), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n230), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n226), .A2(KEYINPUT7), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT86), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n222), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n213), .A3(new_n211), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n255), .A2(KEYINPUT85), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n254), .A2(new_n288), .A3(KEYINPUT5), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n258), .A3(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n290), .B1(new_n246), .B2(new_n247), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n266), .A2(new_n267), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n264), .A2(new_n240), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI22_X1  g108(.A1(new_n291), .A2(new_n292), .B1(new_n294), .B2(new_n259), .ZN(new_n295));
  XOR2_X1   g109(.A(new_n272), .B(KEYINPUT8), .Z(new_n296));
  AOI22_X1  g110(.A1(new_n283), .A2(new_n286), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n297), .B(new_n275), .C1(new_n223), .C2(new_n283), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n189), .B1(new_n282), .B2(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n273), .A2(KEYINPUT6), .A3(new_n275), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n278), .A2(KEYINPUT81), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n281), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n227), .A2(new_n229), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n298), .A2(new_n299), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n306), .A2(new_n307), .A3(new_n188), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n301), .A2(new_n308), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n224), .A2(G952), .ZN(new_n310));
  NAND2_X1  g124(.A1(G234), .A2(G237), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  XOR2_X1   g127(.A(KEYINPUT21), .B(G898), .Z(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n311), .A2(G902), .A3(G953), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n313), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(G214), .B1(G237), .B2(G902), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n309), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G475), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n299), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n323), .B(KEYINPUT89), .ZN(new_n324));
  NOR2_X1   g138(.A1(G237), .A2(G953), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(G143), .A3(G214), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(G143), .B1(new_n325), .B2(G214), .ZN(new_n328));
  NOR2_X1   g142(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT88), .ZN(new_n330));
  INV_X1    g144(.A(G131), .ZN(new_n331));
  NOR3_X1   g145(.A1(new_n329), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n328), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(new_n326), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT88), .B1(new_n334), .B2(G131), .ZN(new_n335));
  OAI21_X1  g149(.A(KEYINPUT17), .B1(new_n332), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n330), .B1(new_n329), .B2(new_n331), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n334), .A2(KEYINPUT88), .A3(G131), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT17), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n329), .A2(new_n331), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n337), .A2(new_n338), .A3(new_n339), .A4(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT16), .ZN(new_n342));
  INV_X1    g156(.A(G140), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n342), .A2(new_n343), .A3(G125), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n208), .A2(G140), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n343), .A2(G125), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(KEYINPUT71), .ZN(new_n347));
  OR3_X1    g161(.A1(new_n343), .A2(KEYINPUT71), .A3(G125), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n344), .B1(new_n350), .B2(new_n342), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n190), .ZN(new_n352));
  OAI211_X1 g166(.A(G146), .B(new_n344), .C1(new_n350), .C2(new_n342), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n336), .A2(new_n341), .A3(new_n352), .A4(new_n353), .ZN(new_n354));
  AND2_X1   g168(.A1(new_n345), .A2(new_n346), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(new_n190), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AND3_X1   g171(.A1(new_n347), .A2(KEYINPUT87), .A3(new_n348), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT87), .B1(new_n347), .B2(new_n348), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n357), .B1(new_n360), .B2(new_n190), .ZN(new_n361));
  NAND2_X1  g175(.A1(KEYINPUT18), .A2(G131), .ZN(new_n362));
  XNOR2_X1  g176(.A(new_n334), .B(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G113), .B(G122), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(new_n231), .ZN(new_n366));
  AND3_X1   g180(.A1(new_n354), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n337), .A2(new_n338), .A3(new_n340), .ZN(new_n368));
  OAI21_X1  g182(.A(KEYINPUT19), .B1(new_n358), .B2(new_n359), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT19), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n355), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  OAI211_X1 g186(.A(new_n353), .B(new_n368), .C1(new_n372), .C2(G146), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n366), .B1(new_n373), .B2(new_n364), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n324), .B1(new_n367), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT20), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n366), .B1(new_n354), .B2(new_n364), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n299), .B1(new_n367), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G475), .ZN(new_n380));
  OAI211_X1 g194(.A(KEYINPUT20), .B(new_n324), .C1(new_n367), .C2(new_n374), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n377), .A2(new_n380), .A3(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(KEYINPUT9), .B(G234), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n383), .B(KEYINPUT73), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(G217), .A3(new_n224), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G116), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n244), .A2(G122), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n387), .A2(new_n388), .A3(new_n234), .ZN(new_n389));
  XNOR2_X1  g203(.A(G128), .B(G143), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n390), .B(G134), .ZN(new_n391));
  OAI21_X1  g205(.A(KEYINPUT14), .B1(new_n386), .B2(G116), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT90), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT90), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n388), .A2(new_n394), .A3(KEYINPUT14), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(new_n387), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT91), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n388), .A2(KEYINPUT14), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n393), .A2(new_n395), .A3(KEYINPUT91), .A4(new_n387), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI211_X1 g215(.A(new_n389), .B(new_n391), .C1(new_n401), .C2(G107), .ZN(new_n402));
  INV_X1    g216(.A(G134), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n216), .A2(KEYINPUT13), .A3(G143), .ZN(new_n404));
  AOI211_X1 g218(.A(new_n403), .B(new_n404), .C1(KEYINPUT13), .C2(new_n390), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n390), .A2(new_n403), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n234), .B1(new_n387), .B2(new_n388), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n406), .B1(new_n389), .B2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n385), .B1(new_n402), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n401), .A2(G107), .ZN(new_n411));
  INV_X1    g225(.A(new_n389), .ZN(new_n412));
  INV_X1    g226(.A(new_n391), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n409), .ZN(new_n415));
  INV_X1    g229(.A(new_n385), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(G902), .B1(new_n410), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G478), .ZN(new_n419));
  OR2_X1    g233(.A1(new_n419), .A2(KEYINPUT15), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n418), .B(new_n420), .ZN(new_n421));
  NOR2_X1   g235(.A1(new_n382), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(G469), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n221), .A2(KEYINPUT76), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT76), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n196), .A2(new_n425), .A3(new_n220), .A4(G128), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n424), .A2(new_n219), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n294), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT10), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT65), .A2(G137), .ZN(new_n431));
  NOR2_X1   g245(.A1(KEYINPUT65), .A2(G137), .ZN(new_n432));
  OAI211_X1 g246(.A(KEYINPUT11), .B(G134), .C1(new_n431), .C2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(G137), .ZN(new_n434));
  OAI21_X1  g248(.A(KEYINPUT11), .B1(new_n434), .B2(G134), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(G134), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(G131), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n433), .A2(new_n437), .A3(new_n331), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n219), .A2(new_n221), .ZN(new_n443));
  OAI211_X1 g257(.A(KEYINPUT10), .B(new_n443), .C1(new_n266), .C2(new_n267), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n212), .A2(new_n250), .A3(new_n241), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n430), .A2(new_n442), .A3(new_n444), .A4(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(G110), .B(G140), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n447), .B(KEYINPUT74), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n224), .A2(G227), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n448), .B(new_n449), .Z(new_n450));
  NAND2_X1  g264(.A1(new_n446), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT77), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n293), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n443), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n453), .A2(new_n454), .A3(new_n265), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT78), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n453), .A2(new_n454), .A3(new_n457), .A4(new_n265), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n456), .A2(new_n428), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n441), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT12), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(KEYINPUT12), .A3(new_n441), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n451), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n430), .A2(new_n445), .A3(new_n444), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n441), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n450), .B1(new_n466), .B2(new_n446), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n423), .B(new_n299), .C1(new_n464), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT79), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n451), .A2(new_n469), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n446), .A2(KEYINPUT79), .A3(new_n450), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n466), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n446), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n473), .B1(new_n462), .B2(new_n463), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n472), .B(G469), .C1(new_n474), .C2(new_n450), .ZN(new_n475));
  NAND2_X1  g289(.A1(G469), .A2(G902), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n468), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(new_n384), .ZN(new_n478));
  OAI21_X1  g292(.A(G221), .B1(new_n478), .B2(G902), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n422), .A2(new_n477), .A3(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n187), .B1(new_n321), .B2(new_n480), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n422), .A2(new_n477), .A3(new_n479), .ZN(new_n482));
  INV_X1    g296(.A(new_n320), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n483), .B1(new_n301), .B2(new_n308), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n482), .A2(KEYINPUT92), .A3(new_n319), .A4(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(KEYINPUT69), .B(KEYINPUT28), .ZN(new_n486));
  INV_X1    g300(.A(new_n248), .ZN(new_n487));
  NOR3_X1   g301(.A1(new_n431), .A2(new_n432), .A3(G134), .ZN(new_n488));
  INV_X1    g302(.A(new_n436), .ZN(new_n489));
  OAI21_X1  g303(.A(G131), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n443), .A2(new_n440), .A3(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n441), .A2(new_n212), .A3(KEYINPUT66), .ZN(new_n492));
  AOI21_X1  g306(.A(KEYINPUT66), .B1(new_n441), .B2(new_n212), .ZN(new_n493));
  OAI211_X1 g307(.A(new_n487), .B(new_n491), .C1(new_n492), .C2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n441), .A2(new_n212), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n491), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n496), .A2(new_n248), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n486), .B1(new_n494), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT28), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n496), .B2(new_n248), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(G101), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n325), .A2(G210), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT68), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n494), .A2(new_n509), .A3(new_n506), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n509), .B1(new_n494), .B2(new_n506), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT30), .ZN(new_n513));
  AOI21_X1  g327(.A(KEYINPUT67), .B1(new_n496), .B2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n515));
  OAI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(new_n513), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT66), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n495), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n441), .A2(new_n212), .A3(KEYINPUT66), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g334(.A1(new_n520), .A2(KEYINPUT67), .A3(KEYINPUT30), .A4(new_n491), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n487), .B1(new_n516), .B2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT31), .ZN(new_n523));
  NOR3_X1   g337(.A1(new_n512), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n516), .A2(new_n521), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n248), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n494), .A2(new_n506), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT68), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n494), .A2(new_n509), .A3(new_n506), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT31), .B1(new_n526), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n508), .B1(new_n524), .B2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(G472), .A2(G902), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n532), .A2(KEYINPUT32), .A3(new_n533), .ZN(new_n534));
  XOR2_X1   g348(.A(KEYINPUT70), .B(KEYINPUT32), .Z(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n523), .B1(new_n512), .B2(new_n522), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n526), .A2(KEYINPUT31), .A3(new_n530), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n507), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n533), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n515), .A2(new_n248), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n499), .B1(new_n542), .B2(new_n494), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  NAND4_X1  g358(.A1(new_n544), .A2(KEYINPUT29), .A3(new_n506), .A4(new_n500), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n506), .B1(new_n526), .B2(new_n494), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT29), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n494), .A2(new_n497), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n500), .B1(new_n548), .B2(new_n486), .ZN(new_n549));
  INV_X1    g363(.A(new_n506), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n547), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n299), .B(new_n545), .C1(new_n546), .C2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(G472), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n534), .A2(new_n541), .A3(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n352), .A2(new_n353), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT23), .B1(new_n242), .B2(G128), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NOR3_X1   g371(.A1(new_n242), .A2(KEYINPUT23), .A3(G128), .ZN(new_n558));
  OAI22_X1  g372(.A1(new_n557), .A2(new_n558), .B1(G119), .B2(new_n216), .ZN(new_n559));
  XNOR2_X1  g373(.A(G119), .B(G128), .ZN(new_n560));
  XOR2_X1   g374(.A(KEYINPUT24), .B(G110), .Z(new_n561));
  AOI22_X1  g375(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n555), .A2(new_n562), .ZN(new_n563));
  OAI22_X1  g377(.A1(new_n559), .A2(G110), .B1(new_n560), .B2(new_n561), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n353), .A2(new_n357), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n224), .A2(G221), .A3(G234), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n568), .B(KEYINPUT22), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(G137), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n570), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n566), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  OAI22_X1  g388(.A1(new_n574), .A2(G902), .B1(KEYINPUT72), .B2(KEYINPUT25), .ZN(new_n575));
  INV_X1    g389(.A(G217), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(G234), .B2(new_n299), .ZN(new_n577));
  NOR2_X1   g391(.A1(KEYINPUT72), .A2(KEYINPUT25), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n571), .A2(new_n299), .A3(new_n573), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n575), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n577), .A2(G902), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n571), .A2(new_n573), .A3(new_n581), .ZN(new_n582));
  AND2_X1   g396(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n481), .A2(new_n485), .A3(new_n554), .A4(new_n583), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(G101), .ZN(G3));
  OR2_X1    g399(.A1(new_n484), .A2(KEYINPUT93), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n389), .B1(new_n401), .B2(G107), .ZN(new_n587));
  AOI211_X1 g401(.A(new_n409), .B(new_n385), .C1(new_n587), .C2(new_n413), .ZN(new_n588));
  AOI21_X1  g402(.A(new_n416), .B1(new_n414), .B2(new_n415), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT33), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n410), .A2(new_n591), .A3(new_n417), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(G478), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n418), .A2(new_n419), .ZN(new_n594));
  NAND2_X1  g408(.A1(G478), .A2(G902), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(KEYINPUT94), .ZN(new_n597));
  INV_X1    g411(.A(KEYINPUT94), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n593), .A2(new_n598), .A3(new_n594), .A4(new_n595), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n597), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n382), .ZN(new_n601));
  INV_X1    g415(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n484), .A2(KEYINPUT93), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n586), .A2(new_n602), .A3(new_n319), .A4(new_n603), .ZN(new_n604));
  AND2_X1   g418(.A1(new_n477), .A2(new_n479), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n539), .B2(G902), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n532), .A2(new_n533), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n605), .A2(new_n606), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n583), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(KEYINPUT34), .B(G104), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  NOR2_X1   g426(.A1(new_n484), .A2(KEYINPUT93), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT93), .ZN(new_n614));
  AOI211_X1 g428(.A(new_n614), .B(new_n483), .C1(new_n301), .C2(new_n308), .ZN(new_n615));
  INV_X1    g429(.A(new_n382), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n421), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n613), .A2(new_n615), .A3(new_n318), .A4(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n583), .A3(new_n608), .ZN(new_n619));
  XOR2_X1   g433(.A(KEYINPUT35), .B(G107), .Z(new_n620));
  XNOR2_X1  g434(.A(new_n619), .B(new_n620), .ZN(G9));
  AND2_X1   g435(.A1(new_n606), .A2(new_n607), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n566), .A2(KEYINPUT95), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n566), .A2(KEYINPUT95), .ZN(new_n624));
  OR4_X1    g438(.A1(KEYINPUT36), .A2(new_n623), .A3(new_n624), .A4(new_n572), .ZN(new_n625));
  OAI22_X1  g439(.A1(new_n623), .A2(new_n624), .B1(KEYINPUT36), .B2(new_n572), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n581), .A3(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n580), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n481), .A2(new_n485), .A3(new_n622), .A4(new_n628), .ZN(new_n629));
  XOR2_X1   g443(.A(new_n629), .B(KEYINPUT37), .Z(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(G110), .ZN(G12));
  NOR2_X1   g445(.A1(new_n613), .A2(new_n615), .ZN(new_n632));
  OR2_X1    g446(.A1(new_n316), .A2(G900), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n617), .B1(new_n312), .B2(new_n633), .ZN(new_n634));
  AND2_X1   g448(.A1(new_n605), .A2(new_n628), .ZN(new_n635));
  NAND4_X1  g449(.A1(new_n632), .A2(new_n554), .A3(new_n634), .A4(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G128), .ZN(G30));
  NOR2_X1   g451(.A1(new_n512), .A2(new_n522), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n506), .B1(new_n542), .B2(new_n494), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n299), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n534), .A2(new_n541), .A3(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n534), .A2(new_n541), .A3(new_n641), .A4(KEYINPUT96), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n633), .A2(new_n312), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT39), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n605), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(KEYINPUT40), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n647), .A2(new_n628), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n382), .A2(new_n421), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n483), .B(new_n653), .C1(new_n650), .C2(KEYINPUT40), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n309), .B(KEYINPUT38), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n652), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n657));
  OR2_X1    g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n656), .A2(new_n657), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n192), .ZN(G45));
  NAND4_X1  g475(.A1(new_n597), .A2(new_n382), .A3(new_n599), .A4(new_n648), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n632), .A2(new_n664), .A3(new_n554), .A4(new_n635), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  INV_X1    g480(.A(new_n464), .ZN(new_n667));
  INV_X1    g481(.A(new_n467), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n423), .B1(new_n669), .B2(new_n299), .ZN(new_n670));
  INV_X1    g484(.A(new_n468), .ZN(new_n671));
  INV_X1    g485(.A(new_n479), .ZN(new_n672));
  NOR3_X1   g486(.A1(new_n670), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n554), .A2(new_n583), .A3(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT99), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n613), .A2(new_n615), .A3(new_n318), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n674), .A2(new_n675), .A3(new_n602), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n554), .A2(new_n583), .A3(new_n673), .ZN(new_n678));
  OAI21_X1  g492(.A(KEYINPUT99), .B1(new_n604), .B2(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(KEYINPUT41), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(G113), .ZN(G15));
  NAND2_X1  g496(.A1(new_n618), .A2(new_n674), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  AND4_X1   g498(.A1(new_n586), .A2(new_n603), .A3(new_n628), .A4(new_n673), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n554), .A2(new_n319), .A3(new_n422), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  AND2_X1   g502(.A1(new_n632), .A2(new_n673), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n544), .A2(KEYINPUT100), .A3(new_n500), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT100), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n691), .B1(new_n543), .B2(new_n501), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n690), .A2(new_n550), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n693), .B1(new_n531), .B2(new_n524), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n533), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n695), .A2(new_n583), .A3(new_n606), .ZN(new_n696));
  INV_X1    g510(.A(new_n653), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n689), .A2(new_n696), .A3(new_n319), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G122), .ZN(G24));
  AND3_X1   g513(.A1(new_n695), .A2(new_n606), .A3(new_n628), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n632), .A2(new_n664), .A3(new_n673), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  AND2_X1   g516(.A1(new_n554), .A2(new_n583), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n301), .A2(new_n308), .A3(new_n320), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(KEYINPUT102), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n476), .B(KEYINPUT101), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n468), .A2(new_n475), .A3(new_n706), .ZN(new_n707));
  AND2_X1   g521(.A1(new_n707), .A2(new_n479), .ZN(new_n708));
  INV_X1    g522(.A(KEYINPUT102), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n301), .A2(new_n308), .A3(new_n709), .A4(new_n320), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n705), .A2(new_n708), .A3(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n703), .A2(new_n664), .A3(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT42), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT32), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n539), .B2(new_n540), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n534), .A2(new_n716), .A3(new_n553), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n583), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n662), .B(KEYINPUT98), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n705), .A2(new_n708), .A3(new_n710), .ZN(new_n720));
  NOR4_X1   g534(.A1(new_n718), .A2(new_n719), .A3(new_n720), .A4(KEYINPUT103), .ZN(new_n721));
  INV_X1    g535(.A(KEYINPUT103), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n717), .A2(KEYINPUT42), .A3(new_n583), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n714), .B1(new_n721), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G131), .ZN(G33));
  NAND3_X1  g541(.A1(new_n703), .A2(new_n634), .A3(new_n711), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G134), .ZN(G36));
  OAI21_X1  g543(.A(new_n472), .B1(new_n474), .B2(new_n450), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(KEYINPUT45), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G469), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n706), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT46), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(KEYINPUT46), .A3(new_n706), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n735), .A2(new_n468), .A3(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n737), .A2(new_n479), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n649), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n705), .A2(new_n710), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n600), .A2(new_n616), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT43), .Z(new_n743));
  INV_X1    g557(.A(new_n622), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n628), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT44), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n741), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n739), .B(new_n747), .C1(new_n746), .C2(new_n745), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n434), .ZN(G39));
  INV_X1    g563(.A(KEYINPUT47), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n737), .A2(new_n479), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n751), .A2(KEYINPUT104), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n750), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(new_n754), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT47), .A3(new_n752), .ZN(new_n757));
  NOR4_X1   g571(.A1(new_n719), .A2(new_n740), .A3(new_n554), .A4(new_n583), .ZN(new_n758));
  AOI22_X1  g572(.A1(new_n755), .A2(new_n757), .B1(KEYINPUT105), .B2(new_n758), .ZN(new_n759));
  OR2_X1    g573(.A1(new_n758), .A2(KEYINPUT105), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G140), .ZN(G42));
  INV_X1    g576(.A(KEYINPUT115), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n743), .A2(new_n763), .A3(new_n313), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n763), .B1(new_n743), .B2(new_n313), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n670), .A2(new_n671), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n740), .A2(new_n672), .A3(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n717), .A2(new_n583), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT48), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n766), .A2(new_n689), .A3(new_n696), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n310), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n647), .A2(new_n583), .A3(new_n313), .A4(new_n769), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(new_n601), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n776), .A2(KEYINPUT118), .A3(new_n778), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n774), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n755), .B(new_n757), .C1(new_n479), .C2(new_n768), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n784), .A2(new_n696), .A3(new_n741), .A4(new_n766), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT50), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n673), .A2(new_n483), .ZN(new_n787));
  OAI221_X1 g601(.A(new_n696), .B1(KEYINPUT116), .B2(new_n787), .C1(new_n764), .C2(new_n765), .ZN(new_n788));
  INV_X1    g602(.A(new_n655), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(KEYINPUT116), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n786), .A2(new_n792), .B1(new_n770), .B2(new_n700), .ZN(new_n793));
  OAI21_X1  g607(.A(KEYINPUT50), .B1(new_n788), .B2(new_n791), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n785), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g609(.A(KEYINPUT51), .B1(new_n785), .B2(KEYINPUT117), .ZN(new_n796));
  OR3_X1    g610(.A1(new_n777), .A2(new_n382), .A3(new_n600), .ZN(new_n797));
  NAND3_X1  g611(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n785), .A2(new_n793), .A3(new_n797), .A4(new_n794), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n785), .A2(KEYINPUT117), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n799), .B1(new_n800), .B2(KEYINPUT51), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n783), .B1(new_n798), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n803));
  AOI22_X1  g617(.A1(new_n685), .A2(new_n686), .B1(new_n618), .B2(new_n674), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n680), .A2(new_n804), .A3(new_n698), .ZN(new_n805));
  XOR2_X1   g619(.A(new_n805), .B(KEYINPUT114), .Z(new_n806));
  INV_X1    g620(.A(new_n321), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n601), .A2(new_n617), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n608), .A2(new_n807), .A3(new_n808), .A4(new_n583), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n584), .A2(new_n629), .A3(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n613), .A2(new_n615), .A3(new_n653), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n627), .A2(new_n580), .A3(new_n648), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT109), .ZN(new_n814));
  NAND4_X1  g628(.A1(new_n646), .A2(new_n708), .A3(new_n812), .A4(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n665), .A2(new_n701), .A3(new_n636), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT110), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n701), .A2(new_n636), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT110), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n819), .A2(new_n820), .A3(new_n665), .A4(new_n815), .ZN(new_n821));
  XNOR2_X1  g635(.A(KEYINPUT111), .B(KEYINPUT52), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n818), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n817), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(KEYINPUT52), .A3(new_n815), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n811), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n664), .A2(new_n700), .A3(new_n708), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n635), .A2(new_n554), .A3(new_n422), .A4(new_n648), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n740), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n726), .A2(new_n728), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n806), .A2(new_n810), .A3(new_n826), .A4(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n680), .A2(new_n810), .A3(new_n804), .A4(new_n698), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n834), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n680), .A2(new_n810), .A3(new_n804), .A4(new_n698), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n711), .A2(new_n664), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT103), .B1(new_n838), .B2(new_n718), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n723), .A2(new_n724), .A3(new_n722), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n829), .B1(new_n841), .B2(new_n714), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n837), .A2(new_n842), .A3(KEYINPUT108), .A4(new_n728), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n818), .B2(new_n821), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n818), .A2(new_n821), .A3(new_n844), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n836), .B(new_n843), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n847), .A2(new_n848), .A3(new_n811), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n848), .B1(new_n847), .B2(new_n811), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n803), .B(new_n833), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n836), .A2(new_n843), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n846), .A2(new_n845), .ZN(new_n853));
  OAI21_X1  g667(.A(KEYINPUT53), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT53), .B1(new_n823), .B2(new_n825), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n855), .A2(new_n836), .A3(new_n843), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n854), .A2(KEYINPUT54), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT112), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n854), .A2(KEYINPUT112), .A3(KEYINPUT54), .A4(new_n856), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n802), .A2(new_n851), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n772), .A2(new_n773), .ZN(new_n863));
  OAI22_X1  g677(.A1(new_n862), .A2(new_n863), .B1(G952), .B2(G953), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT49), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n583), .B1(new_n767), .B2(new_n865), .ZN(new_n866));
  NOR4_X1   g680(.A1(new_n866), .A2(new_n742), .A3(new_n483), .A4(new_n672), .ZN(new_n867));
  XOR2_X1   g681(.A(new_n867), .B(KEYINPUT106), .Z(new_n868));
  NAND2_X1  g682(.A1(new_n767), .A2(new_n865), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n868), .A2(new_n789), .A3(new_n647), .A4(new_n869), .ZN(new_n870));
  XNOR2_X1  g684(.A(new_n870), .B(KEYINPUT107), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n864), .A2(new_n871), .ZN(G75));
  NOR2_X1   g686(.A1(new_n224), .A2(G952), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n833), .B1(new_n849), .B2(new_n850), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n874), .A2(G210), .A3(G902), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n304), .A2(new_n305), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n877), .A2(new_n282), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT55), .ZN(new_n879));
  OR2_X1    g693(.A1(new_n879), .A2(KEYINPUT120), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT56), .B1(new_n880), .B2(KEYINPUT119), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n876), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g696(.A1(KEYINPUT119), .A2(KEYINPUT56), .ZN(new_n883));
  OR2_X1    g697(.A1(new_n883), .A2(KEYINPUT120), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n879), .B1(new_n875), .B2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n873), .B1(new_n882), .B2(new_n885), .ZN(G51));
  NAND2_X1  g700(.A1(new_n874), .A2(KEYINPUT54), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n887), .A2(new_n851), .ZN(new_n888));
  XOR2_X1   g702(.A(new_n706), .B(KEYINPUT57), .Z(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n669), .B(KEYINPUT121), .Z(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n732), .B(KEYINPUT122), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n874), .A2(G902), .A3(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n873), .B1(new_n892), .B2(new_n894), .ZN(G54));
  INV_X1    g709(.A(KEYINPUT123), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n897));
  OAI21_X1  g711(.A(new_n896), .B1(new_n897), .B2(new_n322), .ZN(new_n898));
  NAND3_X1  g712(.A1(KEYINPUT123), .A2(KEYINPUT58), .A3(G475), .ZN(new_n899));
  NAND4_X1  g713(.A1(new_n874), .A2(G902), .A3(new_n898), .A4(new_n899), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n367), .A2(new_n374), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n900), .A2(new_n902), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n903), .A2(new_n904), .A3(new_n873), .ZN(G60));
  INV_X1    g719(.A(new_n873), .ZN(new_n906));
  XOR2_X1   g720(.A(new_n595), .B(KEYINPUT59), .Z(new_n907));
  AOI21_X1  g721(.A(new_n907), .B1(new_n861), .B2(new_n851), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n590), .A2(new_n592), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n906), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT124), .ZN(new_n911));
  INV_X1    g725(.A(new_n909), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n912), .A2(new_n907), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n888), .B2(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n913), .ZN(new_n915));
  AOI211_X1 g729(.A(KEYINPUT124), .B(new_n915), .C1(new_n887), .C2(new_n851), .ZN(new_n916));
  NOR3_X1   g730(.A1(new_n910), .A2(new_n914), .A3(new_n916), .ZN(G63));
  NAND2_X1  g731(.A1(G217), .A2(G902), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  NAND2_X1  g733(.A1(new_n874), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n574), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n874), .A2(new_n625), .A3(new_n626), .A4(new_n919), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n921), .A2(new_n906), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n921), .A2(KEYINPUT61), .A3(new_n906), .A4(new_n922), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n925), .A2(new_n926), .ZN(G66));
  INV_X1    g741(.A(G224), .ZN(new_n928));
  OAI21_X1  g742(.A(G953), .B1(new_n315), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n835), .B(KEYINPUT125), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n929), .B1(new_n930), .B2(G953), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n279), .B(new_n281), .C1(G898), .C2(new_n224), .ZN(new_n932));
  XNOR2_X1  g746(.A(new_n932), .B(KEYINPUT126), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n931), .B(new_n933), .ZN(G69));
  XOR2_X1   g748(.A(new_n525), .B(new_n372), .Z(new_n935));
  NAND2_X1  g749(.A1(G900), .A2(G953), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n748), .B1(new_n759), .B2(new_n760), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n738), .A2(new_n649), .A3(new_n771), .A4(new_n812), .ZN(new_n938));
  AND3_X1   g752(.A1(new_n938), .A2(new_n726), .A3(new_n824), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n937), .A2(new_n728), .A3(new_n939), .ZN(new_n940));
  OAI211_X1 g754(.A(new_n935), .B(new_n936), .C1(new_n940), .C2(G953), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n658), .A2(new_n659), .A3(new_n824), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT62), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n740), .A2(new_n650), .ZN(new_n945));
  NAND3_X1  g759(.A1(new_n703), .A2(new_n945), .A3(new_n808), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n944), .A2(new_n937), .A3(new_n946), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(new_n224), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n941), .B1(new_n948), .B2(new_n935), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n224), .B1(G227), .B2(G900), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n949), .B(new_n950), .ZN(G72));
  NAND2_X1  g765(.A1(G472), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT63), .Z(new_n953));
  INV_X1    g767(.A(new_n930), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n953), .B1(new_n940), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n494), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n522), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n550), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n944), .A2(new_n930), .A3(new_n937), .A4(new_n946), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n959), .A2(KEYINPUT127), .A3(new_n953), .ZN(new_n960));
  INV_X1    g774(.A(new_n957), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n506), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g776(.A(KEYINPUT127), .B1(new_n959), .B2(new_n953), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n906), .B(new_n958), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n546), .A2(new_n638), .ZN(new_n965));
  AND4_X1   g779(.A1(new_n854), .A2(new_n856), .A3(new_n953), .A4(new_n965), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n964), .A2(new_n966), .ZN(G57));
endmodule


