

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(n700), .A2(n920), .ZN(n695) );
  NAND2_X1 U557 ( .A1(n751), .A2(n750), .ZN(n764) );
  AND2_X1 U558 ( .A1(G138), .A2(n873), .ZN(n523) );
  AND2_X1 U559 ( .A1(n529), .A2(n528), .ZN(n524) );
  OR2_X1 U560 ( .A1(n774), .A2(n773), .ZN(n525) );
  AND2_X1 U561 ( .A1(n804), .A2(n1003), .ZN(n526) );
  NOR2_X1 U562 ( .A1(n734), .A2(n971), .ZN(n690) );
  NOR2_X1 U563 ( .A1(n921), .A2(n691), .ZN(n693) );
  INV_X1 U564 ( .A(KEYINPUT97), .ZN(n703) );
  XNOR2_X1 U565 ( .A(n704), .B(n703), .ZN(n711) );
  XNOR2_X1 U566 ( .A(n742), .B(KEYINPUT32), .ZN(n751) );
  NAND2_X1 U567 ( .A1(n776), .A2(n685), .ZN(n734) );
  NOR2_X1 U568 ( .A1(G164), .A2(G1384), .ZN(n776) );
  NOR2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n527) );
  NOR2_X1 U570 ( .A1(n805), .A2(n526), .ZN(n806) );
  XOR2_X1 U571 ( .A(KEYINPUT15), .B(n593), .Z(n920) );
  XOR2_X1 U572 ( .A(KEYINPUT1), .B(n535), .Z(n653) );
  NOR2_X1 U573 ( .A1(G651), .A2(n649), .ZN(n648) );
  NAND2_X1 U574 ( .A1(n524), .A2(n531), .ZN(n532) );
  NOR2_X1 U575 ( .A1(n555), .A2(n554), .ZN(G160) );
  XOR2_X2 U576 ( .A(KEYINPUT17), .B(n527), .Z(n873) );
  AND2_X1 U577 ( .A1(G2104), .A2(G2105), .ZN(n878) );
  NAND2_X1 U578 ( .A1(G114), .A2(n878), .ZN(n529) );
  INV_X1 U579 ( .A(G2104), .ZN(n530) );
  NOR2_X2 U580 ( .A1(G2105), .A2(n530), .ZN(n874) );
  NAND2_X1 U581 ( .A1(G102), .A2(n874), .ZN(n528) );
  AND2_X1 U582 ( .A1(n530), .A2(G2105), .ZN(n881) );
  NAND2_X1 U583 ( .A1(G126), .A2(n881), .ZN(n531) );
  NOR2_X1 U584 ( .A1(n523), .A2(n532), .ZN(n533) );
  XOR2_X1 U585 ( .A(KEYINPUT87), .B(n533), .Z(G164) );
  XNOR2_X1 U586 ( .A(G543), .B(KEYINPUT0), .ZN(n534) );
  XNOR2_X1 U587 ( .A(n534), .B(KEYINPUT65), .ZN(n649) );
  NAND2_X1 U588 ( .A1(n648), .A2(G51), .ZN(n537) );
  XOR2_X1 U589 ( .A(G651), .B(KEYINPUT66), .Z(n540) );
  NOR2_X1 U590 ( .A1(G543), .A2(n540), .ZN(n535) );
  NAND2_X1 U591 ( .A1(G63), .A2(n653), .ZN(n536) );
  NAND2_X1 U592 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U593 ( .A(KEYINPUT6), .B(n538), .ZN(n545) );
  NOR2_X1 U594 ( .A1(G651), .A2(G543), .ZN(n638) );
  NAND2_X1 U595 ( .A1(n638), .A2(G89), .ZN(n539) );
  XNOR2_X1 U596 ( .A(n539), .B(KEYINPUT4), .ZN(n542) );
  NOR2_X1 U597 ( .A1(n649), .A2(n540), .ZN(n642) );
  NAND2_X1 U598 ( .A1(G76), .A2(n642), .ZN(n541) );
  NAND2_X1 U599 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U600 ( .A(n543), .B(KEYINPUT5), .Z(n544) );
  NOR2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U602 ( .A(KEYINPUT7), .B(n546), .Z(n547) );
  XNOR2_X1 U603 ( .A(KEYINPUT76), .B(n547), .ZN(G168) );
  XOR2_X1 U604 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U605 ( .A1(G125), .A2(n881), .ZN(n548) );
  XNOR2_X1 U606 ( .A(n548), .B(KEYINPUT64), .ZN(n551) );
  NAND2_X1 U607 ( .A1(G101), .A2(n874), .ZN(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT23), .B(n549), .Z(n550) );
  NAND2_X1 U609 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G113), .A2(n878), .ZN(n553) );
  NAND2_X1 U611 ( .A1(G137), .A2(n873), .ZN(n552) );
  NAND2_X1 U612 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U613 ( .A1(n648), .A2(G52), .ZN(n557) );
  NAND2_X1 U614 ( .A1(G64), .A2(n653), .ZN(n556) );
  NAND2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n564) );
  NAND2_X1 U616 ( .A1(G77), .A2(n642), .ZN(n558) );
  XNOR2_X1 U617 ( .A(n558), .B(KEYINPUT68), .ZN(n560) );
  NAND2_X1 U618 ( .A1(G90), .A2(n638), .ZN(n559) );
  NAND2_X1 U619 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT9), .B(n561), .ZN(n562) );
  XNOR2_X1 U621 ( .A(KEYINPUT69), .B(n562), .ZN(n563) );
  NOR2_X1 U622 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U623 ( .A(KEYINPUT70), .B(n565), .ZN(G171) );
  INV_X1 U624 ( .A(G171), .ZN(G301) );
  AND2_X1 U625 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U626 ( .A(G57), .ZN(G237) );
  INV_X1 U627 ( .A(G132), .ZN(G219) );
  NAND2_X1 U628 ( .A1(n638), .A2(G88), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G75), .A2(n642), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n648), .A2(G50), .ZN(n569) );
  NAND2_X1 U632 ( .A1(G62), .A2(n653), .ZN(n568) );
  NAND2_X1 U633 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U634 ( .A1(n571), .A2(n570), .ZN(G166) );
  NAND2_X1 U635 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U636 ( .A(n572), .B(KEYINPUT10), .ZN(n573) );
  XNOR2_X1 U637 ( .A(KEYINPUT72), .B(n573), .ZN(G223) );
  INV_X1 U638 ( .A(G223), .ZN(n824) );
  NAND2_X1 U639 ( .A1(n824), .A2(G567), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n574), .B(KEYINPUT11), .ZN(n575) );
  XNOR2_X1 U641 ( .A(KEYINPUT73), .B(n575), .ZN(G234) );
  NAND2_X1 U642 ( .A1(n653), .A2(G56), .ZN(n576) );
  XOR2_X1 U643 ( .A(KEYINPUT14), .B(n576), .Z(n582) );
  NAND2_X1 U644 ( .A1(n638), .A2(G81), .ZN(n577) );
  XNOR2_X1 U645 ( .A(n577), .B(KEYINPUT12), .ZN(n579) );
  NAND2_X1 U646 ( .A1(G68), .A2(n642), .ZN(n578) );
  NAND2_X1 U647 ( .A1(n579), .A2(n578), .ZN(n580) );
  XOR2_X1 U648 ( .A(KEYINPUT13), .B(n580), .Z(n581) );
  NOR2_X1 U649 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U650 ( .A1(n648), .A2(G43), .ZN(n583) );
  NAND2_X1 U651 ( .A1(n584), .A2(n583), .ZN(n921) );
  INV_X1 U652 ( .A(G860), .ZN(n606) );
  OR2_X1 U653 ( .A1(n921), .A2(n606), .ZN(G153) );
  NAND2_X1 U654 ( .A1(n648), .A2(G54), .ZN(n592) );
  NAND2_X1 U655 ( .A1(n638), .A2(G92), .ZN(n586) );
  NAND2_X1 U656 ( .A1(G79), .A2(n642), .ZN(n585) );
  NAND2_X1 U657 ( .A1(n586), .A2(n585), .ZN(n590) );
  INV_X1 U658 ( .A(KEYINPUT74), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n653), .A2(G66), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n588), .B(n587), .ZN(n589) );
  NOR2_X1 U661 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U662 ( .A1(n592), .A2(n591), .ZN(n593) );
  INV_X1 U663 ( .A(n920), .ZN(n621) );
  NOR2_X1 U664 ( .A1(n621), .A2(G868), .ZN(n594) );
  XNOR2_X1 U665 ( .A(n594), .B(KEYINPUT75), .ZN(n596) );
  NAND2_X1 U666 ( .A1(G868), .A2(G301), .ZN(n595) );
  NAND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(G284) );
  NAND2_X1 U668 ( .A1(n648), .A2(G53), .ZN(n598) );
  NAND2_X1 U669 ( .A1(G65), .A2(n653), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n598), .A2(n597), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n638), .A2(G91), .ZN(n600) );
  NAND2_X1 U672 ( .A1(G78), .A2(n642), .ZN(n599) );
  NAND2_X1 U673 ( .A1(n600), .A2(n599), .ZN(n601) );
  NOR2_X1 U674 ( .A1(n602), .A2(n601), .ZN(n926) );
  INV_X1 U675 ( .A(n926), .ZN(G299) );
  XNOR2_X1 U676 ( .A(KEYINPUT77), .B(G868), .ZN(n603) );
  NOR2_X1 U677 ( .A1(G286), .A2(n603), .ZN(n605) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n604) );
  NOR2_X1 U679 ( .A1(n605), .A2(n604), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n606), .A2(G559), .ZN(n607) );
  NAND2_X1 U681 ( .A1(n607), .A2(n621), .ZN(n608) );
  XNOR2_X1 U682 ( .A(n608), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n921), .ZN(n611) );
  NAND2_X1 U684 ( .A1(n621), .A2(G868), .ZN(n609) );
  NOR2_X1 U685 ( .A1(G559), .A2(n609), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n611), .A2(n610), .ZN(G282) );
  NAND2_X1 U687 ( .A1(n881), .A2(G123), .ZN(n612) );
  XNOR2_X1 U688 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G111), .A2(n878), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G135), .A2(n873), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G99), .A2(n874), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  NOR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n998) );
  XNOR2_X1 U695 ( .A(G2096), .B(n998), .ZN(n620) );
  INV_X1 U696 ( .A(G2100), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(G156) );
  NAND2_X1 U698 ( .A1(G559), .A2(n621), .ZN(n622) );
  XNOR2_X1 U699 ( .A(n622), .B(n921), .ZN(n664) );
  NOR2_X1 U700 ( .A1(G860), .A2(n664), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n648), .A2(G55), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G67), .A2(n653), .ZN(n623) );
  NAND2_X1 U703 ( .A1(n624), .A2(n623), .ZN(n628) );
  NAND2_X1 U704 ( .A1(n638), .A2(G93), .ZN(n626) );
  NAND2_X1 U705 ( .A1(G80), .A2(n642), .ZN(n625) );
  NAND2_X1 U706 ( .A1(n626), .A2(n625), .ZN(n627) );
  NOR2_X1 U707 ( .A1(n628), .A2(n627), .ZN(n658) );
  XNOR2_X1 U708 ( .A(n658), .B(KEYINPUT78), .ZN(n629) );
  XNOR2_X1 U709 ( .A(n630), .B(n629), .ZN(G145) );
  NAND2_X1 U710 ( .A1(n648), .A2(G47), .ZN(n632) );
  NAND2_X1 U711 ( .A1(G72), .A2(n642), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(n636) );
  NAND2_X1 U713 ( .A1(n638), .A2(G85), .ZN(n634) );
  NAND2_X1 U714 ( .A1(G60), .A2(n653), .ZN(n633) );
  NAND2_X1 U715 ( .A1(n634), .A2(n633), .ZN(n635) );
  NOR2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U717 ( .A(n637), .B(KEYINPUT67), .ZN(G290) );
  NAND2_X1 U718 ( .A1(n638), .A2(G86), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G61), .A2(n653), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U721 ( .A(KEYINPUT80), .B(n641), .ZN(n645) );
  NAND2_X1 U722 ( .A1(G73), .A2(n642), .ZN(n643) );
  XOR2_X1 U723 ( .A(KEYINPUT2), .B(n643), .Z(n644) );
  NOR2_X1 U724 ( .A1(n645), .A2(n644), .ZN(n647) );
  NAND2_X1 U725 ( .A1(n648), .A2(G48), .ZN(n646) );
  NAND2_X1 U726 ( .A1(n647), .A2(n646), .ZN(G305) );
  NAND2_X1 U727 ( .A1(n648), .A2(G49), .ZN(n655) );
  NAND2_X1 U728 ( .A1(G87), .A2(n649), .ZN(n651) );
  NAND2_X1 U729 ( .A1(G74), .A2(G651), .ZN(n650) );
  NAND2_X1 U730 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U732 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U733 ( .A(KEYINPUT79), .B(n656), .Z(G288) );
  NOR2_X1 U734 ( .A1(G868), .A2(n658), .ZN(n657) );
  XOR2_X1 U735 ( .A(n657), .B(KEYINPUT82), .Z(n668) );
  XNOR2_X1 U736 ( .A(n926), .B(KEYINPUT19), .ZN(n663) );
  XNOR2_X1 U737 ( .A(G166), .B(n658), .ZN(n661) );
  XOR2_X1 U738 ( .A(G305), .B(G288), .Z(n659) );
  XNOR2_X1 U739 ( .A(G290), .B(n659), .ZN(n660) );
  XNOR2_X1 U740 ( .A(n661), .B(n660), .ZN(n662) );
  XNOR2_X1 U741 ( .A(n663), .B(n662), .ZN(n852) );
  XNOR2_X1 U742 ( .A(n852), .B(KEYINPUT81), .ZN(n665) );
  XNOR2_X1 U743 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U744 ( .A1(G868), .A2(n666), .ZN(n667) );
  NAND2_X1 U745 ( .A1(n668), .A2(n667), .ZN(G295) );
  NAND2_X1 U746 ( .A1(G2078), .A2(G2084), .ZN(n669) );
  XNOR2_X1 U747 ( .A(n669), .B(KEYINPUT20), .ZN(n670) );
  XNOR2_X1 U748 ( .A(n670), .B(KEYINPUT83), .ZN(n671) );
  NAND2_X1 U749 ( .A1(n671), .A2(G2090), .ZN(n672) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U751 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XNOR2_X1 U753 ( .A(KEYINPUT71), .B(G82), .ZN(G220) );
  NOR2_X1 U754 ( .A1(G219), .A2(G220), .ZN(n674) );
  XOR2_X1 U755 ( .A(KEYINPUT22), .B(n674), .Z(n675) );
  XNOR2_X1 U756 ( .A(n675), .B(KEYINPUT84), .ZN(n676) );
  NOR2_X1 U757 ( .A1(G218), .A2(n676), .ZN(n677) );
  NAND2_X1 U758 ( .A1(G96), .A2(n677), .ZN(n831) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n831), .ZN(n681) );
  NAND2_X1 U760 ( .A1(G120), .A2(G69), .ZN(n678) );
  NOR2_X1 U761 ( .A1(G237), .A2(n678), .ZN(n679) );
  NAND2_X1 U762 ( .A1(G108), .A2(n679), .ZN(n832) );
  NAND2_X1 U763 ( .A1(G567), .A2(n832), .ZN(n680) );
  NAND2_X1 U764 ( .A1(n681), .A2(n680), .ZN(n682) );
  XOR2_X1 U765 ( .A(KEYINPUT85), .B(n682), .Z(n851) );
  NAND2_X1 U766 ( .A1(G661), .A2(G483), .ZN(n683) );
  NOR2_X1 U767 ( .A1(n851), .A2(n683), .ZN(n828) );
  NAND2_X1 U768 ( .A1(G36), .A2(n828), .ZN(n684) );
  XNOR2_X1 U769 ( .A(n684), .B(KEYINPUT86), .ZN(G176) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NAND2_X1 U771 ( .A1(G160), .A2(G40), .ZN(n775) );
  INV_X1 U772 ( .A(n775), .ZN(n685) );
  NAND2_X1 U773 ( .A1(G8), .A2(n734), .ZN(n765) );
  NOR2_X1 U774 ( .A1(G1981), .A2(G305), .ZN(n686) );
  XOR2_X1 U775 ( .A(n686), .B(KEYINPUT24), .Z(n687) );
  NOR2_X1 U776 ( .A1(n765), .A2(n687), .ZN(n688) );
  XNOR2_X1 U777 ( .A(n688), .B(KEYINPUT91), .ZN(n755) );
  NOR2_X1 U778 ( .A1(G2090), .A2(G303), .ZN(n689) );
  NAND2_X1 U779 ( .A1(G8), .A2(n689), .ZN(n752) );
  XNOR2_X1 U780 ( .A(G1996), .B(KEYINPUT95), .ZN(n971) );
  XNOR2_X1 U781 ( .A(n690), .B(KEYINPUT26), .ZN(n691) );
  NAND2_X1 U782 ( .A1(G1341), .A2(n734), .ZN(n692) );
  NAND2_X1 U783 ( .A1(n693), .A2(n692), .ZN(n700) );
  INV_X1 U784 ( .A(KEYINPUT96), .ZN(n694) );
  XNOR2_X1 U785 ( .A(n695), .B(n694), .ZN(n699) );
  INV_X1 U786 ( .A(n734), .ZN(n718) );
  NOR2_X1 U787 ( .A1(n718), .A2(G1348), .ZN(n697) );
  NOR2_X1 U788 ( .A1(G2067), .A2(n734), .ZN(n696) );
  NOR2_X1 U789 ( .A1(n697), .A2(n696), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n699), .A2(n698), .ZN(n702) );
  NAND2_X1 U791 ( .A1(n700), .A2(n920), .ZN(n701) );
  NAND2_X1 U792 ( .A1(n702), .A2(n701), .ZN(n704) );
  INV_X1 U793 ( .A(G2072), .ZN(n1007) );
  NOR2_X1 U794 ( .A1(n734), .A2(n1007), .ZN(n706) );
  XOR2_X1 U795 ( .A(KEYINPUT27), .B(KEYINPUT93), .Z(n705) );
  XNOR2_X1 U796 ( .A(n706), .B(n705), .ZN(n708) );
  NAND2_X1 U797 ( .A1(n734), .A2(G1956), .ZN(n707) );
  NAND2_X1 U798 ( .A1(n708), .A2(n707), .ZN(n709) );
  XOR2_X1 U799 ( .A(KEYINPUT94), .B(n709), .Z(n712) );
  NAND2_X1 U800 ( .A1(n926), .A2(n712), .ZN(n710) );
  NAND2_X1 U801 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U802 ( .A1(n926), .A2(n712), .ZN(n713) );
  XOR2_X1 U803 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U804 ( .A1(n715), .A2(n714), .ZN(n717) );
  XOR2_X1 U805 ( .A(KEYINPUT98), .B(KEYINPUT29), .Z(n716) );
  XNOR2_X1 U806 ( .A(n717), .B(n716), .ZN(n722) );
  XOR2_X1 U807 ( .A(G2078), .B(KEYINPUT25), .Z(n972) );
  NOR2_X1 U808 ( .A1(n972), .A2(n734), .ZN(n720) );
  NOR2_X1 U809 ( .A1(n718), .A2(G1961), .ZN(n719) );
  NOR2_X1 U810 ( .A1(n720), .A2(n719), .ZN(n728) );
  OR2_X1 U811 ( .A1(G301), .A2(n728), .ZN(n721) );
  NAND2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n733) );
  NOR2_X1 U813 ( .A1(G1966), .A2(n765), .ZN(n747) );
  NOR2_X1 U814 ( .A1(G2084), .A2(n734), .ZN(n723) );
  XOR2_X1 U815 ( .A(KEYINPUT92), .B(n723), .Z(n743) );
  NAND2_X1 U816 ( .A1(G8), .A2(n743), .ZN(n724) );
  NOR2_X1 U817 ( .A1(n747), .A2(n724), .ZN(n725) );
  XOR2_X1 U818 ( .A(KEYINPUT30), .B(n725), .Z(n726) );
  NOR2_X1 U819 ( .A1(G168), .A2(n726), .ZN(n727) );
  XNOR2_X1 U820 ( .A(n727), .B(KEYINPUT99), .ZN(n730) );
  NAND2_X1 U821 ( .A1(n728), .A2(G301), .ZN(n729) );
  NAND2_X1 U822 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U823 ( .A(n731), .B(KEYINPUT31), .ZN(n732) );
  NAND2_X1 U824 ( .A1(n733), .A2(n732), .ZN(n745) );
  NAND2_X1 U825 ( .A1(n745), .A2(G286), .ZN(n740) );
  NOR2_X1 U826 ( .A1(G2090), .A2(n734), .ZN(n735) );
  XNOR2_X1 U827 ( .A(n735), .B(KEYINPUT100), .ZN(n737) );
  NOR2_X1 U828 ( .A1(n765), .A2(G1971), .ZN(n736) );
  NOR2_X1 U829 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U830 ( .A1(n738), .A2(G303), .ZN(n739) );
  NAND2_X1 U831 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U832 ( .A1(n741), .A2(G8), .ZN(n742) );
  INV_X1 U833 ( .A(n743), .ZN(n744) );
  NAND2_X1 U834 ( .A1(n744), .A2(G8), .ZN(n749) );
  INV_X1 U835 ( .A(n745), .ZN(n746) );
  NOR2_X1 U836 ( .A1(n747), .A2(n746), .ZN(n748) );
  NAND2_X1 U837 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n752), .A2(n764), .ZN(n753) );
  NAND2_X1 U839 ( .A1(n753), .A2(n765), .ZN(n754) );
  NAND2_X1 U840 ( .A1(n755), .A2(n754), .ZN(n774) );
  NAND2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n927) );
  NOR2_X1 U842 ( .A1(KEYINPUT101), .A2(n765), .ZN(n758) );
  NAND2_X1 U843 ( .A1(n927), .A2(n758), .ZN(n756) );
  INV_X1 U844 ( .A(KEYINPUT33), .ZN(n757) );
  NAND2_X1 U845 ( .A1(n756), .A2(n757), .ZN(n761) );
  OR2_X1 U846 ( .A1(G1976), .A2(G288), .ZN(n932) );
  NOR2_X1 U847 ( .A1(n932), .A2(n757), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n759), .A2(n758), .ZN(n760) );
  NAND2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n772) );
  NOR2_X1 U850 ( .A1(G1971), .A2(G303), .ZN(n762) );
  NOR2_X1 U851 ( .A1(n762), .A2(KEYINPUT33), .ZN(n763) );
  NAND2_X1 U852 ( .A1(n764), .A2(n763), .ZN(n768) );
  INV_X1 U853 ( .A(n765), .ZN(n766) );
  NAND2_X1 U854 ( .A1(n766), .A2(KEYINPUT101), .ZN(n767) );
  NAND2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n769) );
  NAND2_X1 U856 ( .A1(n769), .A2(n932), .ZN(n770) );
  XOR2_X1 U857 ( .A(G1981), .B(G305), .Z(n917) );
  NAND2_X1 U858 ( .A1(n770), .A2(n917), .ZN(n771) );
  NOR2_X1 U859 ( .A1(n772), .A2(n771), .ZN(n773) );
  NOR2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n818) );
  XNOR2_X1 U861 ( .A(KEYINPUT37), .B(G2067), .ZN(n816) );
  NAND2_X1 U862 ( .A1(G128), .A2(n881), .ZN(n778) );
  NAND2_X1 U863 ( .A1(G116), .A2(n878), .ZN(n777) );
  NAND2_X1 U864 ( .A1(n778), .A2(n777), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(KEYINPUT35), .ZN(n784) );
  NAND2_X1 U866 ( .A1(G140), .A2(n873), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G104), .A2(n874), .ZN(n780) );
  NAND2_X1 U868 ( .A1(n781), .A2(n780), .ZN(n782) );
  XOR2_X1 U869 ( .A(KEYINPUT34), .B(n782), .Z(n783) );
  NAND2_X1 U870 ( .A1(n784), .A2(n783), .ZN(n785) );
  XOR2_X1 U871 ( .A(n785), .B(KEYINPUT36), .Z(n896) );
  OR2_X1 U872 ( .A1(n816), .A2(n896), .ZN(n786) );
  XOR2_X1 U873 ( .A(KEYINPUT88), .B(n786), .Z(n1016) );
  NAND2_X1 U874 ( .A1(n818), .A2(n1016), .ZN(n815) );
  XNOR2_X1 U875 ( .A(G1986), .B(G290), .ZN(n934) );
  NAND2_X1 U876 ( .A1(n818), .A2(n934), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n815), .A2(n787), .ZN(n805) );
  XNOR2_X1 U878 ( .A(KEYINPUT90), .B(n818), .ZN(n804) );
  NAND2_X1 U879 ( .A1(G131), .A2(n873), .ZN(n789) );
  NAND2_X1 U880 ( .A1(G95), .A2(n874), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n789), .A2(n788), .ZN(n793) );
  NAND2_X1 U882 ( .A1(G119), .A2(n881), .ZN(n791) );
  NAND2_X1 U883 ( .A1(G107), .A2(n878), .ZN(n790) );
  NAND2_X1 U884 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U885 ( .A1(n793), .A2(n792), .ZN(n889) );
  NAND2_X1 U886 ( .A1(G1991), .A2(n889), .ZN(n803) );
  NAND2_X1 U887 ( .A1(G105), .A2(n874), .ZN(n794) );
  XNOR2_X1 U888 ( .A(n794), .B(KEYINPUT38), .ZN(n801) );
  NAND2_X1 U889 ( .A1(G129), .A2(n881), .ZN(n796) );
  NAND2_X1 U890 ( .A1(G141), .A2(n873), .ZN(n795) );
  NAND2_X1 U891 ( .A1(n796), .A2(n795), .ZN(n799) );
  NAND2_X1 U892 ( .A1(G117), .A2(n878), .ZN(n797) );
  XNOR2_X1 U893 ( .A(KEYINPUT89), .B(n797), .ZN(n798) );
  NOR2_X1 U894 ( .A1(n799), .A2(n798), .ZN(n800) );
  NAND2_X1 U895 ( .A1(n801), .A2(n800), .ZN(n887) );
  NAND2_X1 U896 ( .A1(G1996), .A2(n887), .ZN(n802) );
  NAND2_X1 U897 ( .A1(n803), .A2(n802), .ZN(n1003) );
  NAND2_X1 U898 ( .A1(n525), .A2(n806), .ZN(n822) );
  XOR2_X1 U899 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n813) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n887), .ZN(n996) );
  NOR2_X1 U901 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U902 ( .A1(G1991), .A2(n889), .ZN(n999) );
  NOR2_X1 U903 ( .A1(n807), .A2(n999), .ZN(n808) );
  NOR2_X1 U904 ( .A1(n526), .A2(n808), .ZN(n809) );
  XNOR2_X1 U905 ( .A(n809), .B(KEYINPUT102), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n996), .A2(n810), .ZN(n811) );
  XNOR2_X1 U907 ( .A(n811), .B(KEYINPUT39), .ZN(n812) );
  XNOR2_X1 U908 ( .A(n813), .B(n812), .ZN(n814) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n817) );
  NAND2_X1 U910 ( .A1(n896), .A2(n816), .ZN(n1013) );
  NAND2_X1 U911 ( .A1(n817), .A2(n1013), .ZN(n819) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  XOR2_X1 U913 ( .A(KEYINPUT105), .B(n820), .Z(n821) );
  NAND2_X1 U914 ( .A1(n822), .A2(n821), .ZN(n823) );
  XNOR2_X1 U915 ( .A(n823), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U916 ( .A1(n824), .A2(G2106), .ZN(n825) );
  XOR2_X1 U917 ( .A(KEYINPUT107), .B(n825), .Z(G217) );
  NAND2_X1 U918 ( .A1(G15), .A2(G2), .ZN(n826) );
  XOR2_X1 U919 ( .A(KEYINPUT108), .B(n826), .Z(n827) );
  NAND2_X1 U920 ( .A1(G661), .A2(n827), .ZN(G259) );
  NAND2_X1 U921 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U922 ( .A1(n829), .A2(n828), .ZN(n830) );
  XOR2_X1 U923 ( .A(KEYINPUT109), .B(n830), .Z(G188) );
  XOR2_X1 U924 ( .A(G69), .B(KEYINPUT110), .Z(G235) );
  INV_X1 U926 ( .A(G120), .ZN(G236) );
  NOR2_X1 U927 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U928 ( .A(G325), .ZN(G261) );
  XOR2_X1 U929 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U930 ( .A(G2072), .B(KEYINPUT42), .ZN(n833) );
  XNOR2_X1 U931 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U932 ( .A(n835), .B(G2678), .Z(n837) );
  XNOR2_X1 U933 ( .A(G2067), .B(G2090), .ZN(n836) );
  XNOR2_X1 U934 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U935 ( .A(KEYINPUT112), .B(G2100), .Z(n839) );
  XNOR2_X1 U936 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U937 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U938 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U939 ( .A(G1986), .B(G1956), .Z(n843) );
  XNOR2_X1 U940 ( .A(G1976), .B(G1971), .ZN(n842) );
  XNOR2_X1 U941 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U942 ( .A(n844), .B(G2474), .Z(n846) );
  XNOR2_X1 U943 ( .A(G1981), .B(G1966), .ZN(n845) );
  XNOR2_X1 U944 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U945 ( .A(KEYINPUT41), .B(G1961), .Z(n848) );
  XNOR2_X1 U946 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U947 ( .A(n848), .B(n847), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(G229) );
  XNOR2_X1 U949 ( .A(KEYINPUT111), .B(n851), .ZN(G319) );
  XNOR2_X1 U950 ( .A(n852), .B(n920), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n853), .B(n921), .ZN(n855) );
  XNOR2_X1 U952 ( .A(G286), .B(G301), .ZN(n854) );
  XNOR2_X1 U953 ( .A(n855), .B(n854), .ZN(n856) );
  NOR2_X1 U954 ( .A1(G37), .A2(n856), .ZN(G397) );
  NAND2_X1 U955 ( .A1(n881), .A2(G124), .ZN(n857) );
  XNOR2_X1 U956 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G112), .A2(n878), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n863) );
  NAND2_X1 U959 ( .A1(G136), .A2(n873), .ZN(n861) );
  NAND2_X1 U960 ( .A1(G100), .A2(n874), .ZN(n860) );
  NAND2_X1 U961 ( .A1(n861), .A2(n860), .ZN(n862) );
  NOR2_X1 U962 ( .A1(n863), .A2(n862), .ZN(G162) );
  NAND2_X1 U963 ( .A1(n881), .A2(G127), .ZN(n864) );
  XOR2_X1 U964 ( .A(KEYINPUT115), .B(n864), .Z(n866) );
  NAND2_X1 U965 ( .A1(n878), .A2(G115), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n867), .B(KEYINPUT47), .ZN(n869) );
  NAND2_X1 U968 ( .A1(G103), .A2(n874), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U970 ( .A1(n873), .A2(G139), .ZN(n870) );
  XOR2_X1 U971 ( .A(KEYINPUT114), .B(n870), .Z(n871) );
  NOR2_X1 U972 ( .A1(n872), .A2(n871), .ZN(n1006) );
  NAND2_X1 U973 ( .A1(G142), .A2(n873), .ZN(n876) );
  NAND2_X1 U974 ( .A1(G106), .A2(n874), .ZN(n875) );
  NAND2_X1 U975 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n877), .B(KEYINPUT45), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U979 ( .A1(G130), .A2(n881), .ZN(n882) );
  XNOR2_X1 U980 ( .A(KEYINPUT113), .B(n882), .ZN(n883) );
  NOR2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U982 ( .A(n1006), .B(n885), .ZN(n895) );
  XOR2_X1 U983 ( .A(G162), .B(n998), .Z(n886) );
  XNOR2_X1 U984 ( .A(n887), .B(n886), .ZN(n891) );
  XOR2_X1 U985 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n888) );
  XNOR2_X1 U986 ( .A(n889), .B(n888), .ZN(n890) );
  XOR2_X1 U987 ( .A(n891), .B(n890), .Z(n893) );
  XNOR2_X1 U988 ( .A(G164), .B(G160), .ZN(n892) );
  XNOR2_X1 U989 ( .A(n893), .B(n892), .ZN(n894) );
  XNOR2_X1 U990 ( .A(n895), .B(n894), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(n896), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(n899) );
  XNOR2_X1 U993 ( .A(KEYINPUT116), .B(n899), .ZN(G395) );
  NOR2_X1 U994 ( .A1(G227), .A2(G229), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n900), .B(KEYINPUT49), .ZN(n913) );
  XOR2_X1 U996 ( .A(KEYINPUT106), .B(G2446), .Z(n902) );
  XNOR2_X1 U997 ( .A(G2443), .B(G2454), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n902), .B(n901), .ZN(n903) );
  XOR2_X1 U999 ( .A(n903), .B(G2451), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G1341), .B(G1348), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1002 ( .A(G2435), .B(G2427), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2430), .B(G2438), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n910) );
  NAND2_X1 U1006 ( .A1(G14), .A2(n910), .ZN(n916) );
  NAND2_X1 U1007 ( .A1(n916), .A2(G319), .ZN(n911) );
  XOR2_X1 U1008 ( .A(KEYINPUT117), .B(n911), .Z(n912) );
  NOR2_X1 U1009 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G397), .A2(G395), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1012 ( .A(G225), .ZN(G308) );
  INV_X1 U1013 ( .A(G96), .ZN(G221) );
  INV_X1 U1014 ( .A(G108), .ZN(G238) );
  INV_X1 U1015 ( .A(n916), .ZN(G401) );
  XNOR2_X1 U1016 ( .A(G16), .B(KEYINPUT56), .ZN(n942) );
  XNOR2_X1 U1017 ( .A(G1961), .B(G171), .ZN(n940) );
  XNOR2_X1 U1018 ( .A(G1966), .B(G168), .ZN(n918) );
  NAND2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(KEYINPUT57), .B(n919), .ZN(n925) );
  XNOR2_X1 U1021 ( .A(G1348), .B(n920), .ZN(n923) );
  XNOR2_X1 U1022 ( .A(G1341), .B(n921), .ZN(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1024 ( .A1(n925), .A2(n924), .ZN(n938) );
  XNOR2_X1 U1025 ( .A(n926), .B(G1956), .ZN(n928) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1027 ( .A(G166), .B(G1971), .Z(n929) );
  XNOR2_X1 U1028 ( .A(KEYINPUT122), .B(n929), .ZN(n930) );
  NOR2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n935) );
  NOR2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(KEYINPUT123), .B(n936), .ZN(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n968) );
  INV_X1 U1036 ( .A(G16), .ZN(n966) );
  XNOR2_X1 U1037 ( .A(G1961), .B(KEYINPUT124), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(n943), .B(G5), .ZN(n950) );
  XNOR2_X1 U1039 ( .A(G1976), .B(G23), .ZN(n945) );
  XNOR2_X1 U1040 ( .A(G1971), .B(G22), .ZN(n944) );
  NOR2_X1 U1041 ( .A1(n945), .A2(n944), .ZN(n947) );
  XOR2_X1 U1042 ( .A(G1986), .B(G24), .Z(n946) );
  NAND2_X1 U1043 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1044 ( .A(KEYINPUT58), .B(n948), .ZN(n949) );
  NOR2_X1 U1045 ( .A1(n950), .A2(n949), .ZN(n961) );
  XNOR2_X1 U1046 ( .A(G1981), .B(G6), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(KEYINPUT59), .B(KEYINPUT125), .ZN(n951) );
  XNOR2_X1 U1048 ( .A(n951), .B(G4), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n952), .B(G1348), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n958) );
  XNOR2_X1 U1051 ( .A(G1956), .B(G20), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G19), .B(G1341), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1054 ( .A1(n958), .A2(n957), .ZN(n959) );
  XOR2_X1 U1055 ( .A(KEYINPUT60), .B(n959), .Z(n960) );
  NAND2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(G21), .B(G1966), .ZN(n962) );
  NOR2_X1 U1058 ( .A1(n963), .A2(n962), .ZN(n964) );
  XNOR2_X1 U1059 ( .A(KEYINPUT61), .B(n964), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  XNOR2_X1 U1062 ( .A(KEYINPUT126), .B(n969), .ZN(n993) );
  XOR2_X1 U1063 ( .A(KEYINPUT55), .B(KEYINPUT121), .Z(n990) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G35), .ZN(n984) );
  XOR2_X1 U1065 ( .A(G1991), .B(G25), .Z(n970) );
  NAND2_X1 U1066 ( .A1(n970), .A2(G28), .ZN(n981) );
  XNOR2_X1 U1067 ( .A(G32), .B(n971), .ZN(n979) );
  XNOR2_X1 U1068 ( .A(n972), .B(G27), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(G2067), .B(G26), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G33), .B(G2072), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1072 ( .A(KEYINPUT119), .B(n975), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  XNOR2_X1 U1076 ( .A(KEYINPUT53), .B(n982), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n988) );
  XOR2_X1 U1078 ( .A(KEYINPUT120), .B(G34), .Z(n986) );
  XNOR2_X1 U1079 ( .A(G2084), .B(KEYINPUT54), .ZN(n985) );
  XNOR2_X1 U1080 ( .A(n986), .B(n985), .ZN(n987) );
  NAND2_X1 U1081 ( .A1(n988), .A2(n987), .ZN(n989) );
  XNOR2_X1 U1082 ( .A(n990), .B(n989), .ZN(n991) );
  NOR2_X1 U1083 ( .A1(G29), .A2(n991), .ZN(n992) );
  NOR2_X1 U1084 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1085 ( .A1(G11), .A2(n994), .ZN(n1023) );
  XOR2_X1 U1086 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  XOR2_X1 U1088 ( .A(KEYINPUT51), .B(n997), .Z(n1005) );
  XNOR2_X1 U1089 ( .A(G160), .B(G2084), .ZN(n1001) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  NAND2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1012) );
  XOR2_X1 U1094 ( .A(G164), .B(G2078), .Z(n1009) );
  XNOR2_X1 U1095 ( .A(n1007), .B(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XOR2_X1 U1097 ( .A(KEYINPUT50), .B(n1010), .Z(n1011) );
  NOR2_X1 U1098 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  NAND2_X1 U1099 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1100 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1101 ( .A(KEYINPUT52), .B(n1017), .ZN(n1019) );
  INV_X1 U1102 ( .A(KEYINPUT55), .ZN(n1018) );
  NAND2_X1 U1103 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NAND2_X1 U1104 ( .A1(n1020), .A2(G29), .ZN(n1021) );
  XOR2_X1 U1105 ( .A(n1021), .B(KEYINPUT118), .Z(n1022) );
  NOR2_X1 U1106 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XOR2_X1 U1107 ( .A(KEYINPUT127), .B(n1024), .Z(n1025) );
  XNOR2_X1 U1108 ( .A(KEYINPUT62), .B(n1025), .ZN(G311) );
  INV_X1 U1109 ( .A(G311), .ZN(G150) );
endmodule

