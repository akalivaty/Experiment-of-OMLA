//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 0 1 1 1 0 0 0 1 1 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n696,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  OAI211_X1 g001(.A(new_n187), .B(G119), .C1(KEYINPUT71), .C2(KEYINPUT23), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT23), .ZN(new_n189));
  INV_X1    g003(.A(G119), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(G128), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  OAI21_X1  g006(.A(new_n192), .B1(new_n190), .B2(G128), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n188), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G110), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n190), .A2(G128), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n187), .A2(G119), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT70), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n187), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n190), .A2(G128), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT70), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n199), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  XOR2_X1   g016(.A(KEYINPUT24), .B(G110), .Z(new_n203));
  NAND3_X1  g017(.A1(new_n198), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  AND2_X1   g018(.A1(G125), .A2(G140), .ZN(new_n205));
  NOR2_X1   g019(.A1(G125), .A2(G140), .ZN(new_n206));
  OAI21_X1  g020(.A(KEYINPUT16), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT16), .ZN(new_n208));
  INV_X1    g022(.A(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(new_n209), .A3(G125), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(G146), .A3(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(G146), .B1(new_n207), .B2(new_n210), .ZN(new_n213));
  OAI211_X1 g027(.A(new_n195), .B(new_n204), .C1(new_n212), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G125), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n215), .A2(new_n209), .ZN(new_n216));
  NAND2_X1  g030(.A1(G125), .A2(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(G146), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n203), .B1(new_n198), .B2(new_n202), .ZN(new_n221));
  INV_X1    g035(.A(G110), .ZN(new_n222));
  OAI211_X1 g036(.A(new_n222), .B(new_n188), .C1(new_n191), .C2(new_n193), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n220), .B1(new_n221), .B2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT72), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n211), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g041(.A1(new_n207), .A2(KEYINPUT72), .A3(G146), .A4(new_n210), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n214), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g044(.A(KEYINPUT22), .B(G137), .ZN(new_n231));
  INV_X1    g045(.A(G953), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(G221), .A3(G234), .ZN(new_n233));
  XNOR2_X1  g047(.A(new_n231), .B(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n214), .B(new_n234), .C1(new_n225), .C2(new_n229), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n236), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT73), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT25), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G217), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n243), .B1(G234), .B2(new_n237), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n239), .A2(new_n241), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n236), .A2(KEYINPUT25), .A3(new_n237), .A4(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT73), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n242), .B(new_n244), .C1(new_n245), .C2(new_n247), .ZN(new_n248));
  OR2_X1    g062(.A1(new_n239), .A2(new_n244), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(G134), .ZN(new_n252));
  NAND2_X1  g066(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OR2_X1    g068(.A1(KEYINPUT65), .A2(KEYINPUT11), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n251), .A2(KEYINPUT65), .A3(KEYINPUT11), .A4(G134), .ZN(new_n256));
  INV_X1    g070(.A(G134), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G137), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n255), .A3(new_n256), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G131), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n251), .A2(G134), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n261), .B1(new_n252), .B2(new_n253), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n262), .A2(new_n263), .A3(new_n255), .A4(new_n256), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT0), .A2(G128), .ZN(new_n268));
  INV_X1    g082(.A(G143), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(KEYINPUT64), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT64), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G143), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n270), .A2(new_n272), .A3(new_n219), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n269), .A2(G146), .ZN(new_n274));
  AOI211_X1 g088(.A(new_n267), .B(new_n268), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n269), .A2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n270), .A2(new_n272), .ZN(new_n277));
  AOI211_X1 g091(.A(new_n276), .B(new_n266), .C1(new_n277), .C2(G146), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n275), .A2(new_n278), .A3(KEYINPUT67), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT67), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n273), .A2(new_n274), .ZN(new_n281));
  INV_X1    g095(.A(new_n268), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n281), .A2(new_n266), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n276), .B1(new_n277), .B2(G146), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n267), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n280), .B1(new_n283), .B2(new_n285), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n265), .B1(new_n279), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n252), .B1(new_n261), .B2(KEYINPUT66), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT66), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n258), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(G131), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT1), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(G128), .ZN(new_n293));
  AOI211_X1 g107(.A(new_n276), .B(new_n293), .C1(new_n277), .C2(G146), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n219), .A2(G143), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT1), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n273), .A2(new_n274), .B1(new_n296), .B2(G128), .ZN(new_n297));
  OAI211_X1 g111(.A(new_n264), .B(new_n291), .C1(new_n294), .C2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n287), .A2(KEYINPUT30), .A3(new_n298), .ZN(new_n299));
  XOR2_X1   g113(.A(G116), .B(G119), .Z(new_n300));
  XNOR2_X1  g114(.A(KEYINPUT2), .B(G113), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n300), .B(new_n301), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n275), .A2(new_n278), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n265), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n298), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT30), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n299), .A2(new_n302), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G237), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n232), .A3(G210), .ZN(new_n310));
  INV_X1    g124(.A(G101), .ZN(new_n311));
  XNOR2_X1  g125(.A(new_n310), .B(new_n311), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n313));
  XOR2_X1   g127(.A(new_n312), .B(new_n313), .Z(new_n314));
  INV_X1    g128(.A(new_n302), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n287), .A2(new_n315), .A3(new_n298), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n308), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT31), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT28), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n305), .A2(new_n302), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n287), .A2(KEYINPUT28), .A3(new_n315), .A4(new_n298), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(new_n314), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT31), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n308), .A2(new_n326), .A3(new_n314), .A4(new_n316), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n318), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NOR2_X1   g142(.A1(G472), .A2(G902), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(KEYINPUT32), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT32), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n332), .A3(new_n329), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n320), .A2(new_n314), .A3(new_n321), .A4(new_n322), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT29), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n287), .A2(new_n315), .A3(new_n298), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT30), .B1(new_n304), .B2(new_n298), .ZN(new_n338));
  INV_X1    g152(.A(new_n298), .ZN(new_n339));
  OAI21_X1  g153(.A(KEYINPUT67), .B1(new_n275), .B2(new_n278), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n283), .A2(new_n285), .A3(new_n280), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n342), .B2(new_n265), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n338), .B1(new_n343), .B2(KEYINPUT30), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n337), .B1(new_n344), .B2(new_n302), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n335), .B(new_n336), .C1(new_n345), .C2(new_n314), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT68), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n287), .A2(new_n298), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n302), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n350), .A2(KEYINPUT69), .A3(new_n316), .ZN(new_n351));
  OR3_X1    g165(.A1(new_n343), .A2(KEYINPUT69), .A3(new_n315), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(KEYINPUT28), .A3(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT29), .A3(new_n314), .A4(new_n320), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n308), .A2(new_n316), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(new_n324), .ZN(new_n356));
  NAND4_X1  g170(.A1(new_n356), .A2(KEYINPUT68), .A3(new_n336), .A4(new_n335), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n348), .A2(new_n237), .A3(new_n354), .A4(new_n357), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(G472), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n250), .B1(new_n334), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(G478), .ZN(new_n361));
  OR2_X1    g175(.A1(new_n361), .A2(KEYINPUT15), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT13), .ZN(new_n363));
  XNOR2_X1  g177(.A(KEYINPUT64), .B(G143), .ZN(new_n364));
  NOR3_X1   g178(.A1(new_n364), .A2(KEYINPUT88), .A3(new_n187), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT88), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n366), .B1(new_n277), .B2(G128), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n363), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n187), .A2(G143), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT88), .B1(new_n364), .B2(new_n187), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n277), .A2(new_n366), .A3(G128), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G134), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n370), .A2(new_n371), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n375), .A2(new_n257), .A3(new_n369), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(KEYINPUT89), .ZN(new_n377));
  XNOR2_X1  g191(.A(G116), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(G107), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n378), .B(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n375), .A2(new_n257), .A3(new_n369), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT89), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n374), .A2(new_n377), .A3(new_n380), .A4(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(G116), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n385), .A2(KEYINPUT14), .A3(G122), .ZN(new_n386));
  INV_X1    g200(.A(new_n378), .ZN(new_n387));
  OAI211_X1 g201(.A(G107), .B(new_n386), .C1(new_n387), .C2(KEYINPUT14), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n257), .B1(new_n375), .B2(new_n369), .ZN(new_n389));
  OAI221_X1 g203(.A(new_n388), .B1(G107), .B2(new_n387), .C1(new_n376), .C2(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(KEYINPUT9), .B(G234), .Z(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(G217), .A3(new_n232), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n393), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n384), .A2(new_n390), .A3(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(G902), .B1(new_n394), .B2(new_n396), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n362), .B1(new_n397), .B2(KEYINPUT90), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n384), .A2(new_n390), .A3(new_n395), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n395), .B1(new_n384), .B2(new_n390), .ZN(new_n401));
  OAI211_X1 g215(.A(new_n399), .B(new_n237), .C1(new_n400), .C2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT90), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n398), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n403), .A3(new_n362), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT87), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  INV_X1    g223(.A(G104), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(new_n229), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n309), .A2(new_n232), .A3(G214), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n413), .A2(new_n270), .A3(new_n272), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n269), .A2(new_n309), .A3(new_n232), .A4(G214), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n263), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n414), .A2(G131), .A3(new_n415), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(new_n218), .B(KEYINPUT19), .Z(new_n420));
  OAI211_X1 g234(.A(new_n412), .B(new_n419), .C1(G146), .C2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT18), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n416), .B1(new_n422), .B2(new_n263), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n218), .B(new_n219), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n423), .B(new_n424), .C1(new_n422), .C2(new_n418), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n411), .B1(new_n421), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n414), .A2(KEYINPUT17), .A3(G131), .A4(new_n415), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n208), .B1(new_n216), .B2(new_n217), .ZN(new_n428));
  INV_X1    g242(.A(new_n210), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n219), .B1(new_n428), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n427), .A2(new_n430), .A3(new_n211), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT85), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT17), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n417), .A2(new_n434), .A3(new_n418), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n427), .A2(new_n430), .A3(KEYINPUT85), .A4(new_n211), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n437), .A2(new_n411), .A3(new_n425), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT86), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n437), .A2(KEYINPUT86), .A3(new_n411), .A4(new_n425), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n426), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  NOR3_X1   g256(.A1(new_n442), .A2(G475), .A3(G902), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n408), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n440), .A2(new_n441), .ZN(new_n446));
  INV_X1    g260(.A(new_n426), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(G475), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n448), .A2(new_n449), .A3(new_n237), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(KEYINPUT87), .A3(KEYINPUT20), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n443), .A2(new_n444), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n411), .B1(new_n437), .B2(new_n425), .ZN(new_n454));
  AOI21_X1  g268(.A(new_n454), .B1(new_n440), .B2(new_n441), .ZN(new_n455));
  OAI21_X1  g269(.A(G475), .B1(new_n455), .B2(G902), .ZN(new_n456));
  XOR2_X1   g270(.A(KEYINPUT21), .B(G898), .Z(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT92), .ZN(new_n458));
  AOI211_X1 g272(.A(new_n237), .B(new_n232), .C1(G234), .C2(G237), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(G952), .ZN(new_n461));
  AOI211_X1 g275(.A(G953), .B(new_n461), .C1(G234), .C2(G237), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  AND4_X1   g278(.A1(new_n407), .A2(new_n453), .A3(new_n456), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n360), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(KEYINPUT3), .B1(new_n410), .B2(G107), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT3), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(new_n379), .A3(G104), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n410), .A2(G107), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT4), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n474), .A3(G101), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT76), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT76), .ZN(new_n477));
  NAND4_X1  g291(.A1(new_n473), .A2(new_n477), .A3(new_n474), .A4(G101), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n473), .A2(G101), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n469), .A2(new_n471), .A3(new_n311), .A4(new_n472), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(KEYINPUT4), .A3(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT75), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n480), .A2(KEYINPUT75), .A3(KEYINPUT4), .A4(new_n481), .ZN(new_n485));
  NAND4_X1  g299(.A1(new_n479), .A2(new_n484), .A3(new_n302), .A4(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT77), .B1(new_n410), .B2(G107), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT77), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n488), .A2(new_n379), .A3(G104), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n487), .A2(new_n489), .A3(new_n472), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G101), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n491), .A2(new_n481), .ZN(new_n492));
  INV_X1    g306(.A(new_n300), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT5), .ZN(new_n494));
  INV_X1    g308(.A(G113), .ZN(new_n495));
  NOR2_X1   g309(.A1(KEYINPUT5), .A2(G119), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n495), .B1(new_n496), .B2(G116), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n300), .A2(new_n301), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n492), .A2(new_n498), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n486), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(G110), .B(G122), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT79), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT80), .ZN(new_n506));
  INV_X1    g320(.A(new_n504), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n486), .A2(new_n507), .A3(new_n501), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(new_n486), .B2(new_n501), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT80), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n506), .A2(new_n508), .A3(KEYINPUT6), .A4(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT81), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT6), .ZN(new_n514));
  AND4_X1   g328(.A1(new_n513), .A2(new_n502), .A3(new_n514), .A4(new_n504), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n513), .B1(new_n509), .B2(new_n514), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n303), .A2(G125), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n296), .A2(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n281), .A2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n293), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n295), .B(new_n521), .C1(new_n364), .C2(new_n219), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n215), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n232), .A2(G224), .ZN(new_n526));
  XOR2_X1   g340(.A(new_n526), .B(KEYINPUT82), .Z(new_n527));
  XNOR2_X1  g341(.A(new_n525), .B(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n512), .A2(new_n517), .A3(new_n528), .ZN(new_n529));
  AOI22_X1  g343(.A1(new_n518), .A2(new_n524), .B1(KEYINPUT84), .B2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(KEYINPUT7), .ZN(new_n531));
  XNOR2_X1  g345(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XOR2_X1   g346(.A(new_n504), .B(KEYINPUT8), .Z(new_n533));
  NAND2_X1  g347(.A1(new_n491), .A2(new_n481), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n497), .B(KEYINPUT83), .Z(new_n535));
  AOI211_X1 g349(.A(new_n499), .B(new_n534), .C1(new_n535), .C2(new_n494), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n492), .B1(new_n500), .B2(new_n498), .ZN(new_n537));
  OAI21_X1  g351(.A(new_n533), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n532), .A2(new_n508), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n529), .A2(new_n539), .A3(new_n237), .ZN(new_n540));
  OAI21_X1  g354(.A(G210), .B1(G237), .B2(G902), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n529), .A2(new_n539), .A3(new_n237), .A4(new_n541), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n468), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(G221), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n392), .B2(new_n237), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT74), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND4_X1  g363(.A1(new_n342), .A2(new_n479), .A3(new_n484), .A4(new_n485), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n187), .B1(new_n273), .B2(KEYINPUT1), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n522), .B1(new_n551), .B2(new_n284), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n492), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT10), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n523), .A2(new_n492), .A3(KEYINPUT10), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n265), .B(KEYINPUT78), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n550), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(G110), .B(G140), .ZN(new_n559));
  INV_X1    g373(.A(G227), .ZN(new_n560));
  NOR2_X1   g374(.A1(new_n560), .A2(G953), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n559), .B(new_n561), .Z(new_n562));
  AND2_X1   g376(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n279), .A2(new_n286), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n479), .A2(new_n484), .A3(new_n485), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n555), .B(new_n556), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n265), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n523), .A2(new_n492), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n295), .B1(new_n364), .B2(new_n219), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n292), .B1(new_n364), .B2(new_n219), .ZN(new_n570));
  OAI21_X1  g384(.A(new_n569), .B1(new_n570), .B2(new_n187), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n534), .B1(new_n571), .B2(new_n522), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n265), .B1(new_n568), .B2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT12), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  OAI211_X1 g389(.A(KEYINPUT12), .B(new_n265), .C1(new_n568), .C2(new_n572), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(new_n558), .ZN(new_n578));
  INV_X1    g392(.A(new_n562), .ZN(new_n579));
  AOI22_X1  g393(.A1(new_n563), .A2(new_n567), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G469), .B1(new_n580), .B2(G902), .ZN(new_n581));
  INV_X1    g395(.A(G469), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n577), .A2(new_n558), .A3(new_n562), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n562), .B1(new_n567), .B2(new_n558), .ZN(new_n584));
  OAI211_X1 g398(.A(new_n582), .B(new_n237), .C1(new_n583), .C2(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n549), .B1(new_n581), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n545), .A2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n466), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(new_n311), .ZN(G3));
  INV_X1    g403(.A(new_n250), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n328), .A2(new_n237), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G472), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n586), .A2(new_n330), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(KEYINPUT93), .ZN(new_n594));
  INV_X1    g408(.A(new_n330), .ZN(new_n595));
  INV_X1    g409(.A(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n596), .B1(new_n328), .B2(new_n237), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT93), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n598), .A2(new_n599), .A3(new_n590), .A4(new_n586), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n594), .A2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n601), .B(KEYINPUT94), .ZN(new_n602));
  INV_X1    g416(.A(new_n545), .ZN(new_n603));
  INV_X1    g417(.A(new_n464), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT33), .B1(new_n400), .B2(new_n401), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT33), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n394), .A2(new_n606), .A3(new_n396), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n605), .A2(new_n607), .A3(G478), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n397), .A2(new_n361), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n361), .A2(new_n237), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  AOI211_X1 g426(.A(new_n604), .B(new_n612), .C1(new_n453), .C2(new_n456), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n602), .A2(new_n603), .A3(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT34), .B(G104), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G6));
  INV_X1    g431(.A(new_n602), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n445), .A2(new_n451), .A3(KEYINPUT95), .ZN(new_n619));
  AOI21_X1  g433(.A(KEYINPUT95), .B1(new_n445), .B2(new_n451), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n452), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  AND3_X1   g435(.A1(new_n402), .A2(new_n403), .A3(new_n362), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n622), .B1(new_n404), .B2(new_n398), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n464), .B(KEYINPUT96), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n621), .A2(new_n623), .A3(new_n456), .A4(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(KEYINPUT97), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n445), .A2(new_n451), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT95), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n445), .A2(new_n451), .A3(KEYINPUT95), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n407), .B1(new_n631), .B2(new_n452), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT97), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n456), .A4(new_n624), .ZN(new_n634));
  AND4_X1   g448(.A1(new_n545), .A2(new_n618), .A3(new_n626), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(new_n379), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT98), .B(KEYINPUT35), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G9));
  INV_X1    g452(.A(new_n585), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n578), .A2(new_n579), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n567), .A2(new_n558), .A3(new_n562), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n640), .A2(G469), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(G469), .A2(G902), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n548), .B1(new_n639), .B2(new_n644), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n645), .A2(new_n595), .A3(new_n597), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT36), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n234), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(new_n230), .Z(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n237), .C1(new_n243), .C2(G234), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n248), .A2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT100), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n248), .A2(new_n651), .A3(KEYINPUT100), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n465), .A2(new_n646), .A3(new_n545), .A4(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G110), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  NAND2_X1  g474(.A1(new_n545), .A2(new_n656), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n331), .A2(new_n333), .B1(new_n358), .B2(G472), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n661), .A2(new_n662), .A3(new_n645), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n462), .B1(new_n459), .B2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n456), .A2(new_n666), .ZN(new_n667));
  AND3_X1   g481(.A1(new_n621), .A2(new_n623), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n663), .A2(new_n668), .A3(KEYINPUT102), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT102), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n334), .A2(new_n359), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n671), .A2(new_n545), .A3(new_n586), .A4(new_n656), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n621), .A2(new_n623), .A3(new_n667), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT103), .B(G128), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(G30));
  NAND2_X1  g491(.A1(new_n543), .A2(new_n544), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT38), .ZN(new_n679));
  INV_X1    g493(.A(new_n652), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n453), .A2(new_n456), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n623), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n665), .B(KEYINPUT39), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n645), .A2(new_n684), .ZN(new_n685));
  OR2_X1    g499(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n685), .A2(KEYINPUT40), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n683), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n355), .A2(new_n314), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n237), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n314), .B1(new_n351), .B2(new_n352), .ZN(new_n691));
  OAI21_X1  g505(.A(G472), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n334), .A2(new_n692), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n681), .A2(new_n688), .A3(new_n467), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(new_n364), .ZN(G45));
  AOI21_X1  g509(.A(new_n645), .B1(new_n334), .B2(new_n359), .ZN(new_n696));
  AOI221_X4 g510(.A(new_n468), .B1(new_n654), .B2(new_n655), .C1(new_n543), .C2(new_n544), .ZN(new_n697));
  AOI211_X1 g511(.A(new_n612), .B(new_n665), .C1(new_n453), .C2(new_n456), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  OAI21_X1  g514(.A(new_n237), .B1(new_n583), .B2(new_n584), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n701), .A2(G469), .ZN(new_n702));
  INV_X1    g516(.A(new_n547), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n703), .A3(new_n585), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT104), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n360), .A2(new_n706), .A3(new_n545), .A4(new_n613), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  NAND2_X1  g523(.A1(new_n671), .A2(new_n590), .ZN(new_n710));
  OR2_X1    g524(.A1(new_n704), .A2(KEYINPUT104), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n704), .A2(KEYINPUT104), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n711), .A2(new_n545), .A3(new_n712), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n710), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n634), .A2(new_n626), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  NAND4_X1  g530(.A1(new_n706), .A2(new_n697), .A3(new_n671), .A4(new_n465), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(new_n329), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n353), .A2(new_n320), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n324), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n318), .A2(new_n327), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NOR3_X1   g537(.A1(new_n723), .A2(new_n597), .A3(new_n250), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n724), .B(new_n725), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n682), .A2(new_n623), .A3(new_n624), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n726), .A2(new_n545), .A3(new_n706), .A4(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G122), .ZN(G24));
  NOR3_X1   g543(.A1(new_n723), .A2(new_n597), .A3(new_n680), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n706), .A2(new_n698), .A3(new_n545), .A4(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G125), .ZN(G27));
  AOI21_X1  g546(.A(new_n547), .B1(new_n581), .B2(new_n585), .ZN(new_n733));
  AND4_X1   g547(.A1(new_n467), .A2(new_n733), .A3(new_n543), .A4(new_n544), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(new_n698), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n710), .A2(KEYINPUT107), .ZN(new_n738));
  OAI211_X1 g552(.A(KEYINPUT42), .B(new_n736), .C1(new_n737), .C2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT106), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n735), .B2(new_n710), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT42), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n734), .A2(new_n360), .A3(KEYINPUT106), .A4(new_n698), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n741), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n739), .A2(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(new_n263), .ZN(G33));
  NAND3_X1  g560(.A1(new_n668), .A2(new_n360), .A3(new_n734), .ZN(new_n747));
  XNOR2_X1  g561(.A(KEYINPUT108), .B(G134), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n747), .B(new_n748), .ZN(G36));
  INV_X1    g563(.A(new_n598), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n453), .A2(new_n456), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  AOI21_X1  g566(.A(KEYINPUT43), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  INV_X1    g567(.A(new_n612), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n753), .A2(new_n755), .ZN(new_n758));
  OAI211_X1 g572(.A(new_n750), .B(new_n652), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT44), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n753), .A2(new_n755), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n756), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n763), .A2(KEYINPUT44), .A3(new_n750), .A4(new_n652), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n678), .A2(new_n468), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n580), .A2(KEYINPUT45), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n580), .A2(KEYINPUT45), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n766), .A2(G469), .A3(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n768), .B2(new_n643), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n769), .A2(new_n639), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(KEYINPUT46), .A3(new_n643), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n547), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n684), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n761), .A2(new_n764), .A3(new_n765), .A4(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NOR2_X1   g590(.A1(new_n671), .A2(new_n590), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n698), .A2(new_n765), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n772), .A2(KEYINPUT47), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT47), .ZN(new_n780));
  AOI211_X1 g594(.A(new_n780), .B(new_n547), .C1(new_n770), .C2(new_n771), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n777), .B(new_n778), .C1(new_n779), .C2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(KEYINPUT110), .B(G140), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n782), .B(new_n783), .ZN(G42));
  AOI21_X1  g598(.A(new_n463), .B1(new_n762), .B2(new_n756), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(new_n468), .A3(new_n706), .A4(new_n726), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n787));
  OR3_X1    g601(.A1(new_n786), .A2(new_n787), .A3(new_n679), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n787), .B1(new_n786), .B2(new_n679), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n726), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n468), .A3(new_n678), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n779), .A2(new_n781), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n702), .A2(new_n585), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n793), .A2(new_n548), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT115), .Z(new_n795));
  OR2_X1    g609(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  AOI22_X1  g610(.A1(new_n788), .A2(new_n789), .B1(new_n791), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n706), .A2(new_n765), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT116), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n801), .A2(new_n785), .ZN(new_n802));
  INV_X1    g616(.A(new_n730), .ZN(new_n803));
  INV_X1    g617(.A(new_n693), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n590), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n799), .A2(new_n462), .A3(new_n800), .A4(new_n806), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n682), .A2(new_n754), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  OAI22_X1  g623(.A1(new_n802), .A2(new_n803), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  INV_X1    g624(.A(new_n810), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT51), .B1(new_n797), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n791), .B1(new_n792), .B2(new_n794), .ZN(new_n813));
  OR2_X1    g627(.A1(new_n810), .A2(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n788), .A2(new_n789), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n816), .B1(new_n810), .B2(KEYINPUT117), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n812), .B1(new_n813), .B2(new_n818), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n790), .A2(KEYINPUT118), .A3(new_n713), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT118), .B1(new_n790), .B2(new_n713), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n461), .A2(G953), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n710), .B(KEYINPUT107), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n801), .A2(new_n824), .A3(new_n785), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT48), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT48), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n801), .A2(new_n827), .A3(new_n824), .A4(new_n785), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n612), .B1(new_n453), .B2(new_n456), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n801), .A2(new_n462), .A3(new_n830), .A4(new_n806), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n822), .A2(new_n823), .A3(new_n829), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT119), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n832), .B(new_n833), .ZN(new_n834));
  AND2_X1   g648(.A1(new_n731), .A2(new_n699), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n603), .A2(new_n683), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n652), .A2(new_n665), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n836), .A2(new_n693), .A3(new_n733), .A4(new_n837), .ZN(new_n838));
  AOI21_X1  g652(.A(KEYINPUT102), .B1(new_n663), .B2(new_n668), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n672), .A2(new_n673), .A3(new_n670), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n835), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n675), .A2(KEYINPUT52), .A3(new_n835), .A4(new_n838), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n745), .B1(new_n843), .B2(new_n844), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n623), .A2(new_n453), .A3(new_n456), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n545), .B(new_n624), .C1(new_n846), .C2(new_n830), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n601), .A2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n657), .B1(new_n466), .B2(new_n587), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g664(.A1(new_n407), .A2(new_n667), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n765), .A2(new_n621), .A3(new_n851), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT113), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT113), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n765), .A2(new_n621), .A3(new_n854), .A4(new_n851), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n853), .A2(new_n656), .A3(new_n696), .A4(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n736), .A2(new_n730), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n850), .A2(new_n747), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n707), .A2(new_n717), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n715), .A2(new_n859), .A3(new_n728), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n715), .A2(new_n859), .A3(new_n728), .A4(KEYINPUT112), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n858), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n845), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n843), .A2(new_n844), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT114), .ZN(new_n867));
  AOI21_X1  g681(.A(KEYINPUT53), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g683(.A(KEYINPUT114), .B1(new_n843), .B2(new_n844), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n845), .B(new_n864), .C1(new_n870), .C2(KEYINPUT53), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT54), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n865), .A2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT54), .ZN(new_n876));
  INV_X1    g690(.A(new_n860), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n858), .A2(new_n874), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n845), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n819), .A2(new_n834), .A3(new_n873), .A4(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n461), .A2(new_n232), .ZN(new_n882));
  XNOR2_X1  g696(.A(new_n882), .B(KEYINPUT120), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR4_X1   g698(.A1(new_n755), .A2(new_n250), .A3(new_n468), .A4(new_n549), .ZN(new_n885));
  XNOR2_X1  g699(.A(new_n885), .B(KEYINPUT111), .ZN(new_n886));
  OR2_X1    g700(.A1(new_n793), .A2(KEYINPUT49), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n679), .B1(KEYINPUT49), .B2(new_n793), .ZN(new_n888));
  NAND4_X1  g702(.A1(new_n886), .A2(new_n804), .A3(new_n887), .A4(new_n888), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n884), .A2(new_n889), .ZN(G75));
  NAND2_X1  g704(.A1(new_n875), .A2(new_n879), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n891), .A2(G210), .A3(G902), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT56), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n892), .A2(KEYINPUT121), .A3(new_n893), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n512), .A2(new_n517), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n528), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT55), .Z(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n232), .A2(G952), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n892), .A2(KEYINPUT121), .A3(new_n893), .A4(new_n897), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(G51));
  INV_X1    g717(.A(new_n768), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n891), .A2(G902), .A3(new_n904), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT122), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n905), .B(new_n906), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n643), .B(KEYINPUT57), .Z(new_n908));
  AND3_X1   g722(.A1(new_n875), .A2(new_n876), .A3(new_n879), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n876), .B1(new_n875), .B2(new_n879), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n908), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n911), .B1(new_n584), .B2(new_n583), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n900), .B1(new_n907), .B2(new_n912), .ZN(G54));
  AOI21_X1  g727(.A(new_n237), .B1(new_n875), .B2(new_n879), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n914), .A2(KEYINPUT58), .A3(G475), .ZN(new_n915));
  AND2_X1   g729(.A1(new_n915), .A2(new_n442), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n442), .ZN(new_n917));
  NOR3_X1   g731(.A1(new_n916), .A2(new_n917), .A3(new_n900), .ZN(G60));
  NAND2_X1  g732(.A1(new_n605), .A2(new_n607), .ZN(new_n919));
  XNOR2_X1  g733(.A(KEYINPUT123), .B(KEYINPUT59), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n611), .B(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n919), .B(new_n922), .C1(new_n909), .C2(new_n910), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(new_n901), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT124), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n921), .B1(new_n873), .B2(new_n880), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n925), .B1(new_n926), .B2(new_n919), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n876), .B1(new_n869), .B2(new_n871), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n922), .B1(new_n909), .B2(new_n928), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n929), .A2(KEYINPUT124), .A3(new_n605), .A4(new_n607), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n924), .B1(new_n927), .B2(new_n930), .ZN(G63));
  NAND2_X1  g745(.A1(G217), .A2(G902), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT60), .Z(new_n933));
  NAND2_X1  g747(.A1(new_n891), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n236), .A2(new_n238), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n891), .A2(new_n650), .A3(new_n933), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n936), .A2(new_n901), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT61), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n936), .A2(KEYINPUT61), .A3(new_n901), .A4(new_n937), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(G66));
  INV_X1    g756(.A(G224), .ZN(new_n943));
  OAI21_X1  g757(.A(G953), .B1(new_n458), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n862), .A2(new_n863), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n946));
  AND3_X1   g760(.A1(new_n945), .A2(new_n946), .A3(new_n850), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n946), .B1(new_n945), .B2(new_n850), .ZN(new_n948));
  OR2_X1    g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n944), .B1(new_n949), .B2(G953), .ZN(new_n950));
  INV_X1    g764(.A(G898), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n895), .B1(new_n951), .B2(G953), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n950), .B(new_n952), .Z(G69));
  NAND3_X1  g767(.A1(new_n694), .A2(new_n675), .A3(new_n835), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT62), .ZN(new_n955));
  OR2_X1    g769(.A1(new_n846), .A2(new_n830), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n360), .A2(new_n956), .A3(new_n685), .A4(new_n765), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n954), .B2(KEYINPUT62), .ZN(new_n958));
  AND4_X1   g772(.A1(new_n775), .A2(new_n955), .A3(new_n782), .A4(new_n958), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(G953), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n344), .B(new_n420), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(G953), .B1(new_n560), .B2(new_n664), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n664), .B2(G227), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n775), .A2(new_n747), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n774), .A2(new_n824), .A3(new_n836), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT126), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n774), .A2(new_n968), .A3(new_n824), .A4(new_n836), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n782), .A2(new_n675), .A3(new_n835), .ZN(new_n971));
  NOR4_X1   g785(.A1(new_n965), .A2(new_n970), .A3(new_n745), .A4(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n961), .B1(new_n972), .B2(new_n232), .ZN(new_n973));
  AOI22_X1  g787(.A1(new_n962), .A2(new_n963), .B1(new_n964), .B2(new_n973), .ZN(G72));
  OAI21_X1  g788(.A(new_n972), .B1(new_n948), .B2(new_n947), .ZN(new_n975));
  NAND2_X1  g789(.A1(G472), .A2(G902), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT63), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n355), .A2(new_n314), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n900), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n872), .A2(new_n689), .A3(new_n977), .A4(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n959), .B1(new_n947), .B2(new_n948), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n689), .B1(new_n983), .B2(new_n977), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT127), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI211_X1 g800(.A(KEYINPUT127), .B(new_n689), .C1(new_n983), .C2(new_n977), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n980), .B(new_n982), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(G57));
endmodule


