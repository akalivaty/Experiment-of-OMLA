//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 0 1 0 0 1 1 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 1 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:11 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932;
  XNOR2_X1  g000(.A(G110), .B(G122), .ZN(new_n187));
  XOR2_X1   g001(.A(new_n187), .B(KEYINPUT78), .Z(new_n188));
  XNOR2_X1  g002(.A(G116), .B(G119), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT2), .B(G113), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT71), .ZN(new_n192));
  INV_X1    g006(.A(G107), .ZN(new_n193));
  OAI22_X1  g007(.A1(new_n192), .A2(KEYINPUT3), .B1(new_n193), .B2(G104), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT3), .ZN(new_n195));
  INV_X1    g009(.A(G104), .ZN(new_n196));
  OAI22_X1  g010(.A1(KEYINPUT71), .A2(new_n195), .B1(new_n196), .B2(G107), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT3), .A4(G104), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n194), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT4), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n191), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI22_X1  g017(.A1(KEYINPUT71), .A2(new_n195), .B1(new_n196), .B2(G107), .ZN(new_n204));
  AND4_X1   g018(.A1(new_n192), .A2(new_n193), .A3(KEYINPUT3), .A4(G104), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n192), .A2(KEYINPUT3), .B1(new_n193), .B2(G104), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n200), .B(new_n204), .C1(new_n205), .C2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT72), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n197), .A2(new_n198), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n210), .A2(KEYINPUT72), .A3(new_n200), .A4(new_n204), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT73), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n210), .A2(new_n204), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n202), .B1(new_n214), .B2(G101), .ZN(new_n215));
  AND3_X1   g029(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n213), .B1(new_n212), .B2(new_n215), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n203), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT76), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n193), .A2(G104), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n196), .A2(G107), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n200), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n222), .B1(new_n209), .B2(new_n211), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n189), .A2(KEYINPUT5), .ZN(new_n224));
  INV_X1    g038(.A(G116), .ZN(new_n225));
  NOR3_X1   g039(.A1(new_n225), .A2(KEYINPUT5), .A3(G119), .ZN(new_n226));
  INV_X1    g040(.A(G113), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(new_n190), .ZN(new_n229));
  AOI22_X1  g043(.A1(new_n224), .A2(new_n228), .B1(new_n229), .B2(new_n189), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n223), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT76), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n232), .B(new_n203), .C1(new_n216), .C2(new_n217), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n219), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT77), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n188), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT6), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n219), .A2(KEYINPUT77), .A3(new_n231), .A4(new_n233), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n236), .A2(KEYINPUT80), .A3(new_n237), .A4(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n233), .A2(new_n231), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT72), .B1(new_n199), .B2(new_n200), .ZN(new_n241));
  AND4_X1   g055(.A1(KEYINPUT72), .A2(new_n210), .A3(new_n200), .A4(new_n204), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n215), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(KEYINPUT73), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n232), .B1(new_n246), .B2(new_n203), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n235), .B1(new_n240), .B2(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(new_n188), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n248), .A2(new_n238), .A3(new_n237), .A4(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT80), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n239), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n248), .A2(new_n238), .A3(new_n249), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT79), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n248), .A2(new_n238), .A3(KEYINPUT79), .A4(new_n249), .ZN(new_n257));
  INV_X1    g071(.A(new_n187), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n234), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n259), .A2(new_n237), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n257), .A3(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G143), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(G146), .ZN(new_n263));
  INV_X1    g077(.A(KEYINPUT64), .ZN(new_n264));
  INV_X1    g078(.A(G146), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n264), .B1(new_n265), .B2(G143), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n262), .A2(KEYINPUT64), .A3(G146), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n263), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT1), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n268), .A2(new_n269), .A3(G128), .ZN(new_n270));
  OAI21_X1  g084(.A(G128), .B1(new_n263), .B2(new_n269), .ZN(new_n271));
  XOR2_X1   g085(.A(G143), .B(G146), .Z(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(G125), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  XOR2_X1   g092(.A(KEYINPUT0), .B(G128), .Z(new_n279));
  AOI22_X1  g093(.A1(new_n268), .A2(new_n278), .B1(new_n279), .B2(new_n272), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n277), .B1(new_n276), .B2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G224), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n282), .A2(G953), .ZN(new_n283));
  XNOR2_X1  g097(.A(new_n283), .B(KEYINPUT81), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n281), .B(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n253), .A2(new_n261), .A3(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n259), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT84), .B1(new_n280), .B2(new_n276), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT7), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n289), .B2(new_n284), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n281), .B(new_n290), .Z(new_n291));
  INV_X1    g105(.A(new_n223), .ZN(new_n292));
  OAI211_X1 g106(.A(KEYINPUT83), .B(new_n230), .C1(new_n292), .C2(KEYINPUT82), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n187), .B(KEYINPUT8), .Z(new_n294));
  OAI21_X1  g108(.A(KEYINPUT83), .B1(new_n292), .B2(KEYINPUT82), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT83), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n230), .B1(new_n223), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n294), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n291), .B1(new_n293), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G902), .B1(new_n287), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n286), .A2(new_n300), .ZN(new_n301));
  OAI21_X1  g115(.A(G210), .B1(G237), .B2(G902), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n286), .A2(new_n300), .A3(new_n302), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT11), .ZN(new_n307));
  INV_X1    g121(.A(G134), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n307), .B1(new_n308), .B2(G137), .ZN(new_n309));
  INV_X1    g123(.A(G137), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n310), .A2(KEYINPUT11), .A3(G134), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(G137), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  OR2_X1    g127(.A1(new_n313), .A2(G131), .ZN(new_n314));
  INV_X1    g128(.A(new_n312), .ZN(new_n315));
  NOR2_X1   g129(.A1(new_n308), .A2(G137), .ZN(new_n316));
  OAI21_X1  g130(.A(G131), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n274), .A2(new_n314), .A3(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(new_n313), .B(G131), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n280), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT65), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT30), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n326));
  INV_X1    g140(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n318), .A2(new_n320), .A3(new_n322), .A4(new_n323), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n191), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n318), .A2(new_n320), .A3(new_n191), .ZN(new_n332));
  XOR2_X1   g146(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n333));
  NOR2_X1   g147(.A1(G237), .A2(G953), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G210), .ZN(new_n335));
  XNOR2_X1  g149(.A(new_n333), .B(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(KEYINPUT26), .B(G101), .ZN(new_n337));
  XNOR2_X1  g151(.A(new_n336), .B(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n331), .A2(new_n332), .A3(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT31), .ZN(new_n340));
  INV_X1    g154(.A(new_n338), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n342));
  INV_X1    g156(.A(new_n191), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n321), .A2(new_n343), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n342), .B1(new_n344), .B2(new_n332), .ZN(new_n345));
  INV_X1    g159(.A(new_n332), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n346), .A2(KEYINPUT28), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n341), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n339), .A2(new_n340), .A3(new_n348), .ZN(new_n349));
  NOR3_X1   g163(.A1(new_n330), .A2(new_n346), .A3(new_n341), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n350), .B2(KEYINPUT31), .ZN(new_n351));
  INV_X1    g165(.A(G472), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n353), .A2(KEYINPUT32), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT32), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n349), .A2(new_n351), .A3(new_n355), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  OR3_X1    g171(.A1(new_n345), .A2(new_n347), .A3(new_n341), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT29), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n330), .A2(new_n346), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n338), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n360), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(G902), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n364), .B1(new_n358), .B2(new_n359), .ZN(new_n365));
  OAI21_X1  g179(.A(G472), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT16), .ZN(new_n368));
  INV_X1    g182(.A(G140), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(G125), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n276), .A2(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n370), .B1(new_n373), .B2(new_n368), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(new_n265), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n265), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(G119), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G128), .ZN(new_n380));
  NAND2_X1  g194(.A1(KEYINPUT23), .A2(G119), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n379), .A2(G128), .ZN(new_n382));
  OAI221_X1 g196(.A(new_n380), .B1(G128), .B2(new_n381), .C1(new_n382), .C2(KEYINPUT23), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT68), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n384), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(G110), .A3(new_n386), .ZN(new_n387));
  OR3_X1    g201(.A1(new_n379), .A2(KEYINPUT67), .A3(G128), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT67), .B1(new_n379), .B2(G128), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n380), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT24), .B(G110), .ZN(new_n391));
  OR2_X1    g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n378), .A2(new_n387), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  OAI21_X1  g208(.A(new_n394), .B1(G110), .B2(new_n383), .ZN(new_n395));
  INV_X1    g209(.A(new_n373), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n265), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n376), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(G953), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(G221), .A3(G234), .ZN(new_n400));
  XNOR2_X1  g214(.A(new_n400), .B(KEYINPUT69), .ZN(new_n401));
  XNOR2_X1  g215(.A(KEYINPUT22), .B(G137), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n401), .B(new_n402), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n393), .A2(new_n398), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n403), .B1(new_n393), .B2(new_n398), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  OAI21_X1  g221(.A(KEYINPUT70), .B1(new_n407), .B2(G902), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT25), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI211_X1 g224(.A(KEYINPUT70), .B(KEYINPUT25), .C1(new_n407), .C2(G902), .ZN(new_n411));
  INV_X1    g225(.A(G217), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(G234), .B2(new_n364), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n410), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n407), .ZN(new_n415));
  NOR2_X1   g229(.A1(new_n413), .A2(G902), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n414), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n367), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g234(.A(G214), .B1(G237), .B2(G902), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT20), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n334), .A2(G143), .A3(G214), .ZN(new_n423));
  AOI21_X1  g237(.A(G143), .B1(new_n334), .B2(G214), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(G131), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT17), .ZN(new_n427));
  AND2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(KEYINPUT17), .B(G131), .C1(new_n423), .C2(new_n424), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n376), .A2(new_n377), .A3(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(G113), .B(G122), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n433), .B(new_n196), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n434), .B(KEYINPUT90), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(KEYINPUT18), .A2(G131), .ZN(new_n437));
  XOR2_X1   g251(.A(new_n425), .B(new_n437), .Z(new_n438));
  NAND2_X1  g252(.A1(new_n396), .A2(KEYINPUT85), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT85), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n373), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n439), .A2(G146), .A3(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n442), .A2(new_n443), .A3(new_n397), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n443), .B1(new_n442), .B2(new_n397), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n438), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT87), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n446), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(new_n444), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT87), .B1(new_n451), .B2(new_n438), .ZN(new_n452));
  OAI211_X1 g266(.A(new_n432), .B(new_n436), .C1(new_n449), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n447), .A2(new_n448), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(KEYINPUT87), .A3(new_n438), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n439), .A2(KEYINPUT19), .A3(new_n441), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT88), .ZN(new_n457));
  OR2_X1    g271(.A1(new_n457), .A2(KEYINPUT19), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(KEYINPUT19), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n396), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n456), .A2(new_n265), .A3(new_n460), .ZN(new_n461));
  XNOR2_X1  g275(.A(new_n461), .B(KEYINPUT89), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n426), .A2(new_n375), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n454), .A2(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n453), .B1(new_n434), .B2(new_n464), .ZN(new_n465));
  NOR2_X1   g279(.A1(G475), .A2(G902), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n422), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n465), .A2(new_n422), .A3(new_n466), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n431), .B1(new_n454), .B2(new_n455), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n470), .A2(new_n434), .ZN(new_n471));
  AOI211_X1 g285(.A(new_n435), .B(new_n431), .C1(new_n454), .C2(new_n455), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n364), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI22_X1  g287(.A1(new_n468), .A2(new_n469), .B1(G475), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n399), .A2(G952), .ZN(new_n475));
  INV_X1    g289(.A(G234), .ZN(new_n476));
  INV_X1    g290(.A(G237), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI211_X1 g293(.A(new_n364), .B(new_n399), .C1(G234), .C2(G237), .ZN(new_n480));
  XNOR2_X1  g294(.A(KEYINPUT21), .B(G898), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  INV_X1    g296(.A(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT9), .B(G234), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n484), .A2(new_n412), .A3(G953), .ZN(new_n485));
  XNOR2_X1  g299(.A(G116), .B(G122), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT14), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n225), .A2(KEYINPUT14), .A3(G122), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n488), .A2(G107), .A3(new_n489), .ZN(new_n490));
  XOR2_X1   g304(.A(new_n490), .B(KEYINPUT93), .Z(new_n491));
  NAND2_X1  g305(.A1(new_n486), .A2(new_n193), .ZN(new_n492));
  XNOR2_X1  g306(.A(G128), .B(G143), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G134), .ZN(new_n494));
  INV_X1    g308(.A(new_n493), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n495), .A2(new_n308), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n491), .A2(new_n492), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n486), .B(G107), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT91), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n500));
  OAI22_X1  g314(.A1(new_n500), .A2(KEYINPUT13), .B1(new_n262), .B2(G128), .ZN(new_n501));
  AND2_X1   g315(.A1(new_n500), .A2(KEYINPUT13), .ZN(new_n502));
  OAI21_X1  g316(.A(G134), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n495), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n499), .A2(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n485), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n497), .A2(new_n505), .A3(new_n485), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n364), .ZN(new_n510));
  INV_X1    g324(.A(G478), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  AOI21_X1  g327(.A(G902), .B1(new_n507), .B2(new_n508), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n514), .B1(KEYINPUT15), .B2(new_n511), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n474), .A2(new_n483), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(G469), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n201), .A2(new_n202), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n520), .A2(new_n280), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n246), .A2(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(new_n319), .ZN(new_n523));
  INV_X1    g337(.A(new_n222), .ZN(new_n524));
  INV_X1    g338(.A(new_n271), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n270), .B1(new_n268), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n212), .A2(new_n524), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT10), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n223), .A2(KEYINPUT10), .A3(new_n274), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n522), .A2(new_n523), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(G110), .B(G140), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n399), .A2(G227), .ZN(new_n533));
  XOR2_X1   g347(.A(new_n532), .B(new_n533), .Z(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n274), .B1(new_n212), .B2(new_n524), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT74), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n523), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  OAI211_X1 g353(.A(new_n527), .B(KEYINPUT74), .C1(new_n274), .C2(new_n223), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT12), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT75), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(KEYINPUT12), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT12), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n544), .B1(new_n545), .B2(KEYINPUT75), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n536), .B1(new_n543), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n246), .A2(new_n521), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n529), .A2(new_n530), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n319), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n535), .B1(new_n550), .B2(new_n531), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n519), .B(new_n364), .C1(new_n547), .C2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n536), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n550), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n548), .A2(new_n319), .A3(new_n549), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n555), .B1(new_n546), .B2(new_n543), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n554), .B(G469), .C1(new_n556), .C2(new_n535), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n519), .A2(new_n364), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n552), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g374(.A(G221), .B1(new_n484), .B2(G902), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n518), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g377(.A1(new_n306), .A2(new_n420), .A3(new_n421), .A4(new_n563), .ZN(new_n564));
  XNOR2_X1  g378(.A(new_n564), .B(G101), .ZN(G3));
  INV_X1    g379(.A(KEYINPUT94), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n566), .B1(new_n306), .B2(new_n421), .ZN(new_n567));
  AND3_X1   g381(.A1(new_n286), .A2(new_n300), .A3(new_n302), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n302), .B1(new_n286), .B2(new_n300), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n566), .B(new_n421), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n349), .A2(new_n351), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(G472), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n353), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n577), .A2(new_n560), .A3(new_n418), .A4(new_n561), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n509), .A2(KEYINPUT33), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n509), .A2(KEYINPUT33), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(G478), .A3(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n511), .A2(new_n364), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n583), .B1(new_n514), .B2(new_n511), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n582), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n473), .A2(G475), .ZN(new_n587));
  AND3_X1   g401(.A1(new_n465), .A2(new_n422), .A3(new_n466), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n587), .B1(new_n588), .B2(new_n467), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(new_n482), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n573), .A2(new_n579), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n592), .B(KEYINPUT95), .Z(new_n593));
  XOR2_X1   g407(.A(KEYINPUT34), .B(G104), .Z(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G6));
  OAI211_X1 g409(.A(new_n516), .B(new_n587), .C1(new_n588), .C2(new_n467), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n482), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n573), .A2(new_n579), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  NAND2_X1  g414(.A1(new_n393), .A2(new_n398), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT96), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT96), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n393), .A2(new_n603), .A3(new_n398), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n605), .B1(KEYINPUT36), .B2(new_n403), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n403), .A2(KEYINPUT36), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n602), .A2(new_n607), .A3(new_n604), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n606), .A2(new_n416), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(KEYINPUT97), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT97), .ZN(new_n611));
  NAND4_X1  g425(.A1(new_n606), .A2(new_n611), .A3(new_n416), .A4(new_n608), .ZN(new_n612));
  AND3_X1   g426(.A1(new_n414), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n613), .A2(new_n576), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n306), .A2(new_n421), .A3(new_n563), .A4(new_n614), .ZN(new_n615));
  XOR2_X1   g429(.A(KEYINPUT37), .B(G110), .Z(new_n616));
  XNOR2_X1  g430(.A(new_n615), .B(new_n616), .ZN(G12));
  AOI21_X1  g431(.A(new_n613), .B1(new_n357), .B2(new_n366), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n572), .A2(new_n562), .A3(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(G900), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n479), .B1(new_n480), .B2(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n596), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  INV_X1    g439(.A(new_n562), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT100), .B(KEYINPUT39), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n622), .B(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n626), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n630), .A2(KEYINPUT101), .ZN(new_n631));
  INV_X1    g445(.A(KEYINPUT40), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(KEYINPUT101), .ZN(new_n633));
  AND3_X1   g447(.A1(new_n631), .A2(new_n632), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n632), .B1(new_n631), .B2(new_n633), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n306), .B(KEYINPUT38), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n338), .B1(new_n344), .B2(new_n332), .ZN(new_n638));
  XOR2_X1   g452(.A(new_n638), .B(KEYINPUT98), .Z(new_n639));
  OAI21_X1  g453(.A(new_n364), .B1(new_n639), .B2(new_n350), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(G472), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n357), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT99), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n474), .A2(new_n517), .ZN(new_n644));
  AND4_X1   g458(.A1(new_n421), .A2(new_n643), .A3(new_n613), .A4(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n636), .A2(new_n637), .A3(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(G143), .ZN(G45));
  NOR2_X1   g461(.A1(new_n590), .A2(new_n622), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n620), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G146), .ZN(G48));
  NAND2_X1  g464(.A1(new_n546), .A2(new_n543), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n551), .B1(new_n651), .B2(new_n553), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(G902), .ZN(new_n653));
  NOR2_X1   g467(.A1(new_n653), .A2(new_n519), .ZN(new_n654));
  INV_X1    g468(.A(new_n552), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n561), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(new_n419), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n658), .B(new_n591), .C1(new_n567), .C2(new_n571), .ZN(new_n659));
  XNOR2_X1  g473(.A(KEYINPUT41), .B(G113), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G15));
  OAI211_X1 g475(.A(new_n658), .B(new_n597), .C1(new_n567), .C2(new_n571), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G116), .ZN(G18));
  INV_X1    g477(.A(new_n657), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n619), .A2(new_n518), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n664), .B(new_n665), .C1(new_n567), .C2(new_n571), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G119), .ZN(G21));
  NAND2_X1  g481(.A1(new_n577), .A2(new_n418), .ZN(new_n668));
  NOR3_X1   g482(.A1(new_n657), .A2(new_n482), .A3(new_n668), .ZN(new_n669));
  OAI211_X1 g483(.A(new_n644), .B(new_n669), .C1(new_n567), .C2(new_n571), .ZN(new_n670));
  XNOR2_X1  g484(.A(KEYINPUT102), .B(G122), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n670), .B(new_n671), .ZN(G24));
  AND2_X1   g486(.A1(new_n648), .A2(new_n614), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n664), .B(new_n673), .C1(new_n567), .C2(new_n571), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G125), .ZN(G27));
  INV_X1    g489(.A(new_n421), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n568), .A2(new_n569), .A3(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n560), .A2(new_n678), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n552), .A2(new_n557), .A3(KEYINPUT103), .A4(new_n559), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n679), .A2(new_n561), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n677), .A2(new_n420), .A3(new_n682), .A4(new_n648), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT104), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n304), .A2(new_n421), .A3(new_n305), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n681), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n687), .A2(KEYINPUT104), .A3(new_n420), .A4(new_n648), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT42), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n419), .B(KEYINPUT105), .Z(new_n691));
  NAND4_X1  g505(.A1(new_n691), .A2(KEYINPUT42), .A3(new_n648), .A4(new_n687), .ZN(new_n692));
  AND2_X1   g506(.A1(new_n690), .A2(new_n692), .ZN(new_n693));
  XOR2_X1   g507(.A(new_n693), .B(G131), .Z(G33));
  XNOR2_X1  g508(.A(new_n623), .B(KEYINPUT106), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n695), .A2(new_n677), .A3(new_n420), .A4(new_n682), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G134), .ZN(G36));
  NAND2_X1  g511(.A1(new_n474), .A2(KEYINPUT110), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n586), .B1(new_n474), .B2(KEYINPUT110), .ZN(new_n700));
  OAI21_X1  g514(.A(KEYINPUT43), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT109), .ZN(new_n702));
  AOI21_X1  g516(.A(KEYINPUT43), .B1(new_n585), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g517(.A(new_n703), .B(new_n474), .C1(new_n702), .C2(new_n585), .ZN(new_n704));
  AND2_X1   g518(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n414), .A2(new_n610), .A3(new_n612), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n576), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(new_n707), .B(KEYINPUT111), .Z(new_n708));
  NAND2_X1  g522(.A1(new_n705), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT44), .Z(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n686), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n651), .A2(new_n531), .ZN(new_n712));
  AOI22_X1  g526(.A1(new_n712), .A2(new_n534), .B1(new_n550), .B2(new_n553), .ZN(new_n713));
  OAI21_X1  g527(.A(G469), .B1(new_n713), .B2(KEYINPUT45), .ZN(new_n714));
  OR2_X1    g528(.A1(new_n714), .A2(KEYINPUT107), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(KEYINPUT45), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n714), .A2(KEYINPUT107), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n715), .A2(KEYINPUT108), .A3(new_n716), .A4(new_n717), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n558), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n552), .B1(new_n722), .B2(KEYINPUT46), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT46), .ZN(new_n724));
  AOI211_X1 g538(.A(new_n724), .B(new_n558), .C1(new_n720), .C2(new_n721), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n561), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n711), .A2(new_n628), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G137), .ZN(G39));
  INV_X1    g543(.A(KEYINPUT47), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n726), .A2(new_n730), .ZN(new_n731));
  OAI211_X1 g545(.A(KEYINPUT47), .B(new_n561), .C1(new_n723), .C2(new_n725), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NOR4_X1   g547(.A1(new_n590), .A2(new_n367), .A3(new_n418), .A4(new_n622), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n677), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G140), .ZN(G42));
  XOR2_X1   g550(.A(new_n656), .B(KEYINPUT49), .Z(new_n737));
  NOR2_X1   g551(.A1(new_n699), .A2(new_n700), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n738), .A2(new_n418), .A3(new_n421), .A4(new_n561), .ZN(new_n739));
  OR4_X1    g553(.A1(new_n637), .A2(new_n737), .A3(new_n643), .A4(new_n739), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n705), .A2(KEYINPUT116), .A3(new_n479), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n701), .A2(new_n704), .A3(new_n479), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT116), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n668), .B1(new_n741), .B2(new_n744), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n637), .A2(new_n421), .A3(new_n657), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT50), .ZN(new_n748));
  AND3_X1   g562(.A1(new_n747), .A2(KEYINPUT118), .A3(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n748), .B1(new_n747), .B2(KEYINPUT118), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n664), .A2(new_n677), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(KEYINPUT119), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n741), .A2(new_n744), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(new_n614), .ZN(new_n756));
  INV_X1    g570(.A(new_n418), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n643), .A2(new_n757), .A3(new_n478), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n474), .A2(new_n585), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n756), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n656), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n731), .B(new_n732), .C1(new_n561), .C2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n745), .A2(new_n677), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT117), .ZN(new_n770));
  AOI211_X1 g584(.A(new_n751), .B(new_n764), .C1(new_n769), .C2(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n766), .A2(KEYINPUT117), .A3(new_n768), .ZN(new_n772));
  AOI21_X1  g586(.A(KEYINPUT51), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT120), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n774), .B1(new_n764), .B2(new_n751), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n763), .B(KEYINPUT120), .C1(new_n750), .C2(new_n749), .ZN(new_n776));
  NAND4_X1  g590(.A1(new_n775), .A2(new_n776), .A3(new_n769), .A4(KEYINPUT51), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n755), .A2(new_n691), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(KEYINPUT48), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n778), .A2(KEYINPUT48), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n759), .A2(new_n589), .A3(new_n586), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n745), .A2(new_n573), .A3(new_n664), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n781), .A2(new_n475), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n777), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT114), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n619), .A2(new_n562), .ZN(new_n787));
  OAI221_X1 g601(.A(new_n787), .B1(new_n623), .B2(new_n648), .C1(new_n567), .C2(new_n571), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n706), .A2(new_n622), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT113), .ZN(new_n790));
  AND3_X1   g604(.A1(new_n682), .A2(new_n790), .A3(new_n642), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n644), .C1(new_n567), .C2(new_n571), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n674), .A3(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n793), .A2(KEYINPUT52), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n662), .A2(new_n666), .A3(new_n670), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n482), .B1(new_n590), .B2(new_n596), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n306), .A2(new_n421), .A3(new_n579), .A4(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n564), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n659), .A2(new_n798), .A3(new_n615), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n795), .A2(new_n799), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n673), .A2(new_n677), .A3(new_n682), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n589), .A2(new_n516), .A3(new_n622), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n618), .A2(new_n561), .A3(new_n802), .A4(new_n560), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g618(.A(KEYINPUT112), .B1(new_n804), .B2(new_n677), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  NOR3_X1   g620(.A1(new_n686), .A2(new_n803), .A3(new_n806), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n696), .B(new_n801), .C1(new_n805), .C2(new_n807), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n808), .B1(new_n690), .B2(new_n692), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT52), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n788), .A2(new_n792), .A3(new_n810), .A4(new_n674), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n794), .A2(new_n800), .A3(new_n809), .A4(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT53), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n786), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n794), .A2(new_n811), .ZN(new_n815));
  AND2_X1   g629(.A1(new_n800), .A2(new_n809), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(KEYINPUT53), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n817), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n815), .A2(new_n816), .A3(new_n786), .A4(KEYINPUT53), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(KEYINPUT54), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n812), .A2(new_n813), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n817), .A2(new_n821), .A3(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n817), .A2(KEYINPUT115), .A3(new_n822), .A4(new_n821), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n820), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n773), .A2(new_n785), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(G952), .A2(G953), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n740), .B1(new_n828), .B2(new_n829), .ZN(G75));
  AOI21_X1  g644(.A(new_n364), .B1(new_n817), .B2(new_n822), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n831), .A2(G210), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT56), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n253), .A2(new_n261), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n285), .ZN(new_n835));
  XNOR2_X1  g649(.A(new_n835), .B(KEYINPUT55), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n832), .A2(new_n833), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n836), .B1(new_n832), .B2(new_n833), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n399), .A2(G952), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(G51));
  XNOR2_X1  g654(.A(new_n558), .B(KEYINPUT57), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n817), .A2(new_n821), .A3(new_n822), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n821), .B1(new_n817), .B2(new_n822), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n841), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n652), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(new_n845), .B2(new_n844), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n831), .A2(new_n720), .A3(new_n721), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n839), .B1(new_n847), .B2(new_n848), .ZN(G54));
  NAND3_X1  g663(.A1(new_n831), .A2(KEYINPUT58), .A3(G475), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n462), .A2(new_n463), .ZN(new_n851));
  OAI21_X1  g665(.A(new_n851), .B1(new_n449), .B2(new_n452), .ZN(new_n852));
  INV_X1    g666(.A(new_n434), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n852), .A2(new_n853), .B1(new_n470), .B2(new_n436), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n850), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n850), .A2(new_n854), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n855), .A2(new_n856), .A3(new_n839), .ZN(G60));
  XNOR2_X1  g671(.A(new_n583), .B(KEYINPUT59), .ZN(new_n858));
  INV_X1    g672(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n827), .A2(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n580), .A2(new_n581), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n860), .A2(KEYINPUT123), .A3(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n858), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n815), .B2(new_n816), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n812), .A2(new_n813), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT54), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n867), .B2(new_n823), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT122), .B1(new_n868), .B2(new_n839), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n863), .B1(new_n842), .B2(new_n843), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n871));
  INV_X1    g685(.A(new_n839), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n869), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT123), .B1(new_n860), .B2(new_n861), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(G63));
  NAND2_X1  g691(.A1(G217), .A2(G902), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT60), .Z(new_n879));
  OAI21_X1  g693(.A(new_n879), .B1(new_n865), .B2(new_n866), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n839), .B1(new_n880), .B2(new_n407), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n606), .A2(new_n608), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(new_n880), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n883), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g698(.A(G953), .B1(new_n481), .B2(new_n282), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n800), .B2(G953), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n834), .B1(G898), .B2(new_n399), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n886), .B(new_n887), .ZN(G69));
  NAND2_X1  g702(.A1(new_n328), .A2(new_n329), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n456), .A2(new_n460), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT124), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n889), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n590), .A2(new_n596), .ZN(new_n893));
  XOR2_X1   g707(.A(new_n893), .B(KEYINPUT125), .Z(new_n894));
  NOR2_X1   g708(.A1(new_n894), .A2(new_n419), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n895), .A2(new_n633), .A3(new_n631), .A4(new_n677), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n728), .A2(new_n896), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(new_n735), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n646), .A2(new_n674), .A3(new_n788), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT62), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  AOI211_X1 g715(.A(G953), .B(new_n892), .C1(new_n898), .C2(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n892), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n573), .A2(new_n644), .A3(new_n691), .ZN(new_n904));
  OAI211_X1 g718(.A(new_n727), .B(new_n628), .C1(new_n711), .C2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n788), .A2(new_n674), .A3(new_n696), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n693), .A2(new_n906), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n735), .A2(new_n905), .A3(new_n399), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(G900), .A2(G953), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n903), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AOI21_X1  g724(.A(new_n399), .B1(G227), .B2(G900), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n902), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n908), .A2(new_n909), .ZN(new_n913));
  NAND2_X1  g727(.A1(G227), .A2(G900), .ZN(new_n914));
  AND4_X1   g728(.A1(G953), .A2(new_n913), .A3(new_n914), .A4(new_n892), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G72));
  NAND2_X1  g730(.A1(G472), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT63), .Z(new_n918));
  NOR2_X1   g732(.A1(new_n350), .A2(KEYINPUT127), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n362), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n818), .A2(new_n819), .A3(new_n918), .A4(new_n920), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n735), .A2(new_n905), .A3(new_n800), .A4(new_n907), .ZN(new_n922));
  AND2_X1   g736(.A1(new_n922), .A2(new_n918), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n361), .A2(new_n341), .ZN(new_n924));
  OAI211_X1 g738(.A(new_n872), .B(new_n921), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n901), .A2(new_n735), .A3(new_n800), .A4(new_n897), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n918), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n361), .A2(new_n341), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n929), .A2(KEYINPUT126), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n927), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n925), .B1(new_n930), .B2(new_n932), .ZN(G57));
endmodule


