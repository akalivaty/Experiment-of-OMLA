

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586;

  NOR2_X1 U326 ( .A1(n549), .A2(n296), .ZN(n571) );
  XNOR2_X2 U327 ( .A(n554), .B(KEYINPUT121), .ZN(n567) );
  BUF_X1 U328 ( .A(n547), .Z(n294) );
  XNOR2_X1 U329 ( .A(n522), .B(KEYINPUT48), .ZN(n547) );
  NOR2_X1 U330 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U331 ( .A(n331), .B(n330), .ZN(n577) );
  AND2_X1 U332 ( .A1(n561), .A2(n555), .ZN(n512) );
  XOR2_X1 U333 ( .A(n326), .B(n325), .Z(n295) );
  XOR2_X1 U334 ( .A(KEYINPUT54), .B(n548), .Z(n296) );
  XOR2_X1 U335 ( .A(G99GAT), .B(G85GAT), .Z(n334) );
  XNOR2_X1 U336 ( .A(G92GAT), .B(G64GAT), .ZN(n315) );
  XOR2_X1 U337 ( .A(G57GAT), .B(KEYINPUT13), .Z(n354) );
  XOR2_X1 U338 ( .A(n314), .B(n313), .Z(n555) );
  XOR2_X1 U339 ( .A(KEYINPUT67), .B(KEYINPUT30), .Z(n298) );
  XNOR2_X1 U340 ( .A(G15GAT), .B(G1GAT), .ZN(n297) );
  XNOR2_X1 U341 ( .A(n298), .B(n297), .ZN(n314) );
  XOR2_X1 U342 ( .A(G113GAT), .B(G197GAT), .Z(n300) );
  XNOR2_X1 U343 ( .A(G141GAT), .B(G22GAT), .ZN(n299) );
  XNOR2_X1 U344 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U345 ( .A(n301), .B(G50GAT), .Z(n303) );
  XOR2_X1 U346 ( .A(G169GAT), .B(G8GAT), .Z(n418) );
  XNOR2_X1 U347 ( .A(n418), .B(G36GAT), .ZN(n302) );
  XNOR2_X1 U348 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U349 ( .A(KEYINPUT29), .B(KEYINPUT70), .Z(n305) );
  NAND2_X1 U350 ( .A1(G229GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U352 ( .A(n307), .B(n306), .Z(n312) );
  XOR2_X1 U353 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n309) );
  XNOR2_X1 U354 ( .A(G43GAT), .B(G29GAT), .ZN(n308) );
  XNOR2_X1 U355 ( .A(n309), .B(n308), .ZN(n310) );
  XOR2_X1 U356 ( .A(KEYINPUT69), .B(n310), .Z(n345) );
  XNOR2_X1 U357 ( .A(n345), .B(KEYINPUT68), .ZN(n311) );
  XNOR2_X1 U358 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G71GAT), .Z(n393) );
  INV_X1 U360 ( .A(n315), .ZN(n317) );
  XNOR2_X1 U361 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n316) );
  XNOR2_X1 U362 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U363 ( .A(G176GAT), .B(n318), .Z(n410) );
  XNOR2_X1 U364 ( .A(n393), .B(n410), .ZN(n320) );
  INV_X1 U365 ( .A(KEYINPUT33), .ZN(n319) );
  XNOR2_X1 U366 ( .A(n320), .B(n319), .ZN(n327) );
  XOR2_X1 U367 ( .A(n354), .B(n334), .Z(n322) );
  NAND2_X1 U368 ( .A1(G230GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U369 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U370 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n324) );
  XNOR2_X1 U371 ( .A(KEYINPUT74), .B(KEYINPUT32), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U373 ( .A(n327), .B(n295), .ZN(n331) );
  XOR2_X1 U374 ( .A(G78GAT), .B(G148GAT), .Z(n329) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(KEYINPUT73), .ZN(n328) );
  XNOR2_X1 U376 ( .A(n329), .B(n328), .ZN(n423) );
  XNOR2_X1 U377 ( .A(n423), .B(KEYINPUT72), .ZN(n330) );
  NAND2_X1 U378 ( .A1(n555), .A2(n577), .ZN(n470) );
  XOR2_X1 U379 ( .A(KEYINPUT10), .B(KEYINPUT76), .Z(n333) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(KEYINPUT9), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n344) );
  XOR2_X1 U382 ( .A(KEYINPUT66), .B(n334), .Z(n336) );
  XOR2_X1 U383 ( .A(G36GAT), .B(G190GAT), .Z(n414) );
  XNOR2_X1 U384 ( .A(G218GAT), .B(n414), .ZN(n335) );
  XNOR2_X1 U385 ( .A(n336), .B(n335), .ZN(n340) );
  XOR2_X1 U386 ( .A(KEYINPUT11), .B(G92GAT), .Z(n338) );
  NAND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U388 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U389 ( .A(n340), .B(n339), .Z(n342) );
  XOR2_X1 U390 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U391 ( .A(G134GAT), .B(KEYINPUT77), .Z(n374) );
  XNOR2_X1 U392 ( .A(n428), .B(n374), .ZN(n341) );
  XNOR2_X1 U393 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U394 ( .A(n344), .B(n343), .ZN(n347) );
  INV_X1 U395 ( .A(n345), .ZN(n346) );
  XOR2_X1 U396 ( .A(n347), .B(n346), .Z(n566) );
  XOR2_X1 U397 ( .A(G71GAT), .B(G183GAT), .Z(n349) );
  XNOR2_X1 U398 ( .A(G1GAT), .B(G8GAT), .ZN(n348) );
  XNOR2_X1 U399 ( .A(n349), .B(n348), .ZN(n353) );
  XOR2_X1 U400 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n351) );
  XNOR2_X1 U401 ( .A(G64GAT), .B(KEYINPUT12), .ZN(n350) );
  XNOR2_X1 U402 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U403 ( .A(n353), .B(n352), .ZN(n364) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G155GAT), .Z(n427) );
  XOR2_X1 U405 ( .A(n354), .B(n427), .Z(n356) );
  XNOR2_X1 U406 ( .A(G211GAT), .B(G78GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U408 ( .A(KEYINPUT78), .B(KEYINPUT14), .Z(n358) );
  NAND2_X1 U409 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U410 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U411 ( .A(n360), .B(n359), .Z(n362) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G127GAT), .Z(n396) );
  XNOR2_X1 U413 ( .A(n396), .B(KEYINPUT15), .ZN(n361) );
  XNOR2_X1 U414 ( .A(n362), .B(n361), .ZN(n363) );
  XNOR2_X1 U415 ( .A(n364), .B(n363), .ZN(n564) );
  INV_X1 U416 ( .A(n564), .ZN(n581) );
  NOR2_X1 U417 ( .A1(n566), .A2(n581), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n365), .B(KEYINPUT16), .ZN(n454) );
  XOR2_X1 U419 ( .A(G57GAT), .B(KEYINPUT1), .Z(n367) );
  XNOR2_X1 U420 ( .A(G1GAT), .B(G120GAT), .ZN(n366) );
  XNOR2_X1 U421 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U422 ( .A(G85GAT), .B(G155GAT), .Z(n369) );
  XNOR2_X1 U423 ( .A(G127GAT), .B(G148GAT), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U425 ( .A(n371), .B(n370), .ZN(n387) );
  XOR2_X1 U426 ( .A(KEYINPUT5), .B(KEYINPUT92), .Z(n373) );
  XNOR2_X1 U427 ( .A(KEYINPUT4), .B(KEYINPUT91), .ZN(n372) );
  XNOR2_X1 U428 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U429 ( .A(n374), .B(G162GAT), .Z(n376) );
  XOR2_X1 U430 ( .A(G113GAT), .B(KEYINPUT0), .Z(n405) );
  XNOR2_X1 U431 ( .A(G29GAT), .B(n405), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U433 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U434 ( .A1(G225GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U435 ( .A(n380), .B(n379), .ZN(n382) );
  INV_X1 U436 ( .A(KEYINPUT90), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n385) );
  XNOR2_X1 U438 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n383), .B(KEYINPUT2), .ZN(n436) );
  XNOR2_X1 U440 ( .A(n436), .B(KEYINPUT6), .ZN(n384) );
  XNOR2_X1 U441 ( .A(n385), .B(n384), .ZN(n386) );
  XNOR2_X1 U442 ( .A(n387), .B(n386), .ZN(n549) );
  XOR2_X1 U443 ( .A(KEYINPUT20), .B(KEYINPUT85), .Z(n389) );
  XNOR2_X1 U444 ( .A(G169GAT), .B(KEYINPUT65), .ZN(n388) );
  XNOR2_X1 U445 ( .A(n389), .B(n388), .ZN(n409) );
  XOR2_X1 U446 ( .A(KEYINPUT84), .B(G176GAT), .Z(n391) );
  XNOR2_X1 U447 ( .A(G134GAT), .B(G190GAT), .ZN(n390) );
  XNOR2_X1 U448 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U449 ( .A(n392), .B(G99GAT), .Z(n395) );
  XNOR2_X1 U450 ( .A(G43GAT), .B(n393), .ZN(n394) );
  XNOR2_X1 U451 ( .A(n395), .B(n394), .ZN(n400) );
  XOR2_X1 U452 ( .A(n396), .B(KEYINPUT81), .Z(n398) );
  NAND2_X1 U453 ( .A1(G227GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U454 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U455 ( .A(n400), .B(n399), .Z(n407) );
  XNOR2_X1 U456 ( .A(KEYINPUT82), .B(KEYINPUT18), .ZN(n401) );
  XNOR2_X1 U457 ( .A(n401), .B(G183GAT), .ZN(n402) );
  XOR2_X1 U458 ( .A(n402), .B(KEYINPUT83), .Z(n404) );
  XNOR2_X1 U459 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n403) );
  XNOR2_X1 U460 ( .A(n404), .B(n403), .ZN(n411) );
  XNOR2_X1 U461 ( .A(n411), .B(n405), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U463 ( .A(n409), .B(n408), .ZN(n552) );
  XNOR2_X1 U464 ( .A(n411), .B(n410), .ZN(n422) );
  XOR2_X1 U465 ( .A(G211GAT), .B(KEYINPUT21), .Z(n413) );
  XNOR2_X1 U466 ( .A(G197GAT), .B(G218GAT), .ZN(n412) );
  XNOR2_X1 U467 ( .A(n413), .B(n412), .ZN(n424) );
  XOR2_X1 U468 ( .A(n414), .B(n424), .Z(n416) );
  NAND2_X1 U469 ( .A1(G226GAT), .A2(G233GAT), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n417) );
  XOR2_X1 U471 ( .A(n417), .B(KEYINPUT94), .Z(n420) );
  XNOR2_X1 U472 ( .A(n418), .B(KEYINPUT93), .ZN(n419) );
  XNOR2_X1 U473 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U474 ( .A(n422), .B(n421), .ZN(n546) );
  INV_X1 U475 ( .A(n546), .ZN(n502) );
  NAND2_X1 U476 ( .A1(n552), .A2(n502), .ZN(n441) );
  XNOR2_X1 U477 ( .A(n424), .B(n423), .ZN(n440) );
  XOR2_X1 U478 ( .A(KEYINPUT23), .B(KEYINPUT86), .Z(n426) );
  XNOR2_X1 U479 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n426), .B(n425), .ZN(n432) );
  XOR2_X1 U481 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n430) );
  XNOR2_X1 U482 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U483 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U484 ( .A(n432), .B(n431), .Z(n434) );
  NAND2_X1 U485 ( .A1(G228GAT), .A2(G233GAT), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U487 ( .A(n435), .B(KEYINPUT24), .Z(n438) );
  XNOR2_X1 U488 ( .A(n436), .B(KEYINPUT22), .ZN(n437) );
  XNOR2_X1 U489 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n550) );
  NAND2_X1 U491 ( .A1(n441), .A2(n550), .ZN(n442) );
  XNOR2_X1 U492 ( .A(n442), .B(KEYINPUT97), .ZN(n443) );
  XOR2_X1 U493 ( .A(KEYINPUT25), .B(n443), .Z(n446) );
  XNOR2_X1 U494 ( .A(n502), .B(KEYINPUT27), .ZN(n448) );
  NOR2_X1 U495 ( .A1(n550), .A2(n552), .ZN(n444) );
  XNOR2_X1 U496 ( .A(KEYINPUT26), .B(n444), .ZN(n570) );
  AND2_X1 U497 ( .A1(n448), .A2(n570), .ZN(n445) );
  NOR2_X1 U498 ( .A1(n446), .A2(n445), .ZN(n447) );
  NOR2_X1 U499 ( .A1(n549), .A2(n447), .ZN(n452) );
  XOR2_X2 U500 ( .A(n550), .B(KEYINPUT28), .Z(n507) );
  NAND2_X1 U501 ( .A1(n549), .A2(n448), .ZN(n536) );
  NOR2_X1 U502 ( .A1(n507), .A2(n536), .ZN(n523) );
  XNOR2_X1 U503 ( .A(KEYINPUT95), .B(n523), .ZN(n449) );
  NOR2_X1 U504 ( .A1(n552), .A2(n449), .ZN(n450) );
  XNOR2_X1 U505 ( .A(n450), .B(KEYINPUT96), .ZN(n451) );
  NOR2_X1 U506 ( .A1(n452), .A2(n451), .ZN(n466) );
  INV_X1 U507 ( .A(n466), .ZN(n453) );
  NAND2_X1 U508 ( .A1(n454), .A2(n453), .ZN(n486) );
  NOR2_X1 U509 ( .A1(n470), .A2(n486), .ZN(n464) );
  NAND2_X1 U510 ( .A1(n464), .A2(n549), .ZN(n458) );
  XOR2_X1 U511 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n456) );
  XNOR2_X1 U512 ( .A(G1GAT), .B(KEYINPUT99), .ZN(n455) );
  XNOR2_X1 U513 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U514 ( .A(n458), .B(n457), .ZN(G1324GAT) );
  NAND2_X1 U515 ( .A1(n502), .A2(n464), .ZN(n459) );
  XNOR2_X1 U516 ( .A(n459), .B(KEYINPUT100), .ZN(n460) );
  XNOR2_X1 U517 ( .A(G8GAT), .B(n460), .ZN(G1325GAT) );
  XOR2_X1 U518 ( .A(KEYINPUT101), .B(KEYINPUT35), .Z(n462) );
  NAND2_X1 U519 ( .A1(n464), .A2(n552), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n462), .B(n461), .ZN(n463) );
  XOR2_X1 U521 ( .A(G15GAT), .B(n463), .Z(G1326GAT) );
  NAND2_X1 U522 ( .A1(n464), .A2(n507), .ZN(n465) );
  XNOR2_X1 U523 ( .A(n465), .B(G22GAT), .ZN(G1327GAT) );
  INV_X1 U524 ( .A(n566), .ZN(n514) );
  XNOR2_X1 U525 ( .A(KEYINPUT36), .B(n514), .ZN(n584) );
  NOR2_X1 U526 ( .A1(n584), .A2(n466), .ZN(n467) );
  NAND2_X1 U527 ( .A1(n581), .A2(n467), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(KEYINPUT37), .ZN(n469) );
  XNOR2_X1 U529 ( .A(KEYINPUT103), .B(n469), .ZN(n497) );
  NOR2_X1 U530 ( .A1(n497), .A2(n470), .ZN(n472) );
  XNOR2_X1 U531 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n471) );
  XNOR2_X1 U532 ( .A(n472), .B(n471), .ZN(n483) );
  NAND2_X1 U533 ( .A1(n483), .A2(n549), .ZN(n475) );
  XOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT102), .Z(n473) );
  XNOR2_X1 U535 ( .A(KEYINPUT39), .B(n473), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(G1328GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n477) );
  NAND2_X1 U538 ( .A1(n483), .A2(n502), .ZN(n476) );
  XNOR2_X1 U539 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U540 ( .A(G36GAT), .B(n478), .ZN(G1329GAT) );
  XNOR2_X1 U541 ( .A(G43GAT), .B(KEYINPUT108), .ZN(n482) );
  XOR2_X1 U542 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n480) );
  NAND2_X1 U543 ( .A1(n483), .A2(n552), .ZN(n479) );
  XNOR2_X1 U544 ( .A(n480), .B(n479), .ZN(n481) );
  XNOR2_X1 U545 ( .A(n482), .B(n481), .ZN(G1330GAT) );
  NAND2_X1 U546 ( .A1(n483), .A2(n507), .ZN(n484) );
  XNOR2_X1 U547 ( .A(n484), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT42), .B(KEYINPUT109), .Z(n488) );
  XNOR2_X1 U549 ( .A(n577), .B(KEYINPUT64), .ZN(n485) );
  XNOR2_X1 U550 ( .A(KEYINPUT41), .B(n485), .ZN(n561) );
  INV_X1 U551 ( .A(n555), .ZN(n572) );
  NAND2_X1 U552 ( .A1(n561), .A2(n572), .ZN(n498) );
  NOR2_X1 U553 ( .A1(n498), .A2(n486), .ZN(n494) );
  NAND2_X1 U554 ( .A1(n494), .A2(n549), .ZN(n487) );
  XNOR2_X1 U555 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U556 ( .A(G57GAT), .B(n489), .ZN(G1332GAT) );
  NAND2_X1 U557 ( .A1(n502), .A2(n494), .ZN(n490) );
  XNOR2_X1 U558 ( .A(n490), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U559 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n492) );
  NAND2_X1 U560 ( .A1(n494), .A2(n552), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U562 ( .A(G71GAT), .B(n493), .ZN(G1334GAT) );
  XOR2_X1 U563 ( .A(G78GAT), .B(KEYINPUT43), .Z(n496) );
  NAND2_X1 U564 ( .A1(n494), .A2(n507), .ZN(n495) );
  XNOR2_X1 U565 ( .A(n496), .B(n495), .ZN(G1335GAT) );
  NOR2_X1 U566 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U567 ( .A(n499), .B(KEYINPUT112), .ZN(n506) );
  NAND2_X1 U568 ( .A1(n549), .A2(n506), .ZN(n501) );
  XOR2_X1 U569 ( .A(G85GAT), .B(KEYINPUT113), .Z(n500) );
  XNOR2_X1 U570 ( .A(n501), .B(n500), .ZN(G1336GAT) );
  NAND2_X1 U571 ( .A1(n506), .A2(n502), .ZN(n503) );
  XNOR2_X1 U572 ( .A(n503), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U573 ( .A1(n506), .A2(n552), .ZN(n504) );
  XNOR2_X1 U574 ( .A(n504), .B(KEYINPUT114), .ZN(n505) );
  XNOR2_X1 U575 ( .A(G99GAT), .B(n505), .ZN(G1338GAT) );
  XOR2_X1 U576 ( .A(KEYINPUT44), .B(KEYINPUT115), .Z(n509) );
  NAND2_X1 U577 ( .A1(n507), .A2(n506), .ZN(n508) );
  XNOR2_X1 U578 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U579 ( .A(G106GAT), .B(n510), .ZN(G1339GAT) );
  XOR2_X1 U580 ( .A(G113GAT), .B(KEYINPUT117), .Z(n526) );
  XNOR2_X1 U581 ( .A(KEYINPUT46), .B(KEYINPUT116), .ZN(n511) );
  XNOR2_X1 U582 ( .A(n512), .B(n511), .ZN(n513) );
  NOR2_X1 U583 ( .A1(n564), .A2(n513), .ZN(n515) );
  NAND2_X1 U584 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U585 ( .A(n516), .B(KEYINPUT47), .ZN(n521) );
  NOR2_X1 U586 ( .A1(n584), .A2(n581), .ZN(n517) );
  XNOR2_X1 U587 ( .A(KEYINPUT45), .B(n517), .ZN(n518) );
  NAND2_X1 U588 ( .A1(n518), .A2(n577), .ZN(n519) );
  NOR2_X1 U589 ( .A1(n519), .A2(n555), .ZN(n520) );
  NAND2_X1 U590 ( .A1(n523), .A2(n552), .ZN(n524) );
  NOR2_X1 U591 ( .A1(n294), .A2(n524), .ZN(n532) );
  NAND2_X1 U592 ( .A1(n532), .A2(n555), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(G120GAT), .B(KEYINPUT49), .Z(n528) );
  NAND2_X1 U595 ( .A1(n532), .A2(n561), .ZN(n527) );
  XNOR2_X1 U596 ( .A(n528), .B(n527), .ZN(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT118), .B(KEYINPUT50), .Z(n530) );
  NAND2_X1 U598 ( .A1(n532), .A2(n564), .ZN(n529) );
  XNOR2_X1 U599 ( .A(n530), .B(n529), .ZN(n531) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n531), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT119), .B(KEYINPUT51), .Z(n534) );
  NAND2_X1 U602 ( .A1(n532), .A2(n566), .ZN(n533) );
  XNOR2_X1 U603 ( .A(n534), .B(n533), .ZN(n535) );
  XOR2_X1 U604 ( .A(G134GAT), .B(n535), .Z(G1343GAT) );
  NOR2_X1 U605 ( .A1(n294), .A2(n536), .ZN(n537) );
  NAND2_X1 U606 ( .A1(n570), .A2(n537), .ZN(n538) );
  XOR2_X1 U607 ( .A(KEYINPUT120), .B(n538), .Z(n544) );
  NAND2_X1 U608 ( .A1(n544), .A2(n555), .ZN(n539) );
  XNOR2_X1 U609 ( .A(n539), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n541) );
  NAND2_X1 U611 ( .A1(n561), .A2(n544), .ZN(n540) );
  XNOR2_X1 U612 ( .A(n541), .B(n540), .ZN(n542) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n542), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n544), .A2(n564), .ZN(n543) );
  XNOR2_X1 U615 ( .A(n543), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n544), .A2(n566), .ZN(n545) );
  XNOR2_X1 U617 ( .A(n545), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(KEYINPUT122), .ZN(n557) );
  NOR2_X1 U619 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U620 ( .A1(n550), .A2(n571), .ZN(n551) );
  XNOR2_X1 U621 ( .A(n551), .B(KEYINPUT55), .ZN(n553) );
  NAND2_X1 U622 ( .A1(n553), .A2(n552), .ZN(n554) );
  NAND2_X1 U623 ( .A1(n555), .A2(n567), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT57), .B(KEYINPUT124), .Z(n559) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(n560) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(n560), .Z(n563) );
  NAND2_X1 U629 ( .A1(n567), .A2(n561), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n563), .B(n562), .ZN(G1349GAT) );
  NAND2_X1 U631 ( .A1(n567), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U633 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n569) );
  NAND2_X1 U634 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(G1351GAT) );
  NAND2_X1 U636 ( .A1(n571), .A2(n570), .ZN(n583) );
  NOR2_X1 U637 ( .A1(n572), .A2(n583), .ZN(n574) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n573) );
  XNOR2_X1 U639 ( .A(n574), .B(n573), .ZN(n576) );
  XOR2_X1 U640 ( .A(KEYINPUT125), .B(KEYINPUT59), .Z(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n583), .ZN(n579) );
  XNOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U646 ( .A1(n581), .A2(n583), .ZN(n582) );
  XOR2_X1 U647 ( .A(G211GAT), .B(n582), .Z(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

