//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:51 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n553,
    new_n554, new_n555, new_n558, new_n559, new_n561, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n587, new_n590,
    new_n592, new_n593, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n609, new_n610, new_n611, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G2105), .ZN(new_n458));
  NAND3_X1  g033(.A1(new_n458), .A2(G101), .A3(G2104), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(new_n458), .ZN(new_n465));
  INV_X1    g040(.A(G137), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n459), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n464), .A2(G125), .ZN(new_n468));
  NAND2_X1  g043(.A1(G113), .A2(G2104), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n458), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n467), .A2(new_n470), .ZN(G160));
  AOI21_X1  g046(.A(new_n458), .B1(new_n462), .B2(new_n463), .ZN(new_n472));
  AOI21_X1  g047(.A(G2105), .B1(new_n462), .B2(new_n463), .ZN(new_n473));
  AOI22_X1  g048(.A1(G124), .A2(new_n472), .B1(new_n473), .B2(G136), .ZN(new_n474));
  OR2_X1    g049(.A1(G100), .A2(G2105), .ZN(new_n475));
  OAI211_X1 g050(.A(new_n475), .B(G2104), .C1(G112), .C2(new_n458), .ZN(new_n476));
  AND2_X1   g051(.A1(new_n476), .A2(KEYINPUT64), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n476), .A2(KEYINPUT64), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  XOR2_X1   g054(.A(new_n479), .B(KEYINPUT65), .Z(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G162));
  AND2_X1   g056(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n482));
  NOR2_X1   g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  OAI211_X1 g058(.A(G126), .B(G2105), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(G114), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(new_n482), .B2(new_n483), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n464), .A2(new_n493), .A3(new_n490), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n488), .B1(new_n492), .B2(new_n494), .ZN(G164));
  NAND2_X1  g070(.A1(KEYINPUT66), .A2(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND3_X1  g073(.A1(KEYINPUT66), .A2(KEYINPUT5), .A3(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XOR2_X1   g080(.A(KEYINPUT67), .B(G88), .Z(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n503), .A2(new_n509), .ZN(G166));
  INV_X1    g085(.A(KEYINPUT71), .ZN(new_n511));
  INV_X1    g086(.A(new_n505), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(G89), .ZN(new_n513));
  XNOR2_X1  g088(.A(KEYINPUT69), .B(KEYINPUT7), .ZN(new_n514));
  XNOR2_X1  g089(.A(new_n514), .B(KEYINPUT70), .ZN(new_n515));
  NAND3_X1  g090(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT70), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n514), .B(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n516), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI211_X1 g096(.A(new_n511), .B(new_n513), .C1(new_n517), .C2(new_n521), .ZN(new_n522));
  AND3_X1   g097(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n507), .B(KEYINPUT68), .ZN(new_n524));
  AOI21_X1  g099(.A(new_n523), .B1(new_n524), .B2(G51), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n515), .B(new_n516), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n511), .B1(new_n527), .B2(new_n513), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n526), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n530), .A2(new_n502), .B1(new_n531), .B2(new_n505), .ZN(new_n532));
  AOI21_X1  g107(.A(new_n532), .B1(G52), .B2(new_n524), .ZN(G171));
  AOI22_X1  g108(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G81), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n534), .A2(new_n502), .B1(new_n535), .B2(new_n505), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n536), .B1(G43), .B2(new_n524), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G860), .ZN(G153));
  NAND4_X1  g113(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g114(.A1(G1), .A2(G3), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT8), .ZN(new_n541));
  NAND4_X1  g116(.A1(G319), .A2(G483), .A3(G661), .A4(new_n541), .ZN(G188));
  AND2_X1   g117(.A1(new_n504), .A2(G543), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G53), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT9), .ZN(new_n545));
  NAND2_X1  g120(.A1(G78), .A2(G543), .ZN(new_n546));
  INV_X1    g121(.A(new_n500), .ZN(new_n547));
  INV_X1    g122(.A(G65), .ZN(new_n548));
  OAI21_X1  g123(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  AOI22_X1  g124(.A1(new_n549), .A2(G651), .B1(new_n512), .B2(G91), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n545), .A2(new_n550), .ZN(G299));
  INV_X1    g126(.A(G171), .ZN(G301));
  AND2_X1   g127(.A1(new_n522), .A2(new_n525), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n527), .A2(new_n513), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(KEYINPUT71), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n553), .A2(new_n555), .ZN(G286));
  INV_X1    g131(.A(G166), .ZN(G303));
  AOI22_X1  g132(.A1(new_n512), .A2(G87), .B1(new_n543), .B2(G49), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n558), .A2(new_n559), .ZN(G288));
  NAND2_X1  g135(.A1(G73), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G61), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n547), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n563), .A2(G651), .B1(new_n512), .B2(G86), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n565));
  INV_X1    g140(.A(KEYINPUT72), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n565), .B(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n564), .A2(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n524), .A2(G47), .B1(G85), .B2(new_n512), .ZN(new_n569));
  INV_X1    g144(.A(KEYINPUT73), .ZN(new_n570));
  AOI22_X1  g145(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n571), .B2(new_n502), .ZN(new_n572));
  OR3_X1    g147(.A1(new_n571), .A2(new_n570), .A3(new_n502), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n569), .A2(new_n572), .A3(new_n573), .ZN(G290));
  INV_X1    g149(.A(G868), .ZN(new_n575));
  NOR2_X1   g150(.A1(G301), .A2(new_n575), .ZN(new_n576));
  AND3_X1   g151(.A1(new_n500), .A2(G92), .A3(new_n504), .ZN(new_n577));
  XNOR2_X1  g152(.A(new_n577), .B(KEYINPUT10), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n524), .A2(G54), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n500), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n580));
  OAI211_X1 g155(.A(new_n578), .B(new_n579), .C1(new_n502), .C2(new_n580), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(KEYINPUT74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(KEYINPUT74), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n576), .B1(new_n584), .B2(new_n575), .ZN(G284));
  XNOR2_X1  g160(.A(G284), .B(KEYINPUT75), .ZN(G321));
  NAND2_X1  g161(.A1(G299), .A2(new_n575), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n587), .B1(G168), .B2(new_n575), .ZN(G297));
  OAI21_X1  g163(.A(new_n587), .B1(G168), .B2(new_n575), .ZN(G280));
  INV_X1    g164(.A(G559), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n584), .B1(new_n590), .B2(G860), .ZN(G148));
  NAND2_X1  g166(.A1(new_n584), .A2(new_n590), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n592), .A2(G868), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n593), .B1(G868), .B2(new_n537), .ZN(G323));
  XNOR2_X1  g169(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g170(.A(KEYINPUT76), .B(KEYINPUT12), .ZN(new_n596));
  NOR3_X1   g171(.A1(new_n460), .A2(new_n461), .A3(G2105), .ZN(new_n597));
  XNOR2_X1  g172(.A(new_n596), .B(new_n597), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n598), .B(KEYINPUT13), .ZN(new_n599));
  OR2_X1    g174(.A1(new_n599), .A2(G2100), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n473), .A2(G135), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n472), .A2(G123), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n458), .A2(G111), .ZN(new_n603));
  OAI21_X1  g178(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n604));
  OAI211_X1 g179(.A(new_n601), .B(new_n602), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(G2096), .Z(new_n606));
  NAND2_X1  g181(.A1(new_n599), .A2(G2100), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n600), .A2(new_n606), .A3(new_n607), .ZN(G156));
  INV_X1    g183(.A(KEYINPUT14), .ZN(new_n609));
  XNOR2_X1  g184(.A(G2427), .B(G2438), .ZN(new_n610));
  XNOR2_X1  g185(.A(new_n610), .B(G2430), .ZN(new_n611));
  XNOR2_X1  g186(.A(KEYINPUT15), .B(G2435), .ZN(new_n612));
  AOI21_X1  g187(.A(new_n609), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n613), .B1(new_n612), .B2(new_n611), .ZN(new_n614));
  XNOR2_X1  g189(.A(G2451), .B(G2454), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT16), .ZN(new_n616));
  XNOR2_X1  g191(.A(G1341), .B(G1348), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n614), .B(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(G2443), .B(G2446), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  NAND3_X1  g197(.A1(new_n621), .A2(new_n622), .A3(G14), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(KEYINPUT77), .Z(G401));
  XOR2_X1   g199(.A(G2072), .B(G2078), .Z(new_n625));
  XOR2_X1   g200(.A(G2084), .B(G2090), .Z(new_n626));
  XNOR2_X1  g201(.A(G2067), .B(G2678), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n625), .B1(new_n628), .B2(KEYINPUT18), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT78), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2100), .ZN(new_n631));
  INV_X1    g206(.A(KEYINPUT18), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n628), .A2(KEYINPUT17), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n626), .A2(new_n627), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(new_n635), .B(G2096), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n631), .B(new_n636), .ZN(G227));
  XOR2_X1   g212(.A(G1971), .B(G1976), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT19), .ZN(new_n639));
  XOR2_X1   g214(.A(G1956), .B(G2474), .Z(new_n640));
  XOR2_X1   g215(.A(G1961), .B(G1966), .Z(new_n641));
  AND2_X1   g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(KEYINPUT79), .B(KEYINPUT20), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n640), .A2(new_n641), .ZN(new_n646));
  AND2_X1   g221(.A1(new_n639), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n639), .A2(new_n642), .A3(new_n646), .ZN(new_n648));
  NOR3_X1   g223(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G1981), .ZN(new_n650));
  INV_X1    g225(.A(G1986), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  AND2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n652), .A2(new_n654), .ZN(new_n656));
  XNOR2_X1  g231(.A(G1991), .B(G1996), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OR3_X1    g233(.A1(new_n655), .A2(new_n656), .A3(new_n658), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n658), .B1(new_n655), .B2(new_n656), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(G229));
  INV_X1    g236(.A(KEYINPUT94), .ZN(new_n662));
  INV_X1    g237(.A(G29), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n663), .A2(G35), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT91), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n665), .B1(new_n480), .B2(G29), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT29), .ZN(new_n667));
  INV_X1    g242(.A(G2090), .ZN(new_n668));
  OR3_X1    g243(.A1(new_n667), .A2(KEYINPUT92), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(KEYINPUT92), .B1(new_n667), .B2(new_n668), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(G16), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n672), .A2(G20), .ZN(new_n673));
  XOR2_X1   g248(.A(new_n673), .B(KEYINPUT23), .Z(new_n674));
  AOI21_X1  g249(.A(new_n674), .B1(G299), .B2(G16), .ZN(new_n675));
  XOR2_X1   g250(.A(KEYINPUT93), .B(G1956), .Z(new_n676));
  XOR2_X1   g251(.A(new_n675), .B(new_n676), .Z(new_n677));
  AOI21_X1  g252(.A(new_n662), .B1(new_n671), .B2(new_n677), .ZN(new_n678));
  INV_X1    g253(.A(G21), .ZN(new_n679));
  AOI21_X1  g254(.A(KEYINPUT87), .B1(new_n672), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n680), .B1(G286), .B2(new_n672), .ZN(new_n681));
  NAND3_X1  g256(.A1(G168), .A2(KEYINPUT87), .A3(G16), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(G1966), .ZN(new_n684));
  INV_X1    g259(.A(G1966), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  XNOR2_X1  g261(.A(KEYINPUT30), .B(G28), .ZN(new_n687));
  OR2_X1    g262(.A1(KEYINPUT31), .A2(G11), .ZN(new_n688));
  NAND2_X1  g263(.A1(KEYINPUT31), .A2(G11), .ZN(new_n689));
  AOI22_X1  g264(.A1(new_n687), .A2(new_n663), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(new_n605), .B2(new_n663), .ZN(new_n691));
  AND2_X1   g266(.A1(new_n672), .A2(G5), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n692), .B1(G301), .B2(G16), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g269(.A(new_n691), .B1(new_n694), .B2(G1961), .ZN(new_n695));
  NAND3_X1  g270(.A1(new_n684), .A2(new_n686), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT88), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(new_n678), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n671), .A2(new_n662), .A3(new_n677), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n672), .A2(G4), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n702), .B1(new_n584), .B2(new_n672), .ZN(new_n703));
  AOI22_X1  g278(.A1(new_n667), .A2(new_n668), .B1(new_n703), .B2(G1348), .ZN(new_n704));
  INV_X1    g279(.A(G1961), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n693), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(KEYINPUT24), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n663), .B1(new_n707), .B2(G34), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n708), .B1(new_n707), .B2(G34), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G160), .B2(G29), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT86), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT26), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(G129), .B2(new_n472), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n458), .A2(G105), .A3(G2104), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT85), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT85), .ZN(new_n718));
  NAND4_X1  g293(.A1(new_n718), .A2(new_n458), .A3(G105), .A4(G2104), .ZN(new_n719));
  AOI22_X1  g294(.A1(new_n473), .A2(G141), .B1(new_n717), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n715), .A2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g297(.A1(new_n722), .A2(new_n663), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n723), .B1(new_n663), .B2(G32), .ZN(new_n724));
  OAI221_X1 g299(.A(new_n706), .B1(G2084), .B2(new_n710), .C1(new_n712), .C2(new_n724), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT89), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g302(.A1(new_n704), .A2(new_n727), .ZN(new_n728));
  OAI22_X1  g303(.A1(new_n725), .A2(new_n726), .B1(new_n703), .B2(G1348), .ZN(new_n729));
  AND2_X1   g304(.A1(new_n710), .A2(G2084), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n458), .A2(G103), .A3(G2104), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT25), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n473), .A2(G139), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n464), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n733), .B(new_n734), .C1(new_n735), .C2(new_n458), .ZN(new_n736));
  MUX2_X1   g311(.A(G33), .B(new_n736), .S(G29), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G2072), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n663), .A2(G27), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT90), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n739), .A2(KEYINPUT90), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n740), .B(new_n741), .C1(G164), .C2(new_n663), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n738), .B1(G2078), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n663), .A2(G26), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT28), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n473), .A2(G140), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n472), .A2(G128), .ZN(new_n747));
  OR2_X1    g322(.A1(G104), .A2(G2105), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n748), .B(G2104), .C1(G116), .C2(new_n458), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n746), .A2(new_n747), .A3(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n745), .B1(new_n751), .B2(new_n663), .ZN(new_n752));
  AOI211_X1 g327(.A(new_n730), .B(new_n743), .C1(G2067), .C2(new_n752), .ZN(new_n753));
  NOR2_X1   g328(.A1(new_n737), .A2(G2072), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT84), .ZN(new_n755));
  NOR2_X1   g330(.A1(new_n752), .A2(G2067), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n742), .A2(G2078), .ZN(new_n757));
  AOI211_X1 g332(.A(new_n756), .B(new_n757), .C1(new_n724), .C2(new_n712), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n753), .A2(new_n755), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n672), .A2(G19), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(new_n537), .B2(new_n672), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G1341), .ZN(new_n762));
  NOR3_X1   g337(.A1(new_n729), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NAND3_X1  g338(.A1(new_n701), .A2(new_n728), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT95), .B1(new_n700), .B2(new_n764), .ZN(new_n765));
  INV_X1    g340(.A(new_n764), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT95), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n766), .A2(new_n699), .A3(new_n767), .ZN(new_n768));
  MUX2_X1   g343(.A(G6), .B(G305), .S(G16), .Z(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT32), .ZN(new_n770));
  INV_X1    g345(.A(G1981), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n672), .A2(G22), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(G166), .B2(new_n672), .ZN(new_n774));
  INV_X1    g349(.A(G1971), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n776), .A2(KEYINPUT83), .ZN(new_n777));
  NOR2_X1   g352(.A1(new_n776), .A2(KEYINPUT83), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n672), .A2(G23), .ZN(new_n779));
  INV_X1    g354(.A(G288), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(new_n672), .ZN(new_n781));
  XOR2_X1   g356(.A(KEYINPUT33), .B(G1976), .Z(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n778), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g359(.A1(new_n772), .A2(new_n777), .A3(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n785), .A2(KEYINPUT34), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G24), .ZN(new_n788));
  XOR2_X1   g363(.A(G290), .B(KEYINPUT82), .Z(new_n789));
  AOI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(G16), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(new_n651), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n473), .A2(G131), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n472), .A2(G119), .ZN(new_n793));
  NOR2_X1   g368(.A1(new_n458), .A2(G107), .ZN(new_n794));
  OAI21_X1  g369(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n795));
  OAI211_X1 g370(.A(new_n792), .B(new_n793), .C1(new_n794), .C2(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G25), .B(new_n796), .S(G29), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT35), .B(G1991), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT81), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n797), .B(new_n799), .Z(new_n800));
  NAND4_X1  g375(.A1(new_n786), .A2(new_n787), .A3(new_n791), .A4(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(KEYINPUT36), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n765), .A2(new_n768), .B1(new_n802), .B2(new_n803), .ZN(G311));
  NAND2_X1  g379(.A1(new_n765), .A2(new_n768), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n802), .A2(new_n803), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(G150));
  NAND2_X1  g382(.A1(new_n584), .A2(G559), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT38), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n810));
  INV_X1    g385(.A(G93), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n810), .A2(new_n502), .B1(new_n811), .B2(new_n505), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G55), .B2(new_n524), .ZN(new_n813));
  XOR2_X1   g388(.A(new_n537), .B(new_n813), .Z(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n809), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(KEYINPUT39), .ZN(new_n817));
  AOI21_X1  g392(.A(G860), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(new_n817), .B2(new_n816), .ZN(new_n819));
  INV_X1    g394(.A(new_n813), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n820), .A2(G860), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT96), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n819), .A2(new_n823), .ZN(G145));
  XNOR2_X1  g399(.A(new_n721), .B(new_n736), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(new_n598), .ZN(new_n826));
  XNOR2_X1  g401(.A(G164), .B(new_n750), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n472), .A2(G130), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n458), .A2(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n832), .B1(G142), .B2(new_n473), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(new_n796), .Z(new_n834));
  OR2_X1    g409(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT97), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n828), .A2(new_n834), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n835), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(G160), .B(new_n605), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n480), .B(new_n839), .Z(new_n840));
  AOI21_X1  g415(.A(G37), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n840), .ZN(new_n842));
  NAND4_X1  g417(.A1(new_n835), .A2(new_n836), .A3(new_n842), .A4(new_n837), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT98), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n841), .A2(KEYINPUT98), .A3(new_n843), .ZN(new_n847));
  AND3_X1   g422(.A1(new_n846), .A2(KEYINPUT40), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(KEYINPUT40), .B1(new_n846), .B2(new_n847), .ZN(new_n849));
  NOR2_X1   g424(.A1(new_n848), .A2(new_n849), .ZN(G395));
  NAND2_X1  g425(.A1(new_n820), .A2(new_n575), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n592), .B(new_n815), .ZN(new_n852));
  OR2_X1    g427(.A1(new_n581), .A2(G299), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n581), .A2(G299), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n852), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(KEYINPUT41), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT41), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n853), .A2(new_n858), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  OAI21_X1  g435(.A(new_n856), .B1(new_n852), .B2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(G290), .B(G305), .ZN(new_n862));
  XNOR2_X1  g437(.A(G303), .B(G288), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n863), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n867), .A2(KEYINPUT42), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n869));
  INV_X1    g444(.A(new_n866), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(new_n864), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n865), .A2(KEYINPUT99), .A3(new_n866), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n868), .B1(new_n873), .B2(KEYINPUT42), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n861), .B(new_n874), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n851), .B1(new_n875), .B2(new_n575), .ZN(G295));
  OAI21_X1  g451(.A(new_n851), .B1(new_n875), .B2(new_n575), .ZN(G331));
  INV_X1    g452(.A(new_n873), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT103), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n857), .A2(new_n879), .A3(new_n859), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n859), .A2(new_n879), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT100), .ZN(new_n883));
  NAND2_X1  g458(.A1(G301), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(G171), .A2(KEYINPUT100), .ZN(new_n885));
  NAND4_X1  g460(.A1(new_n553), .A2(new_n555), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n883), .B(G301), .C1(new_n526), .C2(new_n528), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(KEYINPUT101), .A3(new_n815), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT101), .B1(new_n888), .B2(new_n815), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n886), .A2(new_n887), .A3(new_n814), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT102), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT102), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n886), .A2(new_n887), .A3(new_n814), .A4(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g472(.A(new_n882), .B1(new_n892), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n888), .A2(new_n815), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n893), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT104), .B1(new_n900), .B2(new_n855), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT104), .ZN(new_n902));
  INV_X1    g477(.A(new_n855), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n899), .A2(new_n902), .A3(new_n903), .A4(new_n893), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n901), .A2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n878), .B1(new_n898), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT43), .ZN(new_n907));
  INV_X1    g482(.A(G37), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT101), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n899), .A2(new_n909), .ZN(new_n910));
  NAND4_X1  g485(.A1(new_n897), .A2(new_n910), .A3(new_n903), .A4(new_n889), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n900), .A2(new_n860), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n911), .A2(new_n873), .A3(new_n912), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT44), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n913), .A2(new_n908), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n873), .B1(new_n911), .B2(new_n912), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  AND3_X1   g493(.A1(new_n914), .A2(new_n915), .A3(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(new_n916), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT105), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n911), .A2(new_n912), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n878), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n920), .A2(new_n921), .A3(new_n907), .A4(new_n923), .ZN(new_n924));
  NAND4_X1  g499(.A1(new_n923), .A2(new_n907), .A3(new_n908), .A4(new_n913), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(KEYINPUT105), .ZN(new_n926));
  AND3_X1   g501(.A1(new_n906), .A2(new_n908), .A3(new_n913), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n924), .B(new_n926), .C1(new_n927), .C2(new_n907), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n919), .B1(new_n928), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g504(.A1(new_n492), .A2(new_n494), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n484), .A2(new_n487), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(G1384), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT45), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  XOR2_X1   g511(.A(KEYINPUT106), .B(G40), .Z(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(G160), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n750), .B(G2067), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n942), .B(KEYINPUT108), .Z(new_n943));
  INV_X1    g518(.A(G1996), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n722), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n943), .B1(new_n940), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n940), .A2(new_n944), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n947), .B(KEYINPUT107), .Z(new_n948));
  OR2_X1    g523(.A1(new_n948), .A2(new_n721), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n796), .B(new_n799), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n940), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  XNOR2_X1  g527(.A(G290), .B(G1986), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n952), .B1(new_n940), .B2(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT120), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT109), .B1(G164), .B2(G1384), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n932), .A2(new_n957), .A3(new_n933), .ZN(new_n958));
  AOI21_X1  g533(.A(KEYINPUT45), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n932), .A2(KEYINPUT45), .A3(new_n933), .ZN(new_n960));
  NOR3_X1   g535(.A1(new_n467), .A2(new_n470), .A3(new_n937), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n685), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n939), .B1(KEYINPUT50), .B2(new_n934), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n956), .A2(new_n958), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n964), .B1(KEYINPUT50), .B2(new_n965), .ZN(new_n966));
  XOR2_X1   g541(.A(KEYINPUT114), .B(G2084), .Z(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  OAI211_X1 g543(.A(new_n955), .B(G8), .C1(new_n968), .C2(G286), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT121), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n969), .A2(new_n970), .A3(KEYINPUT51), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n968), .A2(G8), .A3(G286), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n969), .A2(new_n970), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT51), .ZN(new_n975));
  OAI211_X1 g550(.A(KEYINPUT121), .B(G8), .C1(new_n968), .C2(G286), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n966), .A2(new_n705), .ZN(new_n978));
  INV_X1    g553(.A(G2078), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n936), .A2(new_n979), .A3(new_n961), .A4(new_n960), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT53), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT122), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT122), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n980), .A2(new_n984), .A3(new_n981), .ZN(new_n985));
  AND2_X1   g560(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n986));
  NOR2_X1   g561(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n987));
  OAI211_X1 g562(.A(KEYINPUT53), .B(G40), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n467), .A2(new_n470), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n936), .A2(new_n960), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT124), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n936), .A2(KEYINPUT124), .A3(new_n960), .A4(new_n989), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n978), .A2(new_n983), .A3(new_n985), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(G171), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n995), .A2(KEYINPUT127), .A3(G171), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n959), .ZN(new_n1001));
  INV_X1    g576(.A(new_n962), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n1001), .A2(KEYINPUT53), .A3(new_n979), .A4(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n978), .A2(new_n983), .A3(new_n985), .A4(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n1004), .A2(G171), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT54), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  AOI22_X1  g582(.A1(new_n973), .A2(new_n977), .B1(new_n1000), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n780), .A2(G1976), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n956), .A2(new_n961), .A3(new_n958), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1009), .A2(new_n1010), .A3(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT52), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1012), .B1(new_n780), .B2(G1976), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n564), .A2(new_n771), .A3(new_n567), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n771), .B1(new_n564), .B2(new_n567), .ZN(new_n1018));
  OAI21_X1  g593(.A(new_n1015), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1018), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1020), .A2(KEYINPUT49), .A3(new_n1016), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n1019), .A2(new_n1021), .A3(G8), .A4(new_n1010), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1011), .A2(KEYINPUT52), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1014), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G8), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1002), .A2(new_n936), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1026), .A2(new_n775), .ZN(new_n1027));
  XOR2_X1   g602(.A(KEYINPUT110), .B(G2090), .Z(new_n1028));
  OAI211_X1 g603(.A(new_n964), .B(new_n1028), .C1(KEYINPUT50), .C2(new_n965), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(G166), .B2(new_n1025), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1024), .B1(new_n1030), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT113), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT50), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1038), .B1(new_n956), .B2(new_n958), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1037), .B1(new_n1039), .B2(new_n939), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n957), .B1(new_n932), .B2(new_n933), .ZN(new_n1041));
  AOI211_X1 g616(.A(KEYINPUT109), .B(G1384), .C1(new_n930), .C2(new_n931), .ZN(new_n1042));
  OAI21_X1  g617(.A(KEYINPUT50), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1043), .A2(KEYINPUT113), .A3(new_n961), .ZN(new_n1044));
  NOR2_X1   g619(.A1(new_n934), .A2(KEYINPUT50), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1040), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(new_n1028), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1027), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  AND2_X1   g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  OAI211_X1 g625(.A(new_n1036), .B(KEYINPUT126), .C1(new_n1050), .C2(new_n1034), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT126), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1030), .A2(new_n1035), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1053), .A2(new_n1022), .A3(new_n1014), .A4(new_n1023), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1034), .B1(new_n1049), .B2(G8), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1052), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  AND2_X1   g631(.A1(new_n1051), .A2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1004), .A2(G171), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n705), .A2(new_n966), .B1(new_n982), .B2(KEYINPUT122), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(G301), .A3(new_n985), .A4(new_n994), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1006), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(KEYINPUT125), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT125), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1061), .A2(new_n1064), .A3(new_n1006), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1063), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1008), .A2(new_n1057), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT118), .ZN(new_n1068));
  XOR2_X1   g643(.A(KEYINPUT56), .B(G2072), .Z(new_n1069));
  NOR2_X1   g644(.A1(new_n1026), .A2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(G1956), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1070), .B1(new_n1047), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT57), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g651(.A1(G299), .A2(new_n1073), .A3(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n545), .A2(new_n1074), .A3(new_n1075), .A4(new_n550), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(new_n1079), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1068), .B1(new_n1072), .B2(new_n1080), .ZN(new_n1081));
  AOI211_X1 g656(.A(new_n1079), .B(new_n1070), .C1(new_n1047), .C2(new_n1071), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n939), .B1(new_n965), .B2(KEYINPUT50), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1045), .B1(new_n1084), .B2(KEYINPUT113), .ZN(new_n1085));
  AOI21_X1  g660(.A(G1956), .B1(new_n1085), .B2(new_n1040), .ZN(new_n1086));
  OAI211_X1 g661(.A(KEYINPUT118), .B(new_n1079), .C1(new_n1086), .C2(new_n1070), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT61), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1083), .A2(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1079), .B1(new_n1086), .B2(new_n1070), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1072), .A2(new_n1080), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1091), .A2(new_n1092), .A3(KEYINPUT61), .ZN(new_n1093));
  INV_X1    g668(.A(KEYINPUT116), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1010), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n956), .A2(new_n958), .A3(KEYINPUT116), .A4(new_n961), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(KEYINPUT58), .B(G1341), .ZN(new_n1098));
  OAI22_X1  g673(.A1(new_n1097), .A2(new_n1098), .B1(G1996), .B2(new_n1026), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n537), .ZN(new_n1100));
  XOR2_X1   g675(.A(KEYINPUT117), .B(KEYINPUT59), .Z(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1101), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1099), .A2(new_n537), .A3(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1102), .A2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1093), .A2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(KEYINPUT119), .B1(new_n1090), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g682(.A(new_n1088), .B(new_n1087), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT119), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n1108), .A2(new_n1093), .A3(new_n1109), .A4(new_n1105), .ZN(new_n1110));
  INV_X1    g685(.A(G2067), .ZN(new_n1111));
  INV_X1    g686(.A(G1348), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1111), .A2(new_n1097), .B1(new_n966), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n584), .A2(KEYINPUT60), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1113), .B(new_n1114), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1115), .B1(KEYINPUT60), .B2(new_n584), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1107), .A2(new_n1110), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1091), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1113), .B1(new_n583), .B2(new_n582), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1118), .B1(new_n1092), .B2(new_n1119), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1067), .B1(new_n1117), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1058), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n973), .A2(KEYINPUT62), .A3(new_n977), .ZN(new_n1123));
  AOI21_X1  g698(.A(KEYINPUT62), .B1(new_n973), .B2(new_n977), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1057), .B(new_n1122), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1125));
  NOR2_X1   g700(.A1(G288), .A2(G1976), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1017), .B1(new_n1022), .B2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1010), .A2(G8), .ZN(new_n1128));
  XNOR2_X1  g703(.A(new_n1128), .B(KEYINPUT112), .ZN(new_n1129));
  OAI22_X1  g704(.A1(new_n1053), .A2(new_n1024), .B1(new_n1127), .B2(new_n1129), .ZN(new_n1130));
  AND3_X1   g705(.A1(new_n968), .A2(G8), .A3(G168), .ZN(new_n1131));
  OAI211_X1 g706(.A(new_n1036), .B(new_n1131), .C1(new_n1050), .C2(new_n1034), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT63), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OR2_X1    g709(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1135));
  NAND4_X1  g710(.A1(new_n1036), .A2(KEYINPUT63), .A3(new_n1131), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1130), .B1(new_n1134), .B2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1125), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n954), .B1(new_n1121), .B2(new_n1138), .ZN(new_n1139));
  NOR4_X1   g714(.A1(G290), .A2(G1986), .A3(new_n936), .A4(new_n939), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n1140), .B(KEYINPUT48), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n952), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n940), .B1(new_n941), .B2(new_n721), .ZN(new_n1143));
  AND2_X1   g718(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n1144));
  NOR2_X1   g719(.A1(new_n948), .A2(KEYINPUT46), .ZN(new_n1145));
  OAI21_X1  g720(.A(new_n1143), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  XOR2_X1   g721(.A(new_n1146), .B(KEYINPUT47), .Z(new_n1147));
  NAND2_X1  g722(.A1(new_n946), .A2(new_n949), .ZN(new_n1148));
  OR2_X1    g723(.A1(new_n796), .A2(new_n799), .ZN(new_n1149));
  OAI22_X1  g724(.A1(new_n1148), .A2(new_n1149), .B1(G2067), .B2(new_n750), .ZN(new_n1150));
  AOI211_X1 g725(.A(new_n1142), .B(new_n1147), .C1(new_n940), .C2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1139), .A2(new_n1151), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g727(.A(G319), .ZN(new_n1154));
  NOR3_X1   g728(.A1(G401), .A2(new_n1154), .A3(G227), .ZN(new_n1155));
  NAND3_X1  g729(.A1(new_n659), .A2(new_n1155), .A3(new_n660), .ZN(new_n1156));
  INV_X1    g730(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g731(.A1(new_n846), .A2(new_n847), .ZN(new_n1158));
  NAND2_X1  g732(.A1(new_n914), .A2(new_n918), .ZN(new_n1159));
  NAND3_X1  g733(.A1(new_n1157), .A2(new_n1158), .A3(new_n1159), .ZN(G225));
  INV_X1    g734(.A(G225), .ZN(G308));
endmodule


