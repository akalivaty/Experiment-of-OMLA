

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591;

  XNOR2_X1 U327 ( .A(n410), .B(n409), .ZN(n532) );
  XNOR2_X1 U328 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U329 ( .A(n363), .B(n362), .ZN(n369) );
  XNOR2_X1 U330 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n409) );
  XNOR2_X1 U331 ( .A(KEYINPUT55), .B(KEYINPUT118), .ZN(n432) );
  XNOR2_X1 U332 ( .A(n433), .B(n432), .ZN(n451) );
  XNOR2_X1 U333 ( .A(n453), .B(G183GAT), .ZN(n454) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(G1350GAT) );
  XOR2_X1 U335 ( .A(G162GAT), .B(G57GAT), .Z(n296) );
  XNOR2_X1 U336 ( .A(G29GAT), .B(G85GAT), .ZN(n295) );
  XNOR2_X1 U337 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U338 ( .A(G155GAT), .B(G148GAT), .Z(n298) );
  XNOR2_X1 U339 ( .A(G1GAT), .B(G120GAT), .ZN(n297) );
  XNOR2_X1 U340 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U341 ( .A(n300), .B(n299), .Z(n310) );
  XOR2_X1 U342 ( .A(KEYINPUT6), .B(KEYINPUT1), .Z(n302) );
  XNOR2_X1 U343 ( .A(KEYINPUT5), .B(KEYINPUT87), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n308) );
  XOR2_X1 U345 ( .A(KEYINPUT2), .B(KEYINPUT83), .Z(n304) );
  XNOR2_X1 U346 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n424) );
  XOR2_X1 U348 ( .A(G134GAT), .B(KEYINPUT76), .Z(n359) );
  XOR2_X1 U349 ( .A(n424), .B(n359), .Z(n306) );
  NAND2_X1 U350 ( .A1(G225GAT), .A2(G233GAT), .ZN(n305) );
  XNOR2_X1 U351 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U352 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U354 ( .A(n311), .B(KEYINPUT88), .Z(n314) );
  XNOR2_X1 U355 ( .A(G113GAT), .B(G127GAT), .ZN(n312) );
  XNOR2_X1 U356 ( .A(n312), .B(KEYINPUT0), .ZN(n435) );
  XNOR2_X1 U357 ( .A(n435), .B(KEYINPUT4), .ZN(n313) );
  XNOR2_X1 U358 ( .A(n314), .B(n313), .ZN(n502) );
  XOR2_X1 U359 ( .A(KEYINPUT117), .B(KEYINPUT54), .Z(n412) );
  XOR2_X1 U360 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n316) );
  XNOR2_X1 U361 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n316), .B(n315), .ZN(n438) );
  XOR2_X1 U363 ( .A(G204GAT), .B(G64GAT), .Z(n318) );
  XNOR2_X1 U364 ( .A(G176GAT), .B(G92GAT), .ZN(n317) );
  XNOR2_X1 U365 ( .A(n318), .B(n317), .ZN(n349) );
  XOR2_X1 U366 ( .A(KEYINPUT89), .B(n349), .Z(n320) );
  NAND2_X1 U367 ( .A1(G226GAT), .A2(G233GAT), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n323) );
  XOR2_X1 U369 ( .A(KEYINPUT21), .B(G211GAT), .Z(n322) );
  XNOR2_X1 U370 ( .A(G197GAT), .B(G218GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n420) );
  XOR2_X1 U372 ( .A(n323), .B(n420), .Z(n325) );
  XOR2_X1 U373 ( .A(G36GAT), .B(G190GAT), .Z(n361) );
  XOR2_X1 U374 ( .A(G8GAT), .B(G183GAT), .Z(n376) );
  XNOR2_X1 U375 ( .A(n361), .B(n376), .ZN(n324) );
  XNOR2_X1 U376 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U377 ( .A(n438), .B(n326), .ZN(n505) );
  XOR2_X1 U378 ( .A(G197GAT), .B(G141GAT), .Z(n328) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(KEYINPUT72), .ZN(n327) );
  XNOR2_X1 U380 ( .A(n328), .B(n327), .ZN(n344) );
  XOR2_X1 U381 ( .A(KEYINPUT70), .B(G113GAT), .Z(n330) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(G22GAT), .ZN(n329) );
  XNOR2_X1 U383 ( .A(n330), .B(n329), .ZN(n331) );
  XOR2_X1 U384 ( .A(n331), .B(G50GAT), .Z(n333) );
  XOR2_X1 U385 ( .A(G15GAT), .B(G1GAT), .Z(n384) );
  XNOR2_X1 U386 ( .A(n384), .B(G36GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U388 ( .A(KEYINPUT71), .B(KEYINPUT30), .Z(n335) );
  NAND2_X1 U389 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U390 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n342) );
  XOR2_X1 U392 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n339) );
  XNOR2_X1 U393 ( .A(G43GAT), .B(G29GAT), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U395 ( .A(KEYINPUT73), .B(n340), .Z(n372) );
  XOR2_X1 U396 ( .A(n372), .B(KEYINPUT29), .Z(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U398 ( .A(n344), .B(n343), .Z(n562) );
  INV_X1 U399 ( .A(n562), .ZN(n577) );
  XOR2_X1 U400 ( .A(G99GAT), .B(G85GAT), .Z(n367) );
  XOR2_X1 U401 ( .A(KEYINPUT13), .B(G57GAT), .Z(n383) );
  XNOR2_X1 U402 ( .A(n367), .B(n383), .ZN(n356) );
  XOR2_X1 U403 ( .A(KEYINPUT74), .B(KEYINPUT32), .Z(n346) );
  NAND2_X1 U404 ( .A1(G230GAT), .A2(G233GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U406 ( .A(n347), .B(KEYINPUT75), .Z(n351) );
  XNOR2_X1 U407 ( .A(G106GAT), .B(G78GAT), .ZN(n348) );
  XNOR2_X1 U408 ( .A(n348), .B(G148GAT), .ZN(n421) );
  XNOR2_X1 U409 ( .A(n421), .B(n349), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U411 ( .A(KEYINPUT31), .B(n352), .Z(n354) );
  XOR2_X1 U412 ( .A(G71GAT), .B(G120GAT), .Z(n434) );
  XNOR2_X1 U413 ( .A(n434), .B(KEYINPUT33), .ZN(n353) );
  XNOR2_X1 U414 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n580) );
  INV_X1 U416 ( .A(KEYINPUT45), .ZN(n396) );
  INV_X1 U417 ( .A(KEYINPUT36), .ZN(n375) );
  XOR2_X1 U418 ( .A(KEYINPUT9), .B(KEYINPUT10), .Z(n358) );
  XNOR2_X1 U419 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n371) );
  XOR2_X1 U421 ( .A(G50GAT), .B(G162GAT), .Z(n427) );
  XNOR2_X1 U422 ( .A(n427), .B(n359), .ZN(n363) );
  XNOR2_X1 U423 ( .A(KEYINPUT68), .B(G218GAT), .ZN(n360) );
  XOR2_X1 U424 ( .A(KEYINPUT69), .B(G92GAT), .Z(n365) );
  NAND2_X1 U425 ( .A1(G232GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U426 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U427 ( .A(n367), .B(n366), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U429 ( .A(n371), .B(n370), .ZN(n374) );
  INV_X1 U430 ( .A(n372), .ZN(n373) );
  XOR2_X1 U431 ( .A(n374), .B(n373), .Z(n402) );
  XNOR2_X1 U432 ( .A(n375), .B(n402), .ZN(n482) );
  XOR2_X1 U433 ( .A(KEYINPUT14), .B(KEYINPUT12), .Z(n378) );
  XOR2_X1 U434 ( .A(G22GAT), .B(G155GAT), .Z(n426) );
  XNOR2_X1 U435 ( .A(n376), .B(n426), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U437 ( .A(G64GAT), .B(G78GAT), .Z(n380) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n394) );
  XOR2_X1 U443 ( .A(KEYINPUT15), .B(KEYINPUT80), .Z(n388) );
  XNOR2_X1 U444 ( .A(G71GAT), .B(G127GAT), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n388), .B(n387), .ZN(n392) );
  XOR2_X1 U446 ( .A(G211GAT), .B(KEYINPUT79), .Z(n390) );
  XNOR2_X1 U447 ( .A(KEYINPUT77), .B(KEYINPUT78), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n392), .B(n391), .Z(n393) );
  XNOR2_X1 U450 ( .A(n394), .B(n393), .ZN(n584) );
  NOR2_X1 U451 ( .A1(n482), .A2(n584), .ZN(n395) );
  XNOR2_X1 U452 ( .A(n396), .B(n395), .ZN(n397) );
  NOR2_X1 U453 ( .A1(n580), .A2(n397), .ZN(n398) );
  NAND2_X1 U454 ( .A1(n577), .A2(n398), .ZN(n408) );
  XOR2_X1 U455 ( .A(KEYINPUT41), .B(KEYINPUT65), .Z(n399) );
  XNOR2_X1 U456 ( .A(n399), .B(n580), .ZN(n499) );
  NOR2_X1 U457 ( .A1(n577), .A2(n499), .ZN(n401) );
  INV_X1 U458 ( .A(KEYINPUT46), .ZN(n400) );
  XNOR2_X1 U459 ( .A(n401), .B(n400), .ZN(n404) );
  INV_X1 U460 ( .A(n402), .ZN(n560) );
  INV_X1 U461 ( .A(n584), .ZN(n541) );
  NOR2_X1 U462 ( .A1(n402), .A2(n541), .ZN(n403) );
  NAND2_X1 U463 ( .A1(n404), .A2(n403), .ZN(n406) );
  XOR2_X1 U464 ( .A(KEYINPUT47), .B(KEYINPUT108), .Z(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  NAND2_X1 U466 ( .A1(n408), .A2(n407), .ZN(n410) );
  NAND2_X1 U467 ( .A1(n505), .A2(n532), .ZN(n411) );
  XNOR2_X1 U468 ( .A(n412), .B(n411), .ZN(n413) );
  NOR2_X1 U469 ( .A1(n502), .A2(n413), .ZN(n414) );
  XNOR2_X1 U470 ( .A(n414), .B(KEYINPUT66), .ZN(n576) );
  XOR2_X1 U471 ( .A(KEYINPUT84), .B(KEYINPUT23), .Z(n416) );
  XNOR2_X1 U472 ( .A(G204GAT), .B(KEYINPUT85), .ZN(n415) );
  XNOR2_X1 U473 ( .A(n416), .B(n415), .ZN(n431) );
  XOR2_X1 U474 ( .A(KEYINPUT86), .B(KEYINPUT22), .Z(n418) );
  NAND2_X1 U475 ( .A1(G228GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U476 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U477 ( .A(n419), .B(KEYINPUT24), .Z(n423) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U479 ( .A(n423), .B(n422), .ZN(n425) );
  XOR2_X1 U480 ( .A(n425), .B(n424), .Z(n429) );
  XNOR2_X1 U481 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n430) );
  XOR2_X1 U483 ( .A(n431), .B(n430), .Z(n466) );
  NAND2_X1 U484 ( .A1(n576), .A2(n466), .ZN(n433) );
  XOR2_X1 U485 ( .A(n435), .B(n434), .Z(n437) );
  XNOR2_X1 U486 ( .A(G99GAT), .B(G190GAT), .ZN(n436) );
  XNOR2_X1 U487 ( .A(n437), .B(n436), .ZN(n442) );
  XOR2_X1 U488 ( .A(n438), .B(KEYINPUT81), .Z(n440) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U490 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U491 ( .A(n442), .B(n441), .Z(n450) );
  XOR2_X1 U492 ( .A(G183GAT), .B(G134GAT), .Z(n444) );
  XNOR2_X1 U493 ( .A(G43GAT), .B(G15GAT), .ZN(n443) );
  XNOR2_X1 U494 ( .A(n444), .B(n443), .ZN(n448) );
  XOR2_X1 U495 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n446) );
  XNOR2_X1 U496 ( .A(G176GAT), .B(KEYINPUT67), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U498 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U499 ( .A(n450), .B(n449), .ZN(n534) );
  NAND2_X1 U500 ( .A1(n451), .A2(n534), .ZN(n452) );
  XNOR2_X1 U501 ( .A(n452), .B(KEYINPUT119), .ZN(n570) );
  NAND2_X1 U502 ( .A1(n570), .A2(n541), .ZN(n455) );
  XOR2_X1 U503 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n453) );
  INV_X1 U504 ( .A(n502), .ZN(n516) );
  NOR2_X1 U505 ( .A1(n580), .A2(n577), .ZN(n486) );
  NAND2_X1 U506 ( .A1(n534), .A2(n505), .ZN(n456) );
  XOR2_X1 U507 ( .A(KEYINPUT91), .B(n456), .Z(n457) );
  NAND2_X1 U508 ( .A1(n457), .A2(n466), .ZN(n458) );
  XNOR2_X1 U509 ( .A(n458), .B(KEYINPUT92), .ZN(n459) );
  XNOR2_X1 U510 ( .A(KEYINPUT25), .B(n459), .ZN(n463) );
  NOR2_X1 U511 ( .A1(n466), .A2(n534), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT26), .ZN(n575) );
  INV_X1 U513 ( .A(n575), .ZN(n461) );
  XOR2_X1 U514 ( .A(KEYINPUT27), .B(n505), .Z(n465) );
  NOR2_X1 U515 ( .A1(n461), .A2(n465), .ZN(n462) );
  NOR2_X1 U516 ( .A1(n463), .A2(n462), .ZN(n464) );
  NOR2_X1 U517 ( .A1(n502), .A2(n464), .ZN(n470) );
  NOR2_X1 U518 ( .A1(n516), .A2(n465), .ZN(n531) );
  XOR2_X1 U519 ( .A(n466), .B(KEYINPUT28), .Z(n537) );
  INV_X1 U520 ( .A(n537), .ZN(n527) );
  NAND2_X1 U521 ( .A1(n531), .A2(n527), .ZN(n467) );
  XNOR2_X1 U522 ( .A(KEYINPUT90), .B(n467), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n534), .A2(n468), .ZN(n469) );
  NOR2_X1 U524 ( .A1(n470), .A2(n469), .ZN(n483) );
  NOR2_X1 U525 ( .A1(n402), .A2(n584), .ZN(n471) );
  XOR2_X1 U526 ( .A(KEYINPUT16), .B(n471), .Z(n472) );
  NOR2_X1 U527 ( .A1(n483), .A2(n472), .ZN(n500) );
  NAND2_X1 U528 ( .A1(n486), .A2(n500), .ZN(n479) );
  NOR2_X1 U529 ( .A1(n516), .A2(n479), .ZN(n473) );
  XOR2_X1 U530 ( .A(G1GAT), .B(n473), .Z(n474) );
  XNOR2_X1 U531 ( .A(KEYINPUT34), .B(n474), .ZN(G1324GAT) );
  INV_X1 U532 ( .A(n505), .ZN(n519) );
  NOR2_X1 U533 ( .A1(n519), .A2(n479), .ZN(n475) );
  XOR2_X1 U534 ( .A(G8GAT), .B(n475), .Z(G1325GAT) );
  INV_X1 U535 ( .A(n534), .ZN(n523) );
  NOR2_X1 U536 ( .A1(n523), .A2(n479), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT35), .B(KEYINPUT93), .ZN(n476) );
  XNOR2_X1 U538 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U539 ( .A(G15GAT), .B(n478), .Z(G1326GAT) );
  NOR2_X1 U540 ( .A1(n527), .A2(n479), .ZN(n480) );
  XOR2_X1 U541 ( .A(KEYINPUT94), .B(n480), .Z(n481) );
  XNOR2_X1 U542 ( .A(G22GAT), .B(n481), .ZN(G1327GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT38), .B(KEYINPUT95), .Z(n488) );
  NOR2_X1 U544 ( .A1(n482), .A2(n483), .ZN(n484) );
  NAND2_X1 U545 ( .A1(n584), .A2(n484), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n485), .B(KEYINPUT37), .ZN(n515) );
  NAND2_X1 U547 ( .A1(n486), .A2(n515), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n495) );
  NOR2_X1 U549 ( .A1(n495), .A2(n516), .ZN(n490) );
  XNOR2_X1 U550 ( .A(KEYINPUT39), .B(KEYINPUT96), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(n491), .ZN(G1328GAT) );
  NOR2_X1 U553 ( .A1(n519), .A2(n495), .ZN(n492) );
  XOR2_X1 U554 ( .A(G36GAT), .B(n492), .Z(G1329GAT) );
  NOR2_X1 U555 ( .A1(n495), .A2(n523), .ZN(n493) );
  XOR2_X1 U556 ( .A(KEYINPUT40), .B(n493), .Z(n494) );
  XNOR2_X1 U557 ( .A(G43GAT), .B(n494), .ZN(G1330GAT) );
  NOR2_X1 U558 ( .A1(n495), .A2(n527), .ZN(n497) );
  XNOR2_X1 U559 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U561 ( .A(G50GAT), .B(n498), .ZN(G1331GAT) );
  INV_X1 U562 ( .A(n499), .ZN(n565) );
  NOR2_X1 U563 ( .A1(n562), .A2(n499), .ZN(n514) );
  NAND2_X1 U564 ( .A1(n500), .A2(n514), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT99), .ZN(n509) );
  NAND2_X1 U566 ( .A1(n502), .A2(n509), .ZN(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT42), .B(n503), .ZN(n504) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(n504), .ZN(G1332GAT) );
  NAND2_X1 U569 ( .A1(n505), .A2(n509), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n506), .B(KEYINPUT100), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G64GAT), .B(n507), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n534), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT102), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n537), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT101), .Z(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n526) );
  NOR2_X1 U580 ( .A1(n516), .A2(n526), .ZN(n518) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT103), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n519), .A2(n526), .ZN(n521) );
  XNOR2_X1 U584 ( .A(KEYINPUT104), .B(KEYINPUT105), .ZN(n520) );
  XNOR2_X1 U585 ( .A(n521), .B(n520), .ZN(n522) );
  XNOR2_X1 U586 ( .A(G92GAT), .B(n522), .ZN(G1337GAT) );
  NOR2_X1 U587 ( .A1(n523), .A2(n526), .ZN(n524) );
  XOR2_X1 U588 ( .A(KEYINPUT106), .B(n524), .Z(n525) );
  XNOR2_X1 U589 ( .A(G99GAT), .B(n525), .ZN(G1338GAT) );
  NOR2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n529) );
  XNOR2_X1 U591 ( .A(KEYINPUT44), .B(KEYINPUT107), .ZN(n528) );
  XNOR2_X1 U592 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U593 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NAND2_X1 U594 ( .A1(n532), .A2(n531), .ZN(n533) );
  XNOR2_X1 U595 ( .A(n533), .B(KEYINPUT109), .ZN(n550) );
  NAND2_X1 U596 ( .A1(n534), .A2(n550), .ZN(n535) );
  XNOR2_X1 U597 ( .A(KEYINPUT110), .B(n535), .ZN(n536) );
  NOR2_X1 U598 ( .A1(n537), .A2(n536), .ZN(n546) );
  NAND2_X1 U599 ( .A1(n562), .A2(n546), .ZN(n538) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U602 ( .A1(n546), .A2(n565), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(KEYINPUT112), .ZN(n545) );
  XOR2_X1 U605 ( .A(KEYINPUT111), .B(KEYINPUT50), .Z(n543) );
  NAND2_X1 U606 ( .A1(n546), .A2(n541), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n545), .B(n544), .ZN(G1342GAT) );
  XOR2_X1 U609 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n548) );
  NAND2_X1 U610 ( .A1(n546), .A2(n402), .ZN(n547) );
  XNOR2_X1 U611 ( .A(n548), .B(n547), .ZN(n549) );
  XOR2_X1 U612 ( .A(G134GAT), .B(n549), .Z(G1343GAT) );
  NAND2_X1 U613 ( .A1(n550), .A2(n575), .ZN(n559) );
  NOR2_X1 U614 ( .A1(n577), .A2(n559), .ZN(n551) );
  XOR2_X1 U615 ( .A(G141GAT), .B(n551), .Z(n552) );
  XNOR2_X1 U616 ( .A(KEYINPUT114), .B(n552), .ZN(G1344GAT) );
  NOR2_X1 U617 ( .A1(n499), .A2(n559), .ZN(n557) );
  XOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n554) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(n555), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(G1345GAT) );
  NOR2_X1 U623 ( .A1(n584), .A2(n559), .ZN(n558) );
  XOR2_X1 U624 ( .A(G155GAT), .B(n558), .Z(G1346GAT) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U626 ( .A(G162GAT), .B(n561), .Z(G1347GAT) );
  XNOR2_X1 U627 ( .A(G169GAT), .B(KEYINPUT120), .ZN(n564) );
  NAND2_X1 U628 ( .A1(n562), .A2(n570), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n570), .A2(n565), .ZN(n567) );
  XOR2_X1 U631 ( .A(G176GAT), .B(KEYINPUT57), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n569) );
  XOR2_X1 U633 ( .A(KEYINPUT121), .B(KEYINPUT56), .Z(n568) );
  XNOR2_X1 U634 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n572) );
  NAND2_X1 U636 ( .A1(n402), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT124), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n579) );
  NAND2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n589) );
  NOR2_X1 U642 ( .A1(n577), .A2(n589), .ZN(n578) );
  XOR2_X1 U643 ( .A(n579), .B(n578), .Z(G1352GAT) );
  INV_X1 U644 ( .A(n580), .ZN(n581) );
  NOR2_X1 U645 ( .A1(n581), .A2(n589), .ZN(n583) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(G1353GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n589), .ZN(n586) );
  XNOR2_X1 U649 ( .A(G211GAT), .B(KEYINPUT125), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1354GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(KEYINPUT126), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(KEYINPUT127), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n591) );
  NOR2_X1 U654 ( .A1(n482), .A2(n589), .ZN(n590) );
  XOR2_X1 U655 ( .A(n591), .B(n590), .Z(G1355GAT) );
endmodule

