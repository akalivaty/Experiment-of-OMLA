

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754;

  XNOR2_X1 U381 ( .A(n409), .B(n408), .ZN(n495) );
  XNOR2_X1 U382 ( .A(n495), .B(n494), .ZN(n733) );
  OR2_X2 U383 ( .A1(n370), .A2(n507), .ZN(n509) );
  NOR2_X2 U384 ( .A1(n617), .A2(n620), .ZN(n619) );
  XNOR2_X2 U385 ( .A(n579), .B(KEYINPUT33), .ZN(n693) );
  NOR2_X2 U386 ( .A1(G902), .A2(n647), .ZN(n436) );
  INV_X2 U387 ( .A(G953), .ZN(n744) );
  NOR2_X1 U388 ( .A1(n501), .A2(n684), .ZN(n385) );
  OR2_X2 U389 ( .A1(n696), .A2(n695), .ZN(n600) );
  XNOR2_X1 U390 ( .A(n475), .B(n417), .ZN(n739) );
  INV_X1 U391 ( .A(G143), .ZN(n414) );
  AND2_X1 U392 ( .A1(n594), .A2(n591), .ZN(n592) );
  XNOR2_X1 U393 ( .A(n385), .B(KEYINPUT93), .ZN(n560) );
  XNOR2_X1 U394 ( .A(n456), .B(n455), .ZN(n575) );
  XNOR2_X1 U395 ( .A(n486), .B(n485), .ZN(n490) );
  XNOR2_X1 U396 ( .A(n673), .B(n739), .ZN(n432) );
  XNOR2_X1 U397 ( .A(n368), .B(n731), .ZN(n491) );
  XNOR2_X1 U398 ( .A(n429), .B(KEYINPUT74), .ZN(n368) );
  XNOR2_X1 U399 ( .A(n404), .B(G119), .ZN(n406) );
  XNOR2_X1 U400 ( .A(n367), .B(G110), .ZN(n731) );
  XNOR2_X1 U401 ( .A(n414), .B(G128), .ZN(n488) );
  INV_X1 U402 ( .A(KEYINPUT66), .ZN(n369) );
  INV_X1 U403 ( .A(KEYINPUT3), .ZN(n404) );
  XNOR2_X1 U404 ( .A(G107), .B(G104), .ZN(n367) );
  INV_X1 U405 ( .A(KEYINPUT109), .ZN(n360) );
  INV_X1 U406 ( .A(n525), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n499), .B(n498), .ZN(n501) );
  XOR2_X1 U408 ( .A(n360), .B(n361), .Z(n751) );
  NAND2_X1 U409 ( .A1(n527), .A2(n390), .ZN(n361) );
  XNOR2_X2 U410 ( .A(n369), .B(G101), .ZN(n429) );
  NOR2_X1 U411 ( .A1(n608), .A2(n383), .ZN(n540) );
  XNOR2_X1 U412 ( .A(n520), .B(n384), .ZN(n383) );
  INV_X1 U413 ( .A(KEYINPUT69), .ZN(n384) );
  NOR2_X1 U414 ( .A1(G953), .A2(KEYINPUT4), .ZN(n387) );
  NAND2_X1 U415 ( .A1(n386), .A2(KEYINPUT4), .ZN(n389) );
  XNOR2_X1 U416 ( .A(KEYINPUT72), .B(KEYINPUT73), .ZN(n405) );
  XNOR2_X1 U417 ( .A(n740), .B(n463), .ZN(n464) );
  XNOR2_X1 U418 ( .A(n380), .B(KEYINPUT88), .ZN(n402) );
  NOR2_X1 U419 ( .A1(n506), .A2(n364), .ZN(n380) );
  NAND2_X1 U420 ( .A1(n603), .A2(n540), .ZN(n382) );
  NOR2_X1 U421 ( .A1(n713), .A2(G953), .ZN(n506) );
  XNOR2_X1 U422 ( .A(n534), .B(KEYINPUT39), .ZN(n571) );
  XNOR2_X1 U423 ( .A(n560), .B(n502), .ZN(n370) );
  BUF_X1 U424 ( .A(n515), .Z(n698) );
  XNOR2_X1 U425 ( .A(n434), .B(n433), .ZN(n435) );
  NAND2_X1 U426 ( .A1(n379), .A2(KEYINPUT47), .ZN(n378) );
  NAND2_X1 U427 ( .A1(n552), .A2(n672), .ZN(n379) );
  AND2_X1 U428 ( .A1(n549), .A2(n551), .ZN(n377) );
  XOR2_X1 U429 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n485) );
  NAND2_X1 U430 ( .A1(n389), .A2(n388), .ZN(n486) );
  NAND2_X1 U431 ( .A1(n387), .A2(G224), .ZN(n388) );
  NOR2_X1 U432 ( .A1(n754), .A2(n753), .ZN(n544) );
  XNOR2_X1 U433 ( .A(n374), .B(n398), .ZN(n400) );
  XNOR2_X1 U434 ( .A(n375), .B(KEYINPUT14), .ZN(n374) );
  INV_X1 U435 ( .A(KEYINPUT81), .ZN(n375) );
  XNOR2_X1 U436 ( .A(G116), .B(G113), .ZN(n407) );
  XNOR2_X1 U437 ( .A(n469), .B(n468), .ZN(n639) );
  XNOR2_X1 U438 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U439 ( .A(n616), .B(n615), .ZN(n620) );
  INV_X1 U440 ( .A(n621), .ZN(n373) );
  XNOR2_X1 U441 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n538) );
  AND2_X1 U442 ( .A1(n458), .A2(n457), .ZN(n533) );
  XNOR2_X1 U443 ( .A(n382), .B(n381), .ZN(n542) );
  INV_X1 U444 ( .A(KEYINPUT28), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n634), .B(n633), .ZN(n720) );
  NOR2_X1 U446 ( .A1(n577), .A2(n609), .ZN(n390) );
  NOR2_X1 U447 ( .A1(n698), .A2(n600), .ZN(n362) );
  AND2_X1 U448 ( .A1(n625), .A2(n624), .ZN(n363) );
  AND2_X1 U449 ( .A1(G953), .A2(n401), .ZN(n364) );
  AND2_X1 U450 ( .A1(n378), .A2(n376), .ZN(n365) );
  XOR2_X1 U451 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n366) );
  INV_X1 U452 ( .A(G146), .ZN(n673) );
  NOR2_X1 U453 ( .A1(n547), .A2(n370), .ZN(n672) );
  AND2_X2 U454 ( .A1(n371), .A2(n625), .ZN(n721) );
  AND2_X1 U455 ( .A1(n624), .A2(n372), .ZN(n371) );
  INV_X1 U456 ( .A(n626), .ZN(n372) );
  AND2_X2 U457 ( .A1(n527), .A2(n391), .ZN(n530) );
  NAND2_X1 U458 ( .A1(n574), .A2(n373), .ZN(n622) );
  XNOR2_X1 U459 ( .A(n570), .B(n366), .ZN(n574) );
  NAND2_X1 U460 ( .A1(n400), .A2(G952), .ZN(n399) );
  NAND2_X1 U461 ( .A1(n672), .A2(n377), .ZN(n376) );
  INV_X1 U462 ( .A(n501), .ZN(n525) );
  NAND2_X1 U463 ( .A1(n744), .A2(G224), .ZN(n386) );
  NOR2_X1 U464 ( .A1(n528), .A2(n577), .ZN(n391) );
  XNOR2_X2 U465 ( .A(n530), .B(n529), .ZN(n590) );
  XNOR2_X1 U466 ( .A(n410), .B(n495), .ZN(n413) );
  XOR2_X1 U467 ( .A(n412), .B(n411), .Z(n392) );
  NOR2_X1 U468 ( .A1(n510), .A2(n548), .ZN(n393) );
  NOR2_X1 U469 ( .A1(n621), .A2(n573), .ZN(n394) );
  INV_X1 U470 ( .A(KEYINPUT110), .ZN(n576) );
  XNOR2_X1 U471 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U472 ( .A(n452), .B(KEYINPUT84), .ZN(n453) );
  XNOR2_X1 U473 ( .A(n413), .B(n392), .ZN(n418) );
  XNOR2_X1 U474 ( .A(G140), .B(KEYINPUT10), .ZN(n439) );
  INV_X1 U475 ( .A(G134), .ZN(n415) );
  INV_X1 U476 ( .A(KEYINPUT2), .ZN(n618) );
  INV_X1 U477 ( .A(KEYINPUT30), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U479 ( .A(n488), .B(n415), .ZN(n475) );
  XNOR2_X1 U480 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n446), .B(n445), .ZN(n447) );
  NOR2_X1 U482 ( .A1(n606), .A2(n575), .ZN(n457) );
  XNOR2_X1 U483 ( .A(n539), .B(n538), .ZN(n706) );
  INV_X1 U484 ( .A(KEYINPUT32), .ZN(n529) );
  XNOR2_X1 U485 ( .A(KEYINPUT15), .B(G902), .ZN(n626) );
  NAND2_X1 U486 ( .A1(G234), .A2(n626), .ZN(n395) );
  XNOR2_X1 U487 ( .A(KEYINPUT20), .B(n395), .ZN(n451) );
  AND2_X1 U488 ( .A1(n451), .A2(G221), .ZN(n397) );
  INV_X1 U489 ( .A(KEYINPUT21), .ZN(n396) );
  XNOR2_X1 U490 ( .A(n397), .B(n396), .ZN(n700) );
  NAND2_X1 U491 ( .A1(G237), .A2(G234), .ZN(n398) );
  XNOR2_X1 U492 ( .A(n399), .B(KEYINPUT98), .ZN(n713) );
  NAND2_X1 U493 ( .A1(G902), .A2(n400), .ZN(n504) );
  NOR2_X1 U494 ( .A1(G900), .A2(n504), .ZN(n401) );
  OR2_X1 U495 ( .A1(n700), .A2(n402), .ZN(n520) );
  NOR2_X1 U496 ( .A1(G953), .A2(G237), .ZN(n403) );
  XOR2_X1 U497 ( .A(KEYINPUT83), .B(n403), .Z(n465) );
  NAND2_X1 U498 ( .A1(n465), .A2(G210), .ZN(n410) );
  XNOR2_X1 U499 ( .A(n406), .B(n405), .ZN(n409) );
  XNOR2_X1 U500 ( .A(n407), .B(KEYINPUT96), .ZN(n408) );
  XOR2_X1 U501 ( .A(KEYINPUT82), .B(KEYINPUT5), .Z(n412) );
  XNOR2_X1 U502 ( .A(n429), .B(KEYINPUT104), .ZN(n411) );
  XOR2_X1 U503 ( .A(G131), .B(KEYINPUT4), .Z(n416) );
  XNOR2_X1 U504 ( .A(G137), .B(n416), .ZN(n417) );
  XNOR2_X1 U505 ( .A(n418), .B(n432), .ZN(n653) );
  INV_X1 U506 ( .A(G902), .ZN(n482) );
  NAND2_X1 U507 ( .A1(n653), .A2(n482), .ZN(n421) );
  INV_X1 U508 ( .A(KEYINPUT76), .ZN(n419) );
  XNOR2_X1 U509 ( .A(n419), .B(G472), .ZN(n420) );
  XNOR2_X1 U510 ( .A(n421), .B(n420), .ZN(n515) );
  INV_X1 U511 ( .A(G237), .ZN(n422) );
  NAND2_X1 U512 ( .A1(n482), .A2(n422), .ZN(n497) );
  NAND2_X1 U513 ( .A1(n497), .A2(G214), .ZN(n423) );
  XNOR2_X1 U514 ( .A(n423), .B(KEYINPUT97), .ZN(n684) );
  NOR2_X1 U515 ( .A1(n515), .A2(n684), .ZN(n425) );
  NOR2_X1 U516 ( .A1(n520), .A2(n426), .ZN(n458) );
  XOR2_X1 U517 ( .A(G140), .B(KEYINPUT86), .Z(n428) );
  NAND2_X1 U518 ( .A1(G227), .A2(n744), .ZN(n427) );
  XNOR2_X1 U519 ( .A(n428), .B(n427), .ZN(n430) );
  XOR2_X1 U520 ( .A(n430), .B(n491), .Z(n431) );
  XNOR2_X1 U521 ( .A(n432), .B(n431), .ZN(n647) );
  XNOR2_X1 U522 ( .A(KEYINPUT71), .B(KEYINPUT70), .ZN(n434) );
  INV_X1 U523 ( .A(G469), .ZN(n433) );
  XNOR2_X2 U524 ( .A(n436), .B(n435), .ZN(n606) );
  NAND2_X1 U525 ( .A1(n744), .A2(G234), .ZN(n438) );
  XNOR2_X1 U526 ( .A(KEYINPUT67), .B(KEYINPUT8), .ZN(n437) );
  XNOR2_X1 U527 ( .A(n438), .B(n437), .ZN(n476) );
  NAND2_X1 U528 ( .A1(n476), .A2(G221), .ZN(n450) );
  XOR2_X2 U529 ( .A(G146), .B(G125), .Z(n487) );
  XNOR2_X2 U530 ( .A(n487), .B(n439), .ZN(n740) );
  XOR2_X1 U531 ( .A(KEYINPUT85), .B(KEYINPUT23), .Z(n441) );
  XNOR2_X1 U532 ( .A(KEYINPUT102), .B(KEYINPUT24), .ZN(n440) );
  XNOR2_X1 U533 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U534 ( .A(n740), .B(n442), .ZN(n448) );
  XOR2_X1 U535 ( .A(G119), .B(G137), .Z(n444) );
  XNOR2_X1 U536 ( .A(G128), .B(G110), .ZN(n443) );
  XNOR2_X1 U537 ( .A(n444), .B(n443), .ZN(n446) );
  XOR2_X1 U538 ( .A(KEYINPUT101), .B(KEYINPUT100), .Z(n445) );
  XNOR2_X1 U539 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U540 ( .A(n450), .B(n449), .ZN(n722) );
  NOR2_X1 U541 ( .A1(G902), .A2(n722), .ZN(n456) );
  NAND2_X1 U542 ( .A1(n451), .A2(G217), .ZN(n454) );
  XNOR2_X1 U543 ( .A(KEYINPUT103), .B(KEYINPUT25), .ZN(n452) );
  INV_X1 U544 ( .A(n575), .ZN(n608) );
  XOR2_X1 U545 ( .A(KEYINPUT107), .B(G104), .Z(n460) );
  XNOR2_X1 U546 ( .A(G143), .B(G122), .ZN(n459) );
  XNOR2_X1 U547 ( .A(n460), .B(n459), .ZN(n462) );
  XOR2_X1 U548 ( .A(KEYINPUT11), .B(KEYINPUT106), .Z(n461) );
  XNOR2_X1 U549 ( .A(n464), .B(KEYINPUT12), .ZN(n469) );
  AND2_X1 U550 ( .A1(G214), .A2(n465), .ZN(n467) );
  XOR2_X1 U551 ( .A(G131), .B(G113), .Z(n466) );
  NAND2_X1 U552 ( .A1(n639), .A2(n482), .ZN(n471) );
  XOR2_X1 U553 ( .A(KEYINPUT13), .B(G475), .Z(n470) );
  XNOR2_X1 U554 ( .A(n471), .B(n470), .ZN(n510) );
  XOR2_X1 U555 ( .A(KEYINPUT7), .B(G107), .Z(n473) );
  XNOR2_X1 U556 ( .A(G116), .B(G122), .ZN(n472) );
  XNOR2_X1 U557 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U558 ( .A(n475), .B(n474), .Z(n481) );
  NAND2_X1 U559 ( .A1(G217), .A2(n476), .ZN(n479) );
  INV_X1 U560 ( .A(KEYINPUT108), .ZN(n477) );
  XNOR2_X1 U561 ( .A(n477), .B(KEYINPUT9), .ZN(n478) );
  XNOR2_X1 U562 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U563 ( .A(n481), .B(n480), .ZN(n658) );
  NAND2_X1 U564 ( .A1(n658), .A2(n482), .ZN(n483) );
  XNOR2_X1 U565 ( .A(n483), .B(G478), .ZN(n519) );
  NAND2_X1 U566 ( .A1(n510), .A2(n519), .ZN(n484) );
  XNOR2_X1 U567 ( .A(KEYINPUT111), .B(n484), .ZN(n583) );
  NAND2_X1 U568 ( .A1(n533), .A2(n583), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U570 ( .A(n490), .B(n489), .ZN(n492) );
  XNOR2_X1 U571 ( .A(n492), .B(n491), .ZN(n496) );
  XNOR2_X1 U572 ( .A(KEYINPUT16), .B(G122), .ZN(n493) );
  XNOR2_X1 U573 ( .A(n493), .B(KEYINPUT79), .ZN(n494) );
  XNOR2_X1 U574 ( .A(n496), .B(n733), .ZN(n627) );
  NAND2_X1 U575 ( .A1(n627), .A2(n626), .ZN(n499) );
  NAND2_X1 U576 ( .A1(n497), .A2(G210), .ZN(n498) );
  NOR2_X1 U577 ( .A1(n500), .A2(n359), .ZN(n546) );
  XOR2_X1 U578 ( .A(G143), .B(n546), .Z(G45) );
  XNOR2_X1 U579 ( .A(KEYINPUT65), .B(KEYINPUT19), .ZN(n502) );
  NOR2_X1 U580 ( .A1(G898), .A2(n744), .ZN(n503) );
  XNOR2_X1 U581 ( .A(KEYINPUT99), .B(n503), .ZN(n734) );
  NOR2_X1 U582 ( .A1(n504), .A2(n734), .ZN(n505) );
  NOR2_X1 U583 ( .A1(n506), .A2(n505), .ZN(n507) );
  INV_X1 U584 ( .A(KEYINPUT0), .ZN(n508) );
  XNOR2_X2 U585 ( .A(n509), .B(n508), .ZN(n580) );
  OR2_X1 U586 ( .A1(n510), .A2(n519), .ZN(n537) );
  NOR2_X1 U587 ( .A1(n537), .A2(n700), .ZN(n511) );
  NAND2_X1 U588 ( .A1(n580), .A2(n511), .ZN(n514) );
  XNOR2_X1 U589 ( .A(KEYINPUT78), .B(KEYINPUT22), .ZN(n512) );
  XNOR2_X1 U590 ( .A(n512), .B(KEYINPUT77), .ZN(n513) );
  XNOR2_X2 U591 ( .A(n514), .B(n513), .ZN(n527) );
  XNOR2_X2 U592 ( .A(n606), .B(KEYINPUT1), .ZN(n696) );
  INV_X1 U593 ( .A(n696), .ZN(n564) );
  NAND2_X1 U594 ( .A1(n698), .A2(n575), .ZN(n516) );
  NOR2_X1 U595 ( .A1(n564), .A2(n516), .ZN(n517) );
  NAND2_X1 U596 ( .A1(n527), .A2(n517), .ZN(n589) );
  XNOR2_X1 U597 ( .A(G110), .B(KEYINPUT116), .ZN(n518) );
  XNOR2_X1 U598 ( .A(n589), .B(n518), .ZN(G12) );
  INV_X1 U599 ( .A(n519), .ZN(n548) );
  AND2_X1 U600 ( .A1(n510), .A2(n548), .ZN(n675) );
  INV_X1 U601 ( .A(n675), .ZN(n522) );
  XNOR2_X1 U602 ( .A(n698), .B(KEYINPUT6), .ZN(n577) );
  NAND2_X1 U603 ( .A1(n540), .A2(n577), .ZN(n521) );
  NOR2_X1 U604 ( .A1(n522), .A2(n521), .ZN(n562) );
  NAND2_X1 U605 ( .A1(n562), .A2(n696), .ZN(n523) );
  NOR2_X1 U606 ( .A1(n684), .A2(n523), .ZN(n524) );
  XNOR2_X1 U607 ( .A(n524), .B(KEYINPUT43), .ZN(n526) );
  OR2_X1 U608 ( .A1(n526), .A2(n525), .ZN(n572) );
  XNOR2_X1 U609 ( .A(n572), .B(G140), .ZN(G42) );
  NAND2_X1 U610 ( .A1(n564), .A2(n575), .ZN(n528) );
  XNOR2_X1 U611 ( .A(n590), .B(G119), .ZN(G21) );
  INV_X1 U612 ( .A(KEYINPUT38), .ZN(n531) );
  XNOR2_X1 U613 ( .A(n359), .B(n531), .ZN(n685) );
  INV_X1 U614 ( .A(n685), .ZN(n532) );
  NAND2_X1 U615 ( .A1(n533), .A2(n532), .ZN(n534) );
  NAND2_X1 U616 ( .A1(n571), .A2(n675), .ZN(n535) );
  XOR2_X1 U617 ( .A(n535), .B(KEYINPUT40), .Z(n754) );
  NOR2_X1 U618 ( .A1(n685), .A2(n684), .ZN(n536) );
  XNOR2_X1 U619 ( .A(n536), .B(KEYINPUT112), .ZN(n690) );
  INV_X1 U620 ( .A(n537), .ZN(n687) );
  NAND2_X1 U621 ( .A1(n690), .A2(n687), .ZN(n539) );
  INV_X1 U622 ( .A(n698), .ZN(n603) );
  INV_X1 U623 ( .A(n606), .ZN(n541) );
  NAND2_X1 U624 ( .A1(n542), .A2(n541), .ZN(n547) );
  NOR2_X1 U625 ( .A1(n706), .A2(n547), .ZN(n543) );
  XNOR2_X1 U626 ( .A(n543), .B(KEYINPUT42), .ZN(n753) );
  XNOR2_X1 U627 ( .A(KEYINPUT46), .B(n544), .ZN(n556) );
  INV_X1 U628 ( .A(KEYINPUT47), .ZN(n553) );
  AND2_X1 U629 ( .A1(n553), .A2(KEYINPUT89), .ZN(n545) );
  NOR2_X1 U630 ( .A1(n546), .A2(n545), .ZN(n554) );
  INV_X1 U631 ( .A(KEYINPUT80), .ZN(n551) );
  NOR2_X1 U632 ( .A1(n675), .A2(n393), .ZN(n549) );
  INV_X1 U633 ( .A(n549), .ZN(n689) );
  NOR2_X1 U634 ( .A1(KEYINPUT89), .A2(n689), .ZN(n550) );
  NOR2_X1 U635 ( .A1(n551), .A2(n550), .ZN(n552) );
  AND2_X1 U636 ( .A1(n554), .A2(n365), .ZN(n555) );
  AND2_X1 U637 ( .A1(n556), .A2(n555), .ZN(n569) );
  NAND2_X1 U638 ( .A1(n672), .A2(KEYINPUT80), .ZN(n557) );
  NOR2_X1 U639 ( .A1(n557), .A2(KEYINPUT47), .ZN(n558) );
  NOR2_X1 U640 ( .A1(KEYINPUT89), .A2(n558), .ZN(n559) );
  NOR2_X1 U641 ( .A1(n549), .A2(n559), .ZN(n567) );
  INV_X1 U642 ( .A(n560), .ZN(n561) );
  NAND2_X1 U643 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U644 ( .A(KEYINPUT36), .B(n563), .Z(n565) );
  NAND2_X1 U645 ( .A1(n565), .A2(n564), .ZN(n680) );
  XNOR2_X1 U646 ( .A(KEYINPUT91), .B(n680), .ZN(n566) );
  NOR2_X1 U647 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U648 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n571), .A2(n393), .ZN(n683) );
  NAND2_X1 U650 ( .A1(n683), .A2(n572), .ZN(n621) );
  INV_X1 U651 ( .A(KEYINPUT90), .ZN(n573) );
  NAND2_X1 U652 ( .A1(n574), .A2(n394), .ZN(n617) );
  OR2_X1 U653 ( .A1(n700), .A2(n575), .ZN(n695) );
  XNOR2_X1 U654 ( .A(n600), .B(n576), .ZN(n578) );
  NAND2_X1 U655 ( .A1(n578), .A2(n577), .ZN(n579) );
  NAND2_X1 U656 ( .A1(n693), .A2(n580), .ZN(n582) );
  XNOR2_X1 U657 ( .A(KEYINPUT75), .B(KEYINPUT34), .ZN(n581) );
  XNOR2_X1 U658 ( .A(n582), .B(n581), .ZN(n585) );
  XOR2_X1 U659 ( .A(n583), .B(KEYINPUT87), .Z(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n587) );
  INV_X1 U661 ( .A(KEYINPUT35), .ZN(n586) );
  XNOR2_X2 U662 ( .A(n587), .B(n586), .ZN(n752) );
  INV_X1 U663 ( .A(KEYINPUT92), .ZN(n588) );
  NAND2_X1 U664 ( .A1(n752), .A2(n588), .ZN(n593) );
  NAND2_X1 U665 ( .A1(n590), .A2(n589), .ZN(n594) );
  INV_X1 U666 ( .A(KEYINPUT44), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n593), .ZN(n599) );
  INV_X1 U668 ( .A(n594), .ZN(n597) );
  NOR2_X1 U669 ( .A1(n588), .A2(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n752), .A2(n595), .ZN(n596) );
  NAND2_X1 U671 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U672 ( .A1(n599), .A2(n598), .ZN(n614) );
  OR2_X1 U673 ( .A1(n752), .A2(n591), .ZN(n612) );
  NAND2_X1 U674 ( .A1(n580), .A2(n362), .ZN(n602) );
  XOR2_X1 U675 ( .A(KEYINPUT31), .B(KEYINPUT105), .Z(n601) );
  XNOR2_X1 U676 ( .A(n602), .B(n601), .ZN(n678) );
  NOR2_X1 U677 ( .A1(n603), .A2(n695), .ZN(n604) );
  NAND2_X1 U678 ( .A1(n604), .A2(n580), .ZN(n605) );
  NOR2_X1 U679 ( .A1(n606), .A2(n605), .ZN(n664) );
  NOR2_X1 U680 ( .A1(n678), .A2(n664), .ZN(n607) );
  NOR2_X1 U681 ( .A1(n607), .A2(n549), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n696), .A2(n608), .ZN(n609) );
  NOR2_X1 U683 ( .A1(n610), .A2(n751), .ZN(n611) );
  AND2_X1 U684 ( .A1(n612), .A2(n611), .ZN(n613) );
  NAND2_X1 U685 ( .A1(n614), .A2(n613), .ZN(n616) );
  XOR2_X1 U686 ( .A(KEYINPUT64), .B(KEYINPUT45), .Z(n615) );
  XNOR2_X1 U687 ( .A(n619), .B(n618), .ZN(n625) );
  INV_X1 U688 ( .A(n620), .ZN(n726) );
  INV_X1 U689 ( .A(n622), .ZN(n738) );
  NOR2_X1 U690 ( .A1(n738), .A2(KEYINPUT90), .ZN(n623) );
  NAND2_X1 U691 ( .A1(n726), .A2(n623), .ZN(n624) );
  NAND2_X1 U692 ( .A1(n721), .A2(G210), .ZN(n631) );
  XNOR2_X1 U693 ( .A(KEYINPUT122), .B(KEYINPUT54), .ZN(n628) );
  XOR2_X1 U694 ( .A(n628), .B(KEYINPUT55), .Z(n629) );
  XNOR2_X1 U695 ( .A(n627), .B(n629), .ZN(n630) );
  XNOR2_X1 U696 ( .A(n631), .B(n630), .ZN(n635) );
  INV_X1 U697 ( .A(G952), .ZN(n632) );
  NAND2_X1 U698 ( .A1(n632), .A2(G953), .ZN(n634) );
  INV_X1 U699 ( .A(KEYINPUT95), .ZN(n633) );
  NAND2_X1 U700 ( .A1(n635), .A2(n720), .ZN(n637) );
  INV_X1 U701 ( .A(KEYINPUT56), .ZN(n636) );
  XNOR2_X1 U702 ( .A(n637), .B(n636), .ZN(G51) );
  NAND2_X1 U703 ( .A1(n721), .A2(G475), .ZN(n641) );
  XOR2_X1 U704 ( .A(KEYINPUT94), .B(KEYINPUT59), .Z(n638) );
  XNOR2_X1 U705 ( .A(n639), .B(n638), .ZN(n640) );
  XNOR2_X1 U706 ( .A(n641), .B(n640), .ZN(n642) );
  NAND2_X1 U707 ( .A1(n642), .A2(n720), .ZN(n644) );
  INV_X1 U708 ( .A(KEYINPUT60), .ZN(n643) );
  XNOR2_X1 U709 ( .A(n644), .B(n643), .ZN(G60) );
  NAND2_X1 U710 ( .A1(n721), .A2(G469), .ZN(n649) );
  XNOR2_X1 U711 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n645) );
  XOR2_X1 U712 ( .A(n645), .B(KEYINPUT58), .Z(n646) );
  XNOR2_X1 U713 ( .A(n647), .B(n646), .ZN(n648) );
  XNOR2_X1 U714 ( .A(n649), .B(n648), .ZN(n650) );
  NAND2_X1 U715 ( .A1(n650), .A2(n720), .ZN(n652) );
  INV_X1 U716 ( .A(KEYINPUT124), .ZN(n651) );
  XNOR2_X1 U717 ( .A(n652), .B(n651), .ZN(G54) );
  NAND2_X1 U718 ( .A1(n721), .A2(G472), .ZN(n655) );
  XNOR2_X1 U719 ( .A(n653), .B(KEYINPUT62), .ZN(n654) );
  XNOR2_X1 U720 ( .A(n655), .B(n654), .ZN(n656) );
  NAND2_X1 U721 ( .A1(n656), .A2(n720), .ZN(n657) );
  XNOR2_X1 U722 ( .A(n657), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U723 ( .A1(n721), .A2(G478), .ZN(n659) );
  XNOR2_X1 U724 ( .A(n659), .B(n658), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n660), .A2(n720), .ZN(n661) );
  XNOR2_X1 U726 ( .A(n661), .B(KEYINPUT125), .ZN(G63) );
  NAND2_X1 U727 ( .A1(n664), .A2(n675), .ZN(n662) );
  XNOR2_X1 U728 ( .A(n662), .B(KEYINPUT114), .ZN(n663) );
  XNOR2_X1 U729 ( .A(G104), .B(n663), .ZN(G6) );
  XOR2_X1 U730 ( .A(KEYINPUT115), .B(KEYINPUT26), .Z(n666) );
  NAND2_X1 U731 ( .A1(n664), .A2(n393), .ZN(n665) );
  XNOR2_X1 U732 ( .A(n666), .B(n665), .ZN(n668) );
  XOR2_X1 U733 ( .A(G107), .B(KEYINPUT27), .Z(n667) );
  XNOR2_X1 U734 ( .A(n668), .B(n667), .ZN(G9) );
  XOR2_X1 U735 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n670) );
  NAND2_X1 U736 ( .A1(n672), .A2(n393), .ZN(n669) );
  XNOR2_X1 U737 ( .A(n670), .B(n669), .ZN(n671) );
  XOR2_X1 U738 ( .A(G128), .B(n671), .Z(G30) );
  NAND2_X1 U739 ( .A1(n672), .A2(n675), .ZN(n674) );
  XNOR2_X1 U740 ( .A(n674), .B(G146), .ZN(G48) );
  NAND2_X1 U741 ( .A1(n678), .A2(n675), .ZN(n676) );
  XNOR2_X1 U742 ( .A(n676), .B(KEYINPUT118), .ZN(n677) );
  XNOR2_X1 U743 ( .A(G113), .B(n677), .ZN(G15) );
  NAND2_X1 U744 ( .A1(n678), .A2(n393), .ZN(n679) );
  XNOR2_X1 U745 ( .A(n679), .B(G116), .ZN(G18) );
  XNOR2_X1 U746 ( .A(KEYINPUT119), .B(KEYINPUT37), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U748 ( .A(G125), .B(n682), .ZN(G27) );
  XNOR2_X1 U749 ( .A(G134), .B(n683), .ZN(G36) );
  NAND2_X1 U750 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U751 ( .A(KEYINPUT120), .B(n686), .ZN(n688) );
  NAND2_X1 U752 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U753 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U754 ( .A1(n692), .A2(n691), .ZN(n694) );
  NAND2_X1 U755 ( .A1(n694), .A2(n693), .ZN(n709) );
  NAND2_X1 U756 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U757 ( .A(KEYINPUT50), .B(n697), .ZN(n699) );
  NAND2_X1 U758 ( .A1(n699), .A2(n698), .ZN(n703) );
  NAND2_X1 U759 ( .A1(n700), .A2(n575), .ZN(n701) );
  XNOR2_X1 U760 ( .A(KEYINPUT49), .B(n701), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U762 ( .A1(n362), .A2(n704), .ZN(n705) );
  XNOR2_X1 U763 ( .A(KEYINPUT51), .B(n705), .ZN(n707) );
  INV_X1 U764 ( .A(n706), .ZN(n714) );
  NAND2_X1 U765 ( .A1(n707), .A2(n714), .ZN(n708) );
  NAND2_X1 U766 ( .A1(n709), .A2(n708), .ZN(n710) );
  XNOR2_X1 U767 ( .A(n710), .B(KEYINPUT52), .ZN(n711) );
  XNOR2_X1 U768 ( .A(n711), .B(KEYINPUT121), .ZN(n712) );
  NOR2_X1 U769 ( .A1(n713), .A2(n712), .ZN(n716) );
  AND2_X1 U770 ( .A1(n693), .A2(n714), .ZN(n715) );
  NOR2_X1 U771 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U772 ( .A1(n717), .A2(n744), .ZN(n718) );
  NOR2_X1 U773 ( .A1(n363), .A2(n718), .ZN(n719) );
  XNOR2_X1 U774 ( .A(n719), .B(KEYINPUT53), .ZN(G75) );
  INV_X1 U775 ( .A(n720), .ZN(n725) );
  NAND2_X1 U776 ( .A1(n721), .A2(G217), .ZN(n723) );
  XNOR2_X1 U777 ( .A(n723), .B(n722), .ZN(n724) );
  NOR2_X1 U778 ( .A1(n725), .A2(n724), .ZN(G66) );
  NAND2_X1 U779 ( .A1(n726), .A2(n744), .ZN(n730) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U781 ( .A(KEYINPUT61), .B(n727), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n728), .A2(G898), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n737) );
  XNOR2_X1 U784 ( .A(n731), .B(G101), .ZN(n732) );
  XNOR2_X1 U785 ( .A(n733), .B(n732), .ZN(n735) );
  NAND2_X1 U786 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U787 ( .A(n737), .B(n736), .Z(G69) );
  XNOR2_X1 U788 ( .A(KEYINPUT127), .B(n622), .ZN(n743) );
  XOR2_X1 U789 ( .A(n739), .B(n740), .Z(n741) );
  XNOR2_X1 U790 ( .A(KEYINPUT126), .B(n741), .ZN(n746) );
  INV_X1 U791 ( .A(n746), .ZN(n742) );
  XNOR2_X1 U792 ( .A(n743), .B(n742), .ZN(n745) );
  NAND2_X1 U793 ( .A1(n745), .A2(n744), .ZN(n750) );
  XNOR2_X1 U794 ( .A(G227), .B(n746), .ZN(n747) );
  NAND2_X1 U795 ( .A1(n747), .A2(G900), .ZN(n748) );
  NAND2_X1 U796 ( .A1(n748), .A2(G953), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n750), .A2(n749), .ZN(G72) );
  XOR2_X1 U798 ( .A(G101), .B(n751), .Z(G3) );
  XNOR2_X1 U799 ( .A(n752), .B(G122), .ZN(G24) );
  XOR2_X1 U800 ( .A(G137), .B(n753), .Z(G39) );
  XOR2_X1 U801 ( .A(G131), .B(n754), .Z(G33) );
endmodule

