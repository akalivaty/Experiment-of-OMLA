//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:20 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n951, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(KEYINPUT31), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT11), .A3(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(G137), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n192), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT64), .ZN(new_n196));
  INV_X1    g010(.A(G131), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n192), .A3(new_n197), .A4(new_n193), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(KEYINPUT64), .A3(G131), .ZN(new_n200));
  INV_X1    g014(.A(G146), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G143), .ZN(new_n202));
  INV_X1    g016(.A(G143), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G146), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n202), .A2(new_n204), .A3(KEYINPUT0), .A4(G128), .ZN(new_n205));
  XNOR2_X1  g019(.A(G143), .B(G146), .ZN(new_n206));
  XNOR2_X1  g020(.A(KEYINPUT0), .B(G128), .ZN(new_n207));
  OAI21_X1  g021(.A(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n199), .A2(new_n200), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G116), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(KEYINPUT68), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g031(.A(G116), .B(G119), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT68), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT2), .ZN(new_n220));
  INV_X1    g034(.A(G113), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(KEYINPUT66), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT66), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n223), .B1(KEYINPUT2), .B2(G113), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT2), .A2(G113), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND3_X1  g042(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n217), .A2(new_n219), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n225), .A2(new_n230), .A3(new_n218), .ZN(new_n232));
  INV_X1    g046(.A(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n231), .A2(new_n233), .ZN(new_n234));
  OAI21_X1  g048(.A(KEYINPUT1), .B1(new_n203), .B2(G146), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G128), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n202), .A2(new_n204), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n206), .A2(G128), .A3(new_n235), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n193), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n189), .A2(G137), .ZN(new_n242));
  OAI21_X1  g056(.A(G131), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n198), .A3(new_n243), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n210), .A2(new_n234), .A3(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n210), .A2(new_n244), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT30), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(KEYINPUT65), .A2(KEYINPUT30), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n210), .A2(new_n247), .A3(new_n248), .A4(new_n244), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND3_X1   g069(.A1(new_n212), .A2(new_n214), .A3(KEYINPUT68), .ZN(new_n256));
  AOI21_X1  g070(.A(KEYINPUT68), .B1(new_n212), .B2(new_n214), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  AOI22_X1  g072(.A1(new_n224), .A2(new_n222), .B1(new_n228), .B2(new_n229), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n232), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n245), .B1(new_n255), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n187), .B1(new_n261), .B2(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n234), .B1(new_n253), .B2(new_n254), .ZN(new_n268));
  INV_X1    g082(.A(new_n266), .ZN(new_n269));
  NOR4_X1   g083(.A1(new_n268), .A2(KEYINPUT31), .A3(new_n245), .A4(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n266), .B(KEYINPUT69), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n234), .B1(new_n210), .B2(new_n244), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT28), .B1(new_n245), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n210), .A2(new_n234), .A3(new_n244), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n272), .B1(new_n274), .B2(new_n277), .ZN(new_n278));
  NOR3_X1   g092(.A1(new_n267), .A2(new_n270), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g093(.A1(G472), .A2(G902), .ZN(new_n280));
  INV_X1    g094(.A(new_n280), .ZN(new_n281));
  OAI21_X1  g095(.A(KEYINPUT70), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(new_n249), .B(new_n251), .C1(new_n210), .C2(new_n244), .ZN(new_n283));
  AND4_X1   g097(.A1(new_n247), .A2(new_n210), .A3(new_n248), .A4(new_n244), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n260), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n285), .A2(new_n275), .A3(new_n266), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(KEYINPUT31), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n274), .A2(new_n277), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n271), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n285), .A2(new_n187), .A3(new_n275), .A4(new_n266), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n287), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  AND3_X1   g105(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n280), .ZN(new_n292));
  AOI21_X1  g106(.A(KEYINPUT32), .B1(new_n291), .B2(new_n280), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n282), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n295), .B1(new_n274), .B2(new_n277), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n246), .A2(new_n260), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n275), .ZN(new_n298));
  AOI21_X1  g112(.A(KEYINPUT71), .B1(new_n298), .B2(KEYINPUT28), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT29), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n269), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT72), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n306), .A3(new_n302), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n301), .B1(new_n288), .B2(new_n271), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n266), .B1(new_n285), .B2(new_n275), .ZN(new_n309));
  OR2_X1    g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g124(.A1(new_n304), .A2(new_n305), .A3(new_n307), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G472), .ZN(new_n312));
  OAI211_X1 g126(.A(KEYINPUT70), .B(KEYINPUT32), .C1(new_n279), .C2(new_n281), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n294), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n305), .ZN(new_n316));
  INV_X1    g130(.A(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G128), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n318), .A2(KEYINPUT23), .A3(G119), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT73), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(KEYINPUT23), .B1(new_n318), .B2(G119), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT74), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n211), .A2(G128), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n326), .A2(KEYINPUT74), .A3(KEYINPUT23), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n324), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n321), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n326), .ZN(new_n331));
  XNOR2_X1  g145(.A(KEYINPUT24), .B(G110), .ZN(new_n332));
  OR2_X1    g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(G125), .B(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT16), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT16), .ZN(new_n336));
  INV_X1    g150(.A(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n336), .A2(new_n337), .A3(G125), .ZN(new_n338));
  AOI21_X1  g152(.A(G146), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n335), .A2(G146), .A3(new_n338), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n330), .B(new_n333), .C1(new_n339), .C2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(G110), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n328), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n331), .A2(new_n332), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n334), .A2(new_n201), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n346), .A2(new_n340), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n342), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT22), .B(G137), .ZN(new_n350));
  INV_X1    g164(.A(G953), .ZN(new_n351));
  AND3_X1   g165(.A1(new_n351), .A2(G221), .A3(G234), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n350), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n342), .A2(new_n348), .A3(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n305), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT25), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n354), .A2(KEYINPUT25), .A3(new_n356), .A4(new_n305), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n317), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n356), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n355), .B1(new_n342), .B2(new_n348), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n362), .A2(KEYINPUT75), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT75), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n365), .B1(new_n354), .B2(new_n356), .ZN(new_n366));
  NOR2_X1   g180(.A1(new_n316), .A2(G902), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n364), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n361), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  INV_X1    g185(.A(G237), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(new_n351), .A3(G214), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(new_n203), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n371), .B1(new_n376), .B2(G131), .ZN(new_n377));
  AOI211_X1 g191(.A(KEYINPUT85), .B(new_n197), .C1(new_n374), .C2(new_n375), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT17), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  AND4_X1   g193(.A1(G143), .A2(new_n372), .A3(new_n351), .A4(G214), .ZN(new_n380));
  AOI21_X1  g194(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n381));
  OAI21_X1  g195(.A(G131), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(KEYINPUT85), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT17), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n371), .B(G131), .C1(new_n380), .C2(new_n381), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n374), .A2(new_n197), .A3(new_n375), .ZN(new_n386));
  NAND4_X1  g200(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n341), .A2(new_n339), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n379), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  XNOR2_X1  g203(.A(G113), .B(G122), .ZN(new_n390));
  INV_X1    g204(.A(G104), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n337), .A2(G125), .ZN(new_n393));
  INV_X1    g207(.A(G125), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G146), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n347), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT18), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n399), .A2(new_n197), .ZN(new_n400));
  OAI221_X1 g214(.A(new_n398), .B1(new_n376), .B2(new_n400), .C1(new_n382), .C2(new_n399), .ZN(new_n401));
  AND3_X1   g215(.A1(new_n389), .A2(new_n392), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n392), .B1(new_n389), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n305), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(G475), .ZN(new_n405));
  NOR2_X1   g219(.A1(G475), .A2(G902), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n396), .A2(KEYINPUT19), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT19), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n334), .A2(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(new_n411), .A3(new_n201), .ZN(new_n412));
  AND2_X1   g226(.A1(new_n412), .A2(new_n340), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n392), .B1(new_n414), .B2(new_n401), .ZN(new_n415));
  OAI21_X1  g229(.A(KEYINPUT86), .B1(new_n402), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n401), .ZN(new_n417));
  INV_X1    g231(.A(new_n392), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n389), .A2(new_n392), .A3(new_n401), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT86), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n407), .B1(new_n416), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g237(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT87), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n419), .A2(new_n420), .A3(new_n421), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n421), .B1(new_n419), .B2(new_n420), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n406), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT87), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n430), .A3(new_n424), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n407), .A2(KEYINPUT20), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n402), .B2(new_n415), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n434));
  XNOR2_X1  g248(.A(new_n433), .B(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n426), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n351), .A2(G952), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n437), .B1(G234), .B2(G237), .ZN(new_n438));
  XOR2_X1   g252(.A(KEYINPUT21), .B(G898), .Z(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  AOI211_X1 g254(.A(new_n305), .B(new_n351), .C1(G234), .C2(G237), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n318), .A2(G143), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(KEYINPUT13), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n445), .B(new_n446), .C1(G128), .C2(new_n203), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(G134), .ZN(new_n448));
  XNOR2_X1  g262(.A(G116), .B(G122), .ZN(new_n449));
  INV_X1    g263(.A(G107), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G128), .B(G143), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(KEYINPUT89), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n448), .B(new_n451), .C1(G134), .C2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT91), .B1(new_n213), .B2(G122), .ZN(new_n455));
  INV_X1    g269(.A(G122), .ZN(new_n456));
  NOR3_X1   g270(.A1(new_n456), .A2(KEYINPUT14), .A3(G116), .ZN(new_n457));
  MUX2_X1   g271(.A(new_n455), .B(KEYINPUT91), .S(new_n457), .Z(new_n458));
  OAI21_X1  g272(.A(KEYINPUT14), .B1(new_n456), .B2(G116), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(KEYINPUT90), .ZN(new_n460));
  OAI21_X1  g274(.A(G107), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n449), .A2(new_n450), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n453), .B(new_n189), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n454), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  XOR2_X1   g279(.A(KEYINPUT9), .B(G234), .Z(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(new_n467), .A2(new_n315), .A3(G953), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n465), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n454), .B(new_n468), .C1(new_n463), .C2(new_n464), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n305), .ZN(new_n473));
  INV_X1    g287(.A(G478), .ZN(new_n474));
  OR2_X1    g288(.A1(new_n474), .A2(KEYINPUT15), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n473), .B(new_n475), .ZN(new_n476));
  AND4_X1   g290(.A1(new_n405), .A2(new_n436), .A3(new_n443), .A4(new_n476), .ZN(new_n477));
  OAI21_X1  g291(.A(G210), .B1(G237), .B2(G902), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n391), .A2(G107), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n391), .A2(G107), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT76), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n483));
  OAI21_X1  g297(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n450), .A2(G104), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT3), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(KEYINPUT76), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n482), .A2(KEYINPUT3), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  OAI21_X1  g303(.A(G101), .B1(new_n484), .B2(new_n489), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n450), .A2(G104), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n491), .B1(new_n485), .B2(new_n487), .ZN(new_n492));
  NOR2_X1   g306(.A1(new_n486), .A2(KEYINPUT76), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n481), .B1(new_n483), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(G101), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n492), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n490), .A2(new_n496), .A3(KEYINPUT4), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT4), .ZN(new_n498));
  OAI211_X1 g312(.A(new_n498), .B(G101), .C1(new_n484), .C2(new_n489), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n497), .A2(new_n260), .A3(new_n499), .ZN(new_n500));
  XNOR2_X1  g314(.A(KEYINPUT79), .B(KEYINPUT5), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n217), .A2(new_n219), .A3(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n212), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n221), .B1(new_n501), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n503), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G101), .B1(new_n481), .B2(new_n491), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n506), .A2(new_n232), .A3(new_n496), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n500), .A2(new_n508), .ZN(new_n509));
  XNOR2_X1  g323(.A(G110), .B(G122), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n500), .A2(new_n508), .A3(new_n510), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT6), .A3(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n509), .A2(new_n515), .A3(new_n511), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n238), .A2(new_n239), .A3(new_n394), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT80), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n238), .A2(new_n239), .A3(KEYINPUT80), .A4(new_n394), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n208), .A2(G125), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n523), .A2(G224), .A3(new_n351), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n351), .A2(G224), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n521), .A2(new_n525), .A3(new_n522), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n514), .A2(new_n516), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n528), .A2(new_n305), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT1), .ZN(new_n530));
  AND4_X1   g344(.A1(new_n530), .A2(new_n202), .A3(new_n204), .A4(G128), .ZN(new_n531));
  AOI22_X1  g345(.A1(new_n235), .A2(G128), .B1(new_n202), .B2(new_n204), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(KEYINPUT80), .B1(new_n533), .B2(new_n394), .ZN(new_n534));
  INV_X1    g348(.A(new_n520), .ZN(new_n535));
  OAI21_X1  g349(.A(KEYINPUT81), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT81), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n519), .A2(new_n537), .A3(new_n520), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n536), .A2(new_n538), .A3(new_n522), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n539), .A2(KEYINPUT82), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT82), .B1(new_n539), .B2(new_n540), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n496), .A2(new_n507), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n506), .A2(new_n543), .A3(new_n232), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n510), .B(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n218), .A2(KEYINPUT5), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n233), .B1(new_n505), .B2(new_n546), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n544), .B(new_n545), .C1(new_n543), .C2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n521), .A2(KEYINPUT7), .A3(new_n525), .A4(new_n522), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n513), .A3(new_n549), .ZN(new_n550));
  NOR3_X1   g364(.A1(new_n541), .A2(new_n542), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n479), .B1(new_n529), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n542), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n539), .A2(KEYINPUT82), .A3(new_n540), .ZN(new_n554));
  INV_X1    g368(.A(new_n550), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n556), .A2(new_n305), .A3(new_n478), .A4(new_n528), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n552), .A2(KEYINPUT83), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(G214), .B1(G237), .B2(G902), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n529), .A2(new_n551), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT83), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n561), .A3(new_n478), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n558), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G221), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n564), .B1(new_n466), .B2(new_n305), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  XNOR2_X1  g381(.A(G110), .B(G140), .ZN(new_n568));
  AND2_X1   g382(.A1(new_n351), .A2(G227), .ZN(new_n569));
  XOR2_X1   g383(.A(new_n568), .B(new_n569), .Z(new_n570));
  NAND3_X1  g384(.A1(new_n240), .A2(new_n496), .A3(new_n507), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT10), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT77), .ZN(new_n573));
  NAND4_X1  g387(.A1(new_n497), .A2(new_n573), .A3(new_n209), .A4(new_n499), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n497), .A2(new_n209), .A3(new_n499), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT77), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n199), .A2(new_n200), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n572), .A2(new_n578), .A3(new_n576), .A4(new_n574), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n570), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  AND3_X1   g396(.A1(new_n199), .A2(KEYINPUT78), .A3(new_n200), .ZN(new_n583));
  INV_X1    g397(.A(new_n571), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n240), .B1(new_n496), .B2(new_n507), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n583), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT12), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT12), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n583), .B(new_n588), .C1(new_n584), .C2(new_n585), .ZN(new_n589));
  AND4_X1   g403(.A1(new_n581), .A2(new_n570), .A3(new_n587), .A4(new_n589), .ZN(new_n590));
  OAI211_X1 g404(.A(new_n567), .B(new_n305), .C1(new_n582), .C2(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n581), .A2(new_n587), .A3(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(new_n570), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n580), .A2(new_n581), .A3(new_n570), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(G469), .A3(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(G469), .A2(G902), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n566), .B1(new_n592), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g414(.A1(new_n563), .A2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n314), .A2(new_n370), .A3(new_n477), .A4(new_n601), .ZN(new_n602));
  XOR2_X1   g416(.A(KEYINPUT92), .B(G101), .Z(new_n603));
  XNOR2_X1  g417(.A(new_n602), .B(new_n603), .ZN(G3));
  NAND2_X1  g418(.A1(new_n552), .A2(new_n557), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT94), .B1(new_n605), .B2(new_n559), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT94), .ZN(new_n607));
  INV_X1    g421(.A(new_n559), .ZN(new_n608));
  AOI211_X1 g422(.A(new_n607), .B(new_n608), .C1(new_n552), .C2(new_n557), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n606), .A2(new_n609), .A3(new_n442), .ZN(new_n610));
  AOI21_X1  g424(.A(G478), .B1(new_n472), .B2(new_n305), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n471), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n472), .A2(KEYINPUT33), .A3(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT33), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n470), .B(new_n471), .C1(new_n612), .C2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NOR2_X1   g431(.A1(new_n474), .A2(G902), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n611), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n436), .B2(new_n405), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n610), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  AOI211_X1 g438(.A(new_n623), .B(new_n624), .C1(new_n291), .C2(new_n305), .ZN(new_n625));
  OAI21_X1  g439(.A(G472), .B1(new_n279), .B2(G902), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT93), .B1(new_n279), .B2(new_n281), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n370), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n600), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n622), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT34), .B(G104), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G6));
  NAND2_X1  g448(.A1(new_n423), .A2(new_n425), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n426), .A2(new_n635), .A3(new_n431), .ZN(new_n636));
  INV_X1    g450(.A(new_n476), .ZN(new_n637));
  AND3_X1   g451(.A1(new_n636), .A2(new_n637), .A3(new_n405), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n605), .A2(new_n559), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n607), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n605), .A2(KEYINPUT94), .A3(new_n559), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n638), .A2(new_n640), .A3(new_n443), .A4(new_n641), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n642), .A2(KEYINPUT96), .ZN(new_n643));
  INV_X1    g457(.A(KEYINPUT96), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n610), .B2(new_n638), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n631), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT97), .ZN(new_n647));
  XOR2_X1   g461(.A(KEYINPUT35), .B(G107), .Z(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  OR2_X1    g463(.A1(new_n353), .A2(KEYINPUT36), .ZN(new_n650));
  XNOR2_X1  g464(.A(new_n349), .B(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(new_n368), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n361), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n601), .A2(new_n628), .A3(new_n477), .A4(new_n654), .ZN(new_n655));
  XOR2_X1   g469(.A(KEYINPUT37), .B(G110), .Z(new_n656));
  XNOR2_X1  g470(.A(new_n655), .B(new_n656), .ZN(G12));
  AND2_X1   g471(.A1(new_n581), .A2(new_n570), .ZN(new_n658));
  AOI22_X1  g472(.A1(new_n658), .A2(new_n580), .B1(new_n593), .B2(new_n594), .ZN(new_n659));
  OAI21_X1  g473(.A(G469), .B1(new_n659), .B2(G902), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n565), .B1(new_n660), .B2(new_n591), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n314), .A2(new_n661), .A3(new_n654), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT98), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n640), .A2(new_n641), .ZN(new_n664));
  INV_X1    g478(.A(G900), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n441), .A2(new_n665), .ZN(new_n666));
  INV_X1    g480(.A(new_n438), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n636), .A2(new_n637), .A3(new_n405), .A4(new_n668), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n663), .B1(new_n664), .B2(new_n669), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n606), .A2(new_n609), .ZN(new_n671));
  INV_X1    g485(.A(new_n669), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n672), .A3(KEYINPUT98), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n662), .B1(new_n670), .B2(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(new_n318), .ZN(G30));
  NAND2_X1  g489(.A1(new_n271), .A2(new_n298), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n286), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(new_n624), .B1(new_n677), .B2(new_n305), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n294), .A2(new_n313), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n668), .B(KEYINPUT39), .Z(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n661), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT99), .B(KEYINPUT40), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n558), .A2(new_n562), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(KEYINPUT38), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n476), .B1(new_n436), .B2(new_n405), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n689), .A2(new_n559), .A3(new_n653), .ZN(new_n690));
  OR4_X1    g504(.A1(new_n681), .A2(new_n686), .A3(new_n688), .A4(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G143), .ZN(G45));
  INV_X1    g506(.A(new_n662), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n620), .A2(new_n668), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n664), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G146), .ZN(G48));
  NOR2_X1   g511(.A1(new_n582), .A2(new_n590), .ZN(new_n698));
  OAI21_X1  g512(.A(G469), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(new_n566), .A3(new_n591), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n314), .A2(new_n370), .A3(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n622), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT41), .B(G113), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(KEYINPUT100), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n704), .B(new_n706), .ZN(G15));
  NAND2_X1  g521(.A1(new_n642), .A2(KEYINPUT96), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n610), .A2(new_n644), .A3(new_n638), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n702), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n213), .ZN(G18));
  NOR3_X1   g525(.A1(new_n606), .A2(new_n609), .A3(new_n700), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n712), .A2(new_n314), .A3(new_n477), .A4(new_n654), .ZN(new_n713));
  XOR2_X1   g527(.A(KEYINPUT101), .B(G119), .Z(new_n714));
  XNOR2_X1  g528(.A(new_n713), .B(new_n714), .ZN(G21));
  AND2_X1   g529(.A1(new_n689), .A2(new_n443), .ZN(new_n716));
  INV_X1    g530(.A(new_n361), .ZN(new_n717));
  INV_X1    g531(.A(new_n369), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n717), .A2(KEYINPUT104), .A3(new_n718), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT104), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n720), .B1(new_n361), .B2(new_n369), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n300), .A2(KEYINPUT102), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  OAI21_X1  g538(.A(new_n724), .B1(new_n296), .B2(new_n299), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n723), .A2(new_n725), .A3(new_n271), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n267), .A2(new_n270), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n281), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT103), .B(G472), .Z(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n291), .B2(new_n305), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n722), .A2(new_n728), .A3(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n712), .A2(new_n716), .A3(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  NOR3_X1   g547(.A1(new_n728), .A2(new_n653), .A3(new_n730), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n620), .A3(new_n668), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n671), .A2(new_n701), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(new_n394), .ZN(G27));
  INV_X1    g552(.A(KEYINPUT42), .ZN(new_n739));
  AND3_X1   g553(.A1(new_n620), .A2(new_n739), .A3(new_n668), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n687), .A2(new_n559), .A3(new_n661), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n370), .A3(new_n314), .A4(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n608), .B1(new_n558), .B2(new_n562), .ZN(new_n743));
  NAND4_X1  g557(.A1(new_n743), .A2(new_n620), .A3(new_n661), .A4(new_n668), .ZN(new_n744));
  AND2_X1   g558(.A1(new_n719), .A2(new_n721), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT32), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n746), .B1(new_n279), .B2(new_n281), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n280), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n306), .B1(new_n300), .B2(new_n302), .ZN(new_n750));
  OAI21_X1  g564(.A(new_n305), .B1(new_n308), .B2(new_n309), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n624), .B1(new_n752), .B2(new_n307), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n745), .B1(new_n749), .B2(new_n753), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT42), .B1(new_n744), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n742), .A2(new_n755), .A3(KEYINPUT105), .ZN(new_n756));
  INV_X1    g570(.A(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT105), .B1(new_n742), .B2(new_n755), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n197), .ZN(G33));
  NAND4_X1  g574(.A1(new_n314), .A2(new_n741), .A3(new_n370), .A4(new_n672), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT106), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G134), .ZN(G36));
  INV_X1    g578(.A(new_n619), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n765), .A2(new_n436), .A3(new_n405), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  NOR2_X1   g581(.A1(new_n628), .A2(new_n653), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n769), .A2(KEYINPUT44), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(KEYINPUT44), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n743), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT108), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT108), .ZN(new_n774));
  NAND4_X1  g588(.A1(new_n770), .A2(new_n774), .A3(new_n743), .A4(new_n771), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n659), .A2(KEYINPUT45), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n659), .A2(KEYINPUT45), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n776), .A2(G469), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n598), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n591), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  AND2_X1   g595(.A1(new_n781), .A2(KEYINPUT107), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n779), .A2(new_n780), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n783), .B1(new_n781), .B2(KEYINPUT107), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n566), .B1(new_n782), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n785), .A2(new_n682), .ZN(new_n786));
  INV_X1    g600(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n773), .A2(new_n775), .A3(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  NAND2_X1  g603(.A1(new_n785), .A2(KEYINPUT47), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT47), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n566), .C1(new_n782), .C2(new_n784), .ZN(new_n792));
  INV_X1    g606(.A(new_n743), .ZN(new_n793));
  NOR4_X1   g607(.A1(new_n314), .A2(new_n694), .A3(new_n793), .A4(new_n370), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n790), .A2(new_n792), .A3(new_n794), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(KEYINPUT109), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  NAND3_X1  g611(.A1(new_n745), .A2(new_n559), .A3(new_n566), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n699), .A2(new_n591), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n799), .A2(KEYINPUT49), .ZN(new_n801));
  NOR4_X1   g615(.A1(new_n798), .A2(new_n800), .A3(new_n766), .A4(new_n801), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n802), .A2(new_n681), .A3(new_n688), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n767), .A2(new_n438), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n793), .A2(new_n700), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(new_n734), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n681), .A2(new_n805), .A3(new_n370), .A4(new_n438), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n436), .A2(new_n405), .A3(new_n619), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n804), .A2(new_n731), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n688), .A2(new_n608), .A3(new_n701), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT50), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(KEYINPUT50), .A3(new_n812), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n810), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  AOI21_X1  g631(.A(KEYINPUT51), .B1(new_n817), .B2(KEYINPUT116), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n799), .A2(new_n566), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n819), .B1(new_n790), .B2(new_n792), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n811), .A2(new_n743), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n818), .B(new_n822), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n443), .A2(new_n558), .A3(new_n559), .A4(new_n562), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n436), .A2(new_n637), .A3(new_n405), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n628), .A2(new_n824), .A3(new_n630), .A4(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n655), .A2(KEYINPUT110), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT110), .B1(new_n655), .B2(new_n826), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n628), .A2(new_n824), .A3(new_n620), .A4(new_n630), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n602), .A2(new_n829), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n827), .A2(new_n828), .A3(new_n830), .ZN(new_n831));
  OAI211_X1 g645(.A(new_n713), .B(new_n732), .C1(new_n621), .C2(new_n702), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n710), .ZN(new_n833));
  INV_X1    g647(.A(new_n741), .ZN(new_n834));
  AND4_X1   g648(.A1(new_n405), .A2(new_n636), .A3(new_n476), .A4(new_n668), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n314), .A2(new_n654), .A3(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n834), .B1(new_n836), .B2(new_n735), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n831), .A2(new_n833), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n763), .B1(new_n757), .B2(new_n758), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT111), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  INV_X1    g657(.A(KEYINPUT52), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n670), .A2(new_n673), .ZN(new_n845));
  AOI21_X1  g659(.A(new_n737), .B1(new_n845), .B2(new_n693), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n671), .A2(new_n689), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n653), .A2(new_n668), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n848), .B1(new_n600), .B2(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(new_n668), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n361), .A2(new_n652), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n661), .A2(KEYINPUT113), .A3(new_n852), .ZN(new_n853));
  AND2_X1   g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n847), .A2(new_n854), .A3(KEYINPUT114), .A4(new_n680), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT114), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n671), .A2(new_n850), .A3(new_n689), .A4(new_n853), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n856), .B1(new_n857), .B2(new_n681), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  AND4_X1   g673(.A1(new_n844), .A2(new_n846), .A3(new_n859), .A4(new_n696), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT112), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n861), .B1(new_n674), .B2(new_n737), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n735), .A2(new_n736), .ZN(new_n863));
  NOR4_X1   g677(.A1(new_n669), .A2(new_n606), .A3(new_n609), .A4(new_n663), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT98), .B1(new_n671), .B2(new_n672), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(KEYINPUT112), .B(new_n863), .C1(new_n866), .C2(new_n662), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n862), .A2(new_n867), .A3(new_n696), .A4(new_n859), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n860), .B1(KEYINPUT52), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n841), .A2(KEYINPUT111), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n842), .A2(new_n843), .A3(new_n869), .A4(new_n870), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n761), .B(KEYINPUT106), .ZN(new_n872));
  INV_X1    g686(.A(new_n758), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n872), .B1(new_n873), .B2(new_n756), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n874), .A2(new_n831), .A3(new_n833), .A4(new_n838), .ZN(new_n875));
  AOI22_X1  g689(.A1(new_n855), .A2(new_n858), .B1(new_n693), .B2(new_n695), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n846), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT52), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n844), .A3(new_n846), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT53), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n871), .A2(new_n881), .A3(KEYINPUT54), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n843), .B1(new_n875), .B2(new_n880), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n703), .B1(new_n643), .B2(new_n645), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n713), .A2(new_n732), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT115), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n885), .A2(new_n886), .A3(new_n887), .A4(new_n704), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT115), .B1(new_n832), .B2(new_n710), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n742), .A2(new_n755), .A3(KEYINPUT53), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n891), .A2(new_n837), .ZN(new_n892));
  INV_X1    g706(.A(new_n827), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n828), .A2(new_n830), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n892), .A2(new_n763), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n890), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n869), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n883), .A2(new_n884), .A3(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n882), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n754), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n806), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT117), .Z(new_n902));
  OR2_X1    g716(.A1(new_n902), .A2(KEYINPUT48), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(KEYINPUT48), .ZN(new_n904));
  INV_X1    g718(.A(new_n620), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n808), .A2(new_n905), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n437), .B(new_n906), .C1(new_n811), .C2(new_n712), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n903), .A2(new_n904), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n823), .A2(new_n899), .A3(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(G952), .A2(G953), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(KEYINPUT118), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n803), .B1(new_n909), .B2(new_n911), .ZN(G75));
  XNOR2_X1  g726(.A(KEYINPUT119), .B(KEYINPUT55), .ZN(new_n913));
  INV_X1    g727(.A(G210), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n914), .B(new_n305), .C1(new_n883), .C2(new_n897), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n915), .B2(KEYINPUT56), .ZN(new_n916));
  INV_X1    g730(.A(KEYINPUT56), .ZN(new_n917));
  INV_X1    g731(.A(new_n913), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n883), .A2(new_n897), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(G902), .ZN(new_n920));
  OAI211_X1 g734(.A(new_n917), .B(new_n918), .C1(new_n920), .C2(new_n914), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n514), .A2(new_n516), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n527), .ZN(new_n923));
  AND3_X1   g737(.A1(new_n916), .A2(new_n921), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n923), .B1(new_n916), .B2(new_n921), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n351), .A2(G952), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(G51));
  INV_X1    g741(.A(KEYINPUT120), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n920), .A2(new_n778), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n598), .B(KEYINPUT57), .Z(new_n930));
  NAND2_X1  g744(.A1(new_n868), .A2(KEYINPUT52), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n896), .A2(new_n879), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n844), .B1(new_n876), .B2(new_n846), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n860), .A2(new_n933), .ZN(new_n934));
  AOI21_X1  g748(.A(KEYINPUT53), .B1(new_n934), .B2(new_n841), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n932), .A2(new_n935), .A3(KEYINPUT54), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n884), .B1(new_n883), .B2(new_n897), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n930), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n698), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n929), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n928), .B1(new_n940), .B2(new_n926), .ZN(new_n941));
  INV_X1    g755(.A(new_n926), .ZN(new_n942));
  OAI21_X1  g756(.A(KEYINPUT54), .B1(new_n932), .B2(new_n935), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n898), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n698), .B1(new_n944), .B2(new_n930), .ZN(new_n945));
  OAI211_X1 g759(.A(KEYINPUT120), .B(new_n942), .C1(new_n945), .C2(new_n929), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n941), .A2(new_n946), .ZN(G54));
  AND4_X1   g761(.A1(KEYINPUT58), .A2(new_n919), .A3(G475), .A4(G902), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n416), .A2(new_n422), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n949), .ZN(new_n951));
  NOR3_X1   g765(.A1(new_n950), .A2(new_n951), .A3(new_n926), .ZN(G60));
  XNOR2_X1  g766(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n474), .A2(new_n305), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n953), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n617), .B1(new_n899), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n617), .A2(new_n956), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n958), .B1(new_n943), .B2(new_n898), .ZN(new_n959));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n942), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  AOI211_X1 g775(.A(KEYINPUT122), .B(new_n958), .C1(new_n943), .C2(new_n898), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT123), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(new_n958), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n964), .B1(new_n936), .B2(new_n937), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT122), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n944), .A2(new_n960), .A3(new_n964), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n966), .A2(new_n967), .A3(new_n942), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n957), .B1(new_n963), .B2(new_n969), .ZN(G63));
  XNOR2_X1  g784(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n315), .A2(new_n305), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n971), .B(new_n972), .Z(new_n973));
  AOI21_X1  g787(.A(new_n973), .B1(new_n883), .B2(new_n897), .ZN(new_n974));
  INV_X1    g788(.A(new_n651), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n926), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n364), .A2(new_n366), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n976), .B1(new_n977), .B2(new_n974), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT61), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n978), .B(new_n979), .ZN(G66));
  INV_X1    g794(.A(G224), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n440), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n831), .A2(new_n833), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n982), .B1(new_n984), .B2(G953), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n922), .B1(G898), .B2(new_n351), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  AOI21_X1  g801(.A(new_n351), .B1(G227), .B2(G900), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n409), .A2(new_n411), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n255), .B(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(G900), .B2(G953), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n787), .A2(new_n900), .A3(new_n847), .ZN(new_n992));
  AND3_X1   g806(.A1(new_n862), .A2(new_n696), .A3(new_n867), .ZN(new_n993));
  AND2_X1   g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  XNOR2_X1  g808(.A(new_n840), .B(KEYINPUT126), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n994), .A2(new_n788), .A3(new_n796), .A4(new_n995), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n991), .B1(new_n996), .B2(G953), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT127), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n990), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n998), .B1(new_n997), .B2(KEYINPUT125), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n988), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g817(.A1(new_n825), .A2(new_n620), .ZN(new_n1004));
  NOR3_X1   g818(.A1(new_n1004), .A2(new_n684), .A3(new_n793), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n1005), .A2(new_n370), .A3(new_n314), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n788), .A2(new_n796), .A3(new_n1006), .ZN(new_n1007));
  AND2_X1   g821(.A1(new_n993), .A2(new_n691), .ZN(new_n1008));
  OR2_X1    g822(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(KEYINPUT62), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1007), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n990), .B1(new_n1011), .B2(G953), .ZN(new_n1012));
  INV_X1    g826(.A(new_n988), .ZN(new_n1013));
  NAND4_X1  g827(.A1(new_n1012), .A2(KEYINPUT125), .A3(new_n1013), .A4(new_n997), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n1003), .A2(new_n1014), .ZN(G72));
  NAND2_X1  g829(.A1(new_n1011), .A2(new_n984), .ZN(new_n1016));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  AOI211_X1 g832(.A(new_n269), .B(new_n261), .C1(new_n1016), .C2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n996), .B2(new_n983), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n268), .A2(new_n245), .A3(new_n266), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n261), .B(new_n266), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n871), .A2(new_n881), .A3(new_n1018), .A4(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1022), .A2(new_n942), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1019), .A2(new_n1025), .ZN(G57));
endmodule


