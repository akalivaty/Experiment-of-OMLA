//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 0 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n866, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n878, new_n879,
    new_n880, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905;
  INV_X1    g000(.A(KEYINPUT84), .ZN(new_n202));
  XOR2_X1   g001(.A(G211gat), .B(G218gat), .Z(new_n203));
  INV_X1    g002(.A(KEYINPUT68), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g004(.A(G211gat), .B(G218gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT68), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT22), .ZN(new_n210));
  INV_X1    g009(.A(G211gat), .ZN(new_n211));
  INV_X1    g010(.A(G218gat), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n209), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n208), .A2(new_n214), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n205), .A2(new_n213), .A3(new_n209), .A4(new_n207), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NOR2_X1   g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n218), .B(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G183gat), .A2(G190gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT24), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n224), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n228));
  AND2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT25), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT26), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n218), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n222), .A2(new_n231), .A3(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(KEYINPUT27), .B(G183gat), .ZN(new_n235));
  INV_X1    g034(.A(G190gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT28), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT28), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n239), .A3(new_n236), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n234), .A2(new_n238), .A3(new_n226), .A4(new_n240), .ZN(new_n241));
  OR2_X1    g040(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n228), .A2(KEYINPUT64), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n242), .A2(new_n227), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT25), .ZN(new_n245));
  NAND4_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n222), .A4(new_n220), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n230), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(G226gat), .ZN(new_n248));
  INV_X1    g047(.A(G233gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n247), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT29), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n247), .A2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n250), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n252), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AOI211_X1 g055(.A(KEYINPUT69), .B(new_n250), .C1(new_n247), .C2(new_n253), .ZN(new_n257));
  OAI211_X1 g056(.A(new_n217), .B(new_n251), .C1(new_n256), .C2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(new_n251), .ZN(new_n259));
  AOI21_X1  g058(.A(new_n250), .B1(new_n247), .B2(new_n253), .ZN(new_n260));
  OAI211_X1 g059(.A(new_n216), .B(new_n215), .C1(new_n259), .C2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n258), .A2(new_n261), .ZN(new_n262));
  XNOR2_X1  g061(.A(G8gat), .B(G36gat), .ZN(new_n263));
  INV_X1    g062(.A(G92gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT70), .B(G64gat), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n265), .B(new_n266), .Z(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(KEYINPUT30), .B1(new_n262), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(new_n268), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G78gat), .B(G106gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n272), .B(G22gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(new_n273), .B(KEYINPUT81), .ZN(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(KEYINPUT31), .B(G50gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n215), .A2(new_n253), .A3(new_n216), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT79), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT3), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT79), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n215), .A2(new_n281), .A3(new_n253), .A4(new_n216), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n279), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G155gat), .A2(G162gat), .ZN(new_n284));
  INV_X1    g083(.A(G155gat), .ZN(new_n285));
  INV_X1    g084(.A(G162gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n284), .B1(new_n287), .B2(KEYINPUT2), .ZN(new_n288));
  INV_X1    g087(.A(G141gat), .ZN(new_n289));
  INV_X1    g088(.A(G148gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT73), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT73), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G148gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n289), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n290), .A2(G141gat), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n288), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT72), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n284), .A2(new_n297), .A3(KEYINPUT2), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(G141gat), .B(G148gat), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n297), .B1(new_n284), .B2(KEYINPUT2), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n284), .A2(KEYINPUT71), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G155gat), .A3(G162gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(new_n287), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n296), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n283), .A2(new_n308), .ZN(new_n309));
  OAI211_X1 g108(.A(new_n296), .B(new_n280), .C1(new_n302), .C2(new_n307), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n253), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n311), .A2(new_n217), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT80), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n217), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT80), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n309), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G228gat), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n318), .A2(new_n249), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n284), .A2(KEYINPUT2), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n321), .A2(KEYINPUT72), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n322), .A2(new_n298), .ZN(new_n323));
  OAI211_X1 g122(.A(new_n287), .B(new_n306), .C1(new_n323), .C2(new_n300), .ZN(new_n324));
  AOI22_X1  g123(.A1(new_n278), .A2(new_n280), .B1(new_n296), .B2(new_n324), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n325), .A2(new_n312), .A3(new_n319), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n277), .B1(new_n320), .B2(new_n327), .ZN(new_n328));
  AOI211_X1 g127(.A(new_n276), .B(new_n326), .C1(new_n317), .C2(new_n319), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n275), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n319), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n314), .A2(new_n316), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n331), .B1(new_n332), .B2(new_n309), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n276), .B1(new_n333), .B2(new_n326), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n320), .A2(new_n277), .A3(new_n327), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n334), .A2(new_n274), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(G15gat), .B(G43gat), .ZN(new_n337));
  INV_X1    g136(.A(G71gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT67), .ZN(new_n340));
  INV_X1    g139(.A(G99gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(G227gat), .A2(G233gat), .ZN(new_n343));
  XOR2_X1   g142(.A(G127gat), .B(G134gat), .Z(new_n344));
  XNOR2_X1  g143(.A(G113gat), .B(G120gat), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n344), .B1(KEYINPUT1), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G113gat), .B(G120gat), .Z(new_n347));
  INV_X1    g146(.A(KEYINPUT1), .ZN(new_n348));
  XNOR2_X1  g147(.A(G127gat), .B(G134gat), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n247), .A2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(new_n346), .A2(new_n350), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n230), .A2(new_n241), .A3(new_n353), .A4(new_n246), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n343), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n342), .B(KEYINPUT66), .C1(new_n355), .C2(KEYINPUT33), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n352), .A2(new_n343), .A3(new_n354), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT32), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT34), .B1(new_n355), .B2(new_n360), .ZN(new_n361));
  OR3_X1    g160(.A1(new_n355), .A2(new_n360), .A3(KEYINPUT34), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n356), .A2(new_n357), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n359), .A2(new_n361), .A3(new_n362), .A4(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n362), .A2(new_n361), .ZN(new_n365));
  INV_X1    g164(.A(new_n363), .ZN(new_n366));
  OAI21_X1  g165(.A(new_n365), .B1(new_n366), .B2(new_n358), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n330), .A2(new_n336), .A3(new_n364), .A4(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(G225gat), .A2(G233gat), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n308), .A2(new_n351), .ZN(new_n371));
  AOI22_X1  g170(.A1(new_n324), .A2(new_n296), .B1(new_n350), .B2(new_n346), .ZN(new_n372));
  OAI211_X1 g171(.A(KEYINPUT74), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT4), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n308), .B2(new_n351), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n353), .A2(KEYINPUT4), .A3(new_n324), .A4(new_n296), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n310), .A2(new_n351), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n280), .B1(new_n324), .B2(new_n296), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n375), .B(new_n376), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n373), .B1(new_n379), .B2(new_n370), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n353), .A2(new_n296), .A3(new_n324), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n308), .A2(new_n351), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n369), .B1(new_n381), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT5), .B1(new_n383), .B2(KEYINPUT74), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT75), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT5), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT74), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT75), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n308), .A2(KEYINPUT3), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n391), .A2(new_n351), .A3(new_n310), .ZN(new_n392));
  NAND4_X1  g191(.A1(new_n392), .A2(new_n369), .A3(new_n375), .A4(new_n376), .ZN(new_n393));
  NAND4_X1  g192(.A1(new_n389), .A2(new_n390), .A3(new_n393), .A4(new_n373), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n385), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n375), .A2(new_n376), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n377), .A2(new_n378), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n398), .A2(new_n399), .A3(new_n386), .A4(new_n369), .ZN(new_n400));
  OAI21_X1  g199(.A(KEYINPUT76), .B1(new_n393), .B2(KEYINPUT5), .ZN(new_n401));
  AND2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G1gat), .B(G29gat), .ZN(new_n403));
  XNOR2_X1  g202(.A(new_n403), .B(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT0), .B(G57gat), .ZN(new_n405));
  XOR2_X1   g204(.A(new_n404), .B(new_n405), .Z(new_n406));
  NAND3_X1  g205(.A1(new_n395), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT6), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT77), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT77), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n407), .A2(new_n411), .A3(new_n408), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n400), .A2(new_n401), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n413), .B1(new_n385), .B2(new_n394), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT78), .B1(new_n414), .B2(new_n406), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n395), .A2(new_n402), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT78), .ZN(new_n417));
  INV_X1    g216(.A(new_n406), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND4_X1  g218(.A1(new_n410), .A2(new_n412), .A3(new_n415), .A4(new_n419), .ZN(new_n420));
  NOR3_X1   g219(.A1(new_n414), .A2(new_n408), .A3(new_n406), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AOI211_X1 g221(.A(new_n271), .B(new_n368), .C1(new_n420), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT35), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n202), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  AND3_X1   g224(.A1(new_n416), .A2(KEYINPUT82), .A3(new_n418), .ZN(new_n426));
  AOI21_X1  g225(.A(KEYINPUT82), .B1(new_n416), .B2(new_n418), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n408), .B(new_n407), .C1(new_n426), .C2(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n428), .A2(new_n422), .ZN(new_n429));
  INV_X1    g228(.A(new_n271), .ZN(new_n430));
  INV_X1    g229(.A(new_n368), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n429), .A2(new_n424), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n419), .ZN(new_n433));
  AND3_X1   g232(.A1(new_n407), .A2(new_n411), .A3(new_n408), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n411), .B1(new_n407), .B2(new_n408), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n430), .B(new_n431), .C1(new_n436), .C2(new_n421), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n437), .A2(KEYINPUT84), .A3(KEYINPUT35), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n425), .A2(new_n432), .A3(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n270), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n258), .A2(KEYINPUT37), .A3(new_n261), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n267), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT83), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n441), .A2(new_n444), .A3(new_n267), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n262), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n443), .A2(new_n445), .A3(new_n447), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n440), .B1(new_n448), .B2(KEYINPUT38), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n259), .A2(new_n260), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n217), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n256), .A2(new_n257), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n452), .A2(new_n259), .ZN(new_n453));
  OAI211_X1 g252(.A(KEYINPUT37), .B(new_n451), .C1(new_n453), .C2(new_n217), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT38), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n454), .A2(new_n455), .A3(new_n267), .A4(new_n447), .ZN(new_n456));
  NAND4_X1  g255(.A1(new_n449), .A2(new_n428), .A3(new_n422), .A4(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n330), .A2(new_n336), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  OAI211_X1 g258(.A(KEYINPUT39), .B(new_n369), .C1(new_n371), .C2(new_n372), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n379), .B(KEYINPUT39), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n406), .B(new_n460), .C1(new_n461), .C2(new_n369), .ZN(new_n462));
  XNOR2_X1  g261(.A(new_n462), .B(KEYINPUT40), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n271), .B(new_n463), .C1(new_n427), .C2(new_n426), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n457), .A2(new_n459), .A3(new_n464), .ZN(new_n465));
  AND2_X1   g264(.A1(new_n364), .A2(new_n367), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT36), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n271), .B1(new_n420), .B2(new_n422), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n465), .B(new_n467), .C1(new_n459), .C2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n439), .A2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(G43gat), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n471), .A2(G50gat), .ZN(new_n472));
  XOR2_X1   g271(.A(KEYINPUT86), .B(G50gat), .Z(new_n473));
  OAI21_X1  g272(.A(new_n472), .B1(new_n473), .B2(G43gat), .ZN(new_n474));
  XOR2_X1   g273(.A(KEYINPUT85), .B(KEYINPUT15), .Z(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n471), .A2(G50gat), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n472), .A2(KEYINPUT15), .A3(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT14), .ZN(new_n479));
  INV_X1    g278(.A(G29gat), .ZN(new_n480));
  INV_X1    g279(.A(G36gat), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT87), .ZN(new_n483));
  OR2_X1    g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n483), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G29gat), .A2(G36gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT88), .Z(new_n489));
  NAND4_X1  g288(.A1(new_n476), .A2(new_n478), .A3(new_n487), .A4(new_n489), .ZN(new_n490));
  AOI22_X1  g289(.A1(new_n482), .A2(new_n485), .B1(G29gat), .B2(G36gat), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(new_n478), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT17), .ZN(new_n494));
  XNOR2_X1  g293(.A(G15gat), .B(G22gat), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT16), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n495), .B1(new_n496), .B2(G1gat), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT89), .ZN(new_n498));
  INV_X1    g297(.A(G8gat), .ZN(new_n499));
  OAI221_X1 g298(.A(new_n497), .B1(new_n498), .B2(new_n499), .C1(G1gat), .C2(new_n495), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n497), .B2(new_n498), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n497), .B1(G1gat), .B2(new_n495), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n494), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n500), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n493), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(G229gat), .A2(G233gat), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT90), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n510), .B1(new_n511), .B2(KEYINPUT18), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT18), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n512), .B1(KEYINPUT90), .B2(new_n513), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n493), .A2(new_n505), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT91), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(new_n506), .ZN(new_n517));
  XOR2_X1   g316(.A(new_n508), .B(KEYINPUT13), .Z(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n519), .B(KEYINPUT92), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT18), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  XNOR2_X1  g321(.A(G113gat), .B(G141gat), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(G197gat), .ZN(new_n524));
  XNOR2_X1  g323(.A(KEYINPUT11), .B(G169gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(new_n524), .B(new_n525), .ZN(new_n526));
  XOR2_X1   g325(.A(new_n526), .B(KEYINPUT12), .Z(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n522), .B(new_n528), .ZN(new_n529));
  OR2_X1    g328(.A1(G57gat), .A2(G64gat), .ZN(new_n530));
  NAND2_X1  g329(.A1(G57gat), .A2(G64gat), .ZN(new_n531));
  AND2_X1   g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  OAI211_X1 g331(.A(new_n530), .B(new_n531), .C1(new_n532), .C2(KEYINPUT9), .ZN(new_n533));
  OAI21_X1  g332(.A(KEYINPUT93), .B1(G71gat), .B2(G78gat), .ZN(new_n534));
  AND2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(G71gat), .A2(G78gat), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n532), .A2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OR2_X1    g337(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n535), .A2(new_n538), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n505), .B1(new_n541), .B2(KEYINPUT21), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(KEYINPUT95), .ZN(new_n543));
  NAND2_X1  g342(.A1(G231gat), .A2(G233gat), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n543), .B(new_n544), .ZN(new_n545));
  XOR2_X1   g344(.A(G127gat), .B(G155gat), .Z(new_n546));
  XNOR2_X1  g345(.A(new_n546), .B(KEYINPUT20), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  XNOR2_X1  g347(.A(new_n545), .B(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n541), .A2(KEYINPUT21), .ZN(new_n550));
  XOR2_X1   g349(.A(G183gat), .B(G211gat), .Z(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT94), .ZN(new_n552));
  XOR2_X1   g351(.A(new_n552), .B(KEYINPUT19), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n550), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n549), .B(new_n554), .ZN(new_n555));
  XOR2_X1   g354(.A(KEYINPUT97), .B(KEYINPUT7), .Z(new_n556));
  INV_X1    g355(.A(G85gat), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n557), .A2(new_n264), .ZN(new_n558));
  NAND2_X1  g357(.A1(G99gat), .A2(G106gat), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n556), .A2(new_n558), .B1(KEYINPUT8), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n264), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n560), .B(new_n561), .C1(new_n558), .C2(new_n556), .ZN(new_n562));
  XOR2_X1   g361(.A(G99gat), .B(G106gat), .Z(new_n563));
  XOR2_X1   g362(.A(new_n562), .B(new_n563), .Z(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n494), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G232gat), .A2(G233gat), .ZN(new_n567));
  XOR2_X1   g366(.A(new_n567), .B(KEYINPUT96), .Z(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n564), .A2(new_n493), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n566), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  XOR2_X1   g371(.A(G190gat), .B(G218gat), .Z(new_n573));
  XNOR2_X1  g372(.A(new_n572), .B(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n569), .A2(KEYINPUT41), .ZN(new_n575));
  XOR2_X1   g374(.A(G134gat), .B(G162gat), .Z(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  XOR2_X1   g376(.A(new_n574), .B(new_n577), .Z(new_n578));
  NOR2_X1   g377(.A1(new_n555), .A2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(KEYINPUT99), .B1(new_n562), .B2(KEYINPUT98), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT98), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT99), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n581), .B1(new_n563), .B2(new_n582), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n580), .A2(new_n563), .B1(new_n562), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n541), .ZN(new_n585));
  MUX2_X1   g384(.A(new_n584), .B(new_n564), .S(new_n585), .Z(new_n586));
  INV_X1    g385(.A(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT100), .ZN(new_n589));
  NOR3_X1   g388(.A1(new_n565), .A2(new_n587), .A3(new_n585), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(G230gat), .ZN(new_n593));
  NOR2_X1   g392(.A1(new_n593), .A2(new_n249), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  OR2_X1    g395(.A1(new_n586), .A2(new_n595), .ZN(new_n597));
  XNOR2_X1  g396(.A(G120gat), .B(G148gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(G176gat), .B(G204gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n596), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n588), .A2(KEYINPUT100), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n588), .A2(KEYINPUT100), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n590), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n597), .B1(new_n605), .B2(new_n594), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(new_n600), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n602), .A2(new_n607), .A3(KEYINPUT101), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(KEYINPUT101), .B1(new_n602), .B2(new_n607), .ZN(new_n610));
  NOR2_X1   g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n470), .A2(new_n529), .A3(new_n579), .A4(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT102), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n436), .A2(new_n421), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g415(.A1(new_n613), .A2(new_n271), .ZN(new_n617));
  NAND2_X1  g416(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n496), .A2(new_n499), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n617), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(KEYINPUT42), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n620), .A2(new_n621), .ZN(new_n623));
  OAI211_X1 g422(.A(new_n622), .B(new_n623), .C1(new_n499), .C2(new_n617), .ZN(G1325gat));
  AOI21_X1  g423(.A(G15gat), .B1(new_n613), .B2(new_n466), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n467), .B(KEYINPUT103), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AND2_X1   g426(.A1(new_n613), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n625), .B1(G15gat), .B2(new_n628), .ZN(G1326gat));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n458), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT43), .B(G22gat), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n630), .B(new_n631), .ZN(G1327gat));
  INV_X1    g431(.A(new_n578), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n439), .B2(new_n469), .ZN(new_n634));
  OR2_X1    g433(.A1(new_n634), .A2(KEYINPUT44), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(KEYINPUT44), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n611), .A2(new_n529), .A3(new_n555), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  INV_X1    g439(.A(new_n614), .ZN(new_n641));
  OAI21_X1  g440(.A(G29gat), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n470), .A2(new_n578), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n638), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n644), .A2(new_n480), .A3(new_n614), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(KEYINPUT45), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n642), .A2(new_n646), .ZN(G1328gat));
  NAND3_X1  g446(.A1(new_n644), .A2(new_n481), .A3(new_n271), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT104), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n648), .B1(new_n649), .B2(KEYINPUT46), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(KEYINPUT46), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  AND2_X1   g451(.A1(new_n637), .A2(new_n639), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(new_n271), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT105), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n652), .B1(new_n655), .B2(new_n481), .ZN(G1329gat));
  OR3_X1    g455(.A1(new_n640), .A2(KEYINPUT106), .A3(new_n467), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT106), .B1(new_n640), .B2(new_n467), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(G43gat), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n644), .A2(new_n471), .A3(new_n466), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n659), .A2(KEYINPUT47), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT47), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n471), .B1(new_n653), .B2(new_n627), .ZN(new_n663));
  INV_X1    g462(.A(new_n660), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n662), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n661), .A2(new_n665), .ZN(G1330gat));
  INV_X1    g465(.A(new_n473), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(new_n640), .B2(new_n459), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n644), .A2(new_n473), .A3(new_n458), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(KEYINPUT48), .A3(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(KEYINPUT107), .ZN(new_n671));
  AOI21_X1  g470(.A(KEYINPUT48), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT108), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AOI211_X1 g473(.A(KEYINPUT108), .B(KEYINPUT48), .C1(new_n668), .C2(new_n671), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n670), .B1(new_n674), .B2(new_n675), .ZN(G1331gat));
  NOR2_X1   g475(.A1(new_n611), .A2(new_n529), .ZN(new_n677));
  AND3_X1   g476(.A1(new_n470), .A2(new_n579), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n678), .A2(new_n614), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n271), .ZN(new_n681));
  OAI21_X1  g480(.A(new_n681), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT49), .B(G64gat), .Z(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n681), .B2(new_n683), .ZN(G1333gat));
  AOI21_X1  g483(.A(G71gat), .B1(new_n678), .B2(new_n466), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n626), .A2(new_n338), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n685), .B1(new_n678), .B2(new_n686), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g487(.A1(new_n678), .A2(new_n458), .ZN(new_n689));
  XOR2_X1   g488(.A(KEYINPUT109), .B(G78gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n689), .B(new_n690), .ZN(G1335gat));
  NAND4_X1  g490(.A1(new_n635), .A2(new_n555), .A3(new_n636), .A4(new_n677), .ZN(new_n692));
  OAI21_X1  g491(.A(G85gat), .B1(new_n692), .B2(new_n641), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT51), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n470), .A2(KEYINPUT110), .A3(new_n578), .ZN(new_n695));
  INV_X1    g494(.A(new_n529), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n555), .B1(new_n634), .B2(KEYINPUT110), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n694), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n529), .B1(new_n634), .B2(KEYINPUT110), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT110), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n467), .B1(new_n468), .B2(new_n459), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n457), .A2(new_n464), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n703), .B1(new_n459), .B2(new_n704), .ZN(new_n705));
  AOI211_X1 g504(.A(new_n202), .B(new_n424), .C1(new_n468), .C2(new_n431), .ZN(new_n706));
  AOI21_X1  g505(.A(KEYINPUT84), .B1(new_n437), .B2(KEYINPUT35), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n705), .B1(new_n708), .B2(new_n432), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n702), .B1(new_n709), .B2(new_n633), .ZN(new_n710));
  NAND4_X1  g509(.A1(new_n701), .A2(new_n710), .A3(KEYINPUT51), .A4(new_n555), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n700), .A2(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n713), .A2(KEYINPUT111), .ZN(new_n714));
  INV_X1    g513(.A(new_n611), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n700), .B2(new_n712), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n714), .A2(new_n557), .A3(new_n715), .A4(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n693), .B1(new_n718), .B2(new_n641), .ZN(G1336gat));
  INV_X1    g518(.A(KEYINPUT52), .ZN(new_n720));
  OAI21_X1  g519(.A(G92gat), .B1(new_n692), .B2(new_n430), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n715), .A2(new_n264), .A3(new_n271), .ZN(new_n722));
  OAI211_X1 g521(.A(new_n720), .B(new_n721), .C1(new_n713), .C2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT113), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n699), .A2(new_n711), .A3(KEYINPUT112), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT112), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n726), .B(new_n694), .C1(new_n697), .C2(new_n698), .ZN(new_n727));
  INV_X1    g526(.A(new_n722), .ZN(new_n728));
  NAND3_X1  g527(.A1(new_n725), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n721), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n724), .B1(new_n730), .B2(KEYINPUT52), .ZN(new_n731));
  AOI211_X1 g530(.A(KEYINPUT113), .B(new_n720), .C1(new_n729), .C2(new_n721), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n723), .B1(new_n731), .B2(new_n732), .ZN(G1337gat));
  XNOR2_X1  g532(.A(KEYINPUT114), .B(G99gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n715), .A3(new_n717), .A4(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(new_n466), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n692), .A2(new_n626), .ZN(new_n737));
  OAI22_X1  g536(.A1(new_n735), .A2(new_n736), .B1(new_n737), .B2(new_n734), .ZN(G1338gat));
  INV_X1    g537(.A(G106gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n715), .A2(new_n739), .A3(new_n458), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n727), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(G106gat), .B1(new_n692), .B2(new_n459), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(KEYINPUT53), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT115), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT53), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n743), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g547(.A(new_n740), .B1(new_n699), .B2(new_n711), .ZN(new_n749));
  OR2_X1    g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n745), .A2(new_n746), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n747), .B1(new_n742), .B2(new_n743), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n748), .A2(new_n749), .ZN(new_n753));
  OAI21_X1  g552(.A(KEYINPUT115), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n754), .ZN(G1339gat));
  NOR2_X1   g554(.A1(new_n641), .A2(new_n271), .ZN(new_n756));
  INV_X1    g555(.A(new_n610), .ZN(new_n757));
  AND4_X1   g556(.A1(new_n696), .A2(new_n757), .A3(new_n579), .A4(new_n608), .ZN(new_n758));
  INV_X1    g557(.A(new_n555), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n605), .A2(new_n594), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT54), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n601), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n605), .B2(new_n594), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(new_n596), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT55), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OR2_X1    g566(.A1(new_n517), .A2(new_n518), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n507), .A2(new_n509), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n526), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(new_n522), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n770), .B1(new_n771), .B2(new_n527), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n762), .A2(new_n764), .A3(KEYINPUT55), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n767), .A2(new_n602), .A3(new_n772), .A4(new_n773), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n759), .B1(new_n774), .B2(new_n578), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n767), .A2(new_n529), .A3(new_n602), .A4(new_n773), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n772), .B1(new_n609), .B2(new_n610), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n776), .A2(new_n777), .A3(new_n633), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n758), .B1(new_n775), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(KEYINPUT116), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI211_X1 g580(.A(KEYINPUT116), .B(new_n758), .C1(new_n775), .C2(new_n778), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n431), .B(new_n756), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(G113gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n529), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n779), .B(new_n780), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n787), .A2(KEYINPUT117), .A3(new_n431), .A4(new_n756), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT117), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n783), .A2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n696), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n786), .B1(new_n791), .B2(new_n785), .ZN(G1340gat));
  INV_X1    g591(.A(G120gat), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n784), .A2(new_n793), .A3(new_n715), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n788), .A2(new_n790), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(new_n715), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT118), .B1(new_n796), .B2(G120gat), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT118), .ZN(new_n798));
  AOI211_X1 g597(.A(new_n798), .B(new_n793), .C1(new_n795), .C2(new_n715), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n794), .B1(new_n797), .B2(new_n799), .ZN(G1341gat));
  NAND3_X1  g599(.A1(new_n795), .A2(G127gat), .A3(new_n759), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(KEYINPUT119), .ZN(new_n802));
  INV_X1    g601(.A(G127gat), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n803), .B1(new_n783), .B2(new_n555), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT119), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n795), .A2(new_n805), .A3(G127gat), .A4(new_n759), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n802), .A2(new_n804), .A3(new_n806), .ZN(G1342gat));
  NOR3_X1   g606(.A1(new_n783), .A2(G134gat), .A3(new_n633), .ZN(new_n808));
  XNOR2_X1  g607(.A(new_n808), .B(KEYINPUT56), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n795), .A2(new_n578), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT120), .B1(new_n810), .B2(G134gat), .ZN(new_n811));
  INV_X1    g610(.A(KEYINPUT120), .ZN(new_n812));
  INV_X1    g611(.A(G134gat), .ZN(new_n813));
  AOI211_X1 g612(.A(new_n812), .B(new_n813), .C1(new_n795), .C2(new_n578), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n809), .B1(new_n811), .B2(new_n814), .ZN(G1343gat));
  NOR2_X1   g614(.A1(new_n627), .A2(new_n459), .ZN(new_n816));
  OR2_X1    g615(.A1(new_n816), .A2(KEYINPUT121), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n787), .A2(new_n756), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n816), .A2(KEYINPUT121), .ZN(new_n820));
  NAND4_X1  g619(.A1(new_n819), .A2(new_n289), .A3(new_n529), .A4(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n822));
  OAI211_X1 g621(.A(new_n822), .B(new_n458), .C1(new_n781), .C2(new_n782), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n756), .A2(new_n467), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  OAI21_X1  g624(.A(KEYINPUT57), .B1(new_n779), .B2(new_n459), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G141gat), .B1(new_n827), .B2(new_n696), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n821), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n821), .A2(new_n831), .A3(new_n828), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  NAND2_X1  g632(.A1(new_n291), .A2(new_n293), .ZN(new_n834));
  NAND4_X1  g633(.A1(new_n819), .A2(new_n834), .A3(new_n715), .A4(new_n820), .ZN(new_n835));
  INV_X1    g634(.A(new_n827), .ZN(new_n836));
  AOI211_X1 g635(.A(KEYINPUT59), .B(new_n834), .C1(new_n836), .C2(new_n715), .ZN(new_n837));
  XOR2_X1   g636(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n838));
  OAI211_X1 g637(.A(KEYINPUT57), .B(new_n458), .C1(new_n781), .C2(new_n782), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n822), .B1(new_n779), .B2(new_n459), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n841), .A2(new_n715), .A3(new_n825), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n838), .B1(new_n842), .B2(G148gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n835), .B1(new_n837), .B2(new_n843), .ZN(G1345gat));
  NOR2_X1   g643(.A1(new_n781), .A2(new_n782), .ZN(new_n845));
  INV_X1    g644(.A(new_n756), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n847), .A2(new_n759), .A3(new_n820), .A4(new_n817), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT123), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n819), .A2(KEYINPUT123), .A3(new_n759), .A4(new_n820), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n850), .A2(new_n851), .A3(new_n285), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n836), .A2(G155gat), .A3(new_n759), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n852), .A2(new_n853), .ZN(G1346gat));
  NOR3_X1   g653(.A1(new_n827), .A2(new_n286), .A3(new_n633), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n819), .A2(new_n578), .A3(new_n820), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n855), .B1(new_n286), .B2(new_n856), .ZN(G1347gat));
  NOR2_X1   g656(.A1(new_n614), .A2(new_n430), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n787), .A2(new_n431), .A3(new_n858), .ZN(new_n859));
  NOR3_X1   g658(.A1(new_n859), .A2(G169gat), .A3(new_n696), .ZN(new_n860));
  XNOR2_X1  g659(.A(new_n860), .B(KEYINPUT124), .ZN(new_n861));
  OAI21_X1  g660(.A(G169gat), .B1(new_n859), .B2(new_n696), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT125), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n861), .A2(new_n864), .ZN(G1348gat));
  NOR2_X1   g664(.A1(new_n859), .A2(new_n611), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(G176gat), .Z(G1349gat));
  INV_X1    g666(.A(G183gat), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n868), .B1(new_n859), .B2(new_n555), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n845), .A2(new_n368), .ZN(new_n870));
  INV_X1    g669(.A(new_n235), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n870), .A2(new_n759), .A3(new_n871), .A4(new_n858), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT60), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(KEYINPUT126), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n873), .A2(KEYINPUT126), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n875), .B(new_n876), .ZN(G1350gat));
  XNOR2_X1  g676(.A(KEYINPUT61), .B(G190gat), .ZN(new_n878));
  NAND2_X1  g677(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n859), .A2(new_n633), .ZN(new_n880));
  MUX2_X1   g679(.A(new_n878), .B(new_n879), .S(new_n880), .Z(G1351gat));
  NAND2_X1  g680(.A1(new_n816), .A2(new_n271), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT127), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n787), .A2(new_n883), .A3(new_n641), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(G197gat), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n885), .A2(new_n886), .A3(new_n529), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n626), .A2(new_n858), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n888), .B1(new_n839), .B2(new_n840), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n889), .A2(new_n529), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n887), .B1(new_n890), .B2(new_n886), .ZN(G1352gat));
  NOR3_X1   g690(.A1(new_n884), .A2(G204gat), .A3(new_n611), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n892), .A2(new_n893), .ZN(new_n895));
  INV_X1    g694(.A(G204gat), .ZN(new_n896));
  AOI211_X1 g695(.A(new_n611), .B(new_n888), .C1(new_n839), .C2(new_n840), .ZN(new_n897));
  OAI211_X1 g696(.A(new_n894), .B(new_n895), .C1(new_n896), .C2(new_n897), .ZN(G1353gat));
  NAND3_X1  g697(.A1(new_n885), .A2(new_n211), .A3(new_n759), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n889), .A2(new_n759), .ZN(new_n900));
  AND3_X1   g699(.A1(new_n900), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n901));
  AOI21_X1  g700(.A(KEYINPUT63), .B1(new_n900), .B2(G211gat), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(G1354gat));
  NAND3_X1  g702(.A1(new_n885), .A2(new_n212), .A3(new_n578), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n889), .A2(new_n578), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(new_n212), .ZN(G1355gat));
endmodule


