//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n204, new_n205, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1289, new_n1290,
    new_n1292, new_n1293, new_n1294, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370, new_n1371,
    new_n1372, new_n1373, new_n1374, new_n1375;
  NOR3_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .ZN(new_n201));
  XNOR2_X1  g0001(.A(new_n201), .B(KEYINPUT64), .ZN(new_n202));
  NOR2_X1   g0002(.A1(new_n202), .A2(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(new_n204));
  XNOR2_X1  g0004(.A(new_n204), .B(KEYINPUT65), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(KEYINPUT66), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n208), .ZN(new_n216));
  OAI21_X1  g0016(.A(G50), .B1(G58), .B2(G68), .ZN(new_n217));
  INV_X1    g0017(.A(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(new_n213), .A2(new_n214), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n219), .B1(new_n213), .B2(new_n214), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n221));
  INV_X1    g0021(.A(G68), .ZN(new_n222));
  INV_X1    g0022(.A(G238), .ZN(new_n223));
  INV_X1    g0023(.A(G87), .ZN(new_n224));
  INV_X1    g0024(.A(G250), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n210), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT1), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n220), .A2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G264), .B(G270), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n235), .B(KEYINPUT67), .Z(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G87), .B(G97), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT68), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G50), .B(G68), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G58), .B(G77), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND2_X1  g0050(.A1(new_n202), .A2(G20), .ZN(new_n251));
  INV_X1    g0051(.A(G150), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n208), .A2(G33), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI221_X1 g0056(.A(new_n251), .B1(new_n252), .B2(new_n254), .C1(new_n255), .C2(new_n256), .ZN(new_n257));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(new_n215), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g0060(.A1(new_n258), .A2(new_n215), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n207), .A2(G13), .A3(G20), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(G50), .B1(new_n208), .B2(G1), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n263), .A2(new_n264), .B1(G50), .B2(new_n262), .ZN(new_n265));
  XOR2_X1   g0065(.A(new_n265), .B(KEYINPUT70), .Z(new_n266));
  NAND2_X1  g0066(.A1(new_n260), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  INV_X1    g0068(.A(G1698), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n268), .A2(G222), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G77), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n268), .A2(G1698), .ZN(new_n272));
  INV_X1    g0072(.A(G223), .ZN(new_n273));
  OAI221_X1 g0073(.A(new_n270), .B1(new_n271), .B2(new_n268), .C1(new_n272), .C2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(G33), .A2(G41), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n275), .A2(G1), .A3(G13), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n274), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G179), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT69), .A2(G41), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT69), .A2(G41), .ZN(new_n281));
  NOR3_X1   g0081(.A1(new_n280), .A2(new_n281), .A3(G45), .ZN(new_n282));
  INV_X1    g0082(.A(G274), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G1), .ZN(new_n284));
  INV_X1    g0084(.A(new_n284), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n287));
  AND2_X1   g0087(.A1(new_n276), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n286), .B1(G226), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n278), .A2(new_n279), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n278), .A2(new_n289), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n267), .A2(new_n290), .A3(new_n293), .ZN(new_n294));
  INV_X1    g0094(.A(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT75), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n296), .B1(new_n291), .B2(G200), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  OAI221_X1 g0099(.A(new_n297), .B1(new_n298), .B2(new_n291), .C1(new_n267), .C2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n267), .A2(new_n299), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(KEYINPUT74), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT74), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n267), .A2(new_n304), .A3(new_n299), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n301), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n304), .B1(new_n267), .B2(new_n299), .ZN(new_n309));
  AOI211_X1 g0109(.A(KEYINPUT74), .B(KEYINPUT9), .C1(new_n260), .C2(new_n266), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT10), .B1(new_n311), .B2(new_n300), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n295), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT18), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n256), .B1(new_n207), .B2(G20), .ZN(new_n315));
  INV_X1    g0115(.A(new_n262), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n316), .A2(new_n259), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n315), .A2(new_n317), .B1(new_n316), .B2(new_n256), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(KEYINPUT3), .A2(G33), .ZN(new_n320));
  NOR2_X1   g0120(.A1(KEYINPUT3), .A2(G33), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(KEYINPUT7), .B1(new_n322), .B2(new_n208), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT3), .ZN(new_n324));
  INV_X1    g0124(.A(G33), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(KEYINPUT3), .A2(G33), .ZN(new_n327));
  NAND4_X1  g0127(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  OAI21_X1  g0129(.A(G68), .B1(new_n323), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(G58), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(new_n222), .ZN(new_n332));
  NOR2_X1   g0132(.A1(G58), .A2(G68), .ZN(new_n333));
  OAI21_X1  g0133(.A(G20), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n253), .A2(G159), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n334), .A2(KEYINPUT16), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n261), .B1(new_n330), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT16), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n326), .A2(new_n208), .A3(new_n327), .ZN(new_n340));
  INV_X1    g0140(.A(KEYINPUT7), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n222), .B1(new_n342), .B2(new_n328), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n334), .A2(new_n335), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n339), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n319), .B1(new_n338), .B2(new_n345), .ZN(new_n346));
  OAI211_X1 g0146(.A(G223), .B(new_n269), .C1(new_n320), .C2(new_n321), .ZN(new_n347));
  OAI211_X1 g0147(.A(G226), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n348));
  NAND2_X1  g0148(.A1(G33), .A2(G87), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n347), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n277), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT69), .ZN(new_n352));
  INV_X1    g0152(.A(G41), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(G45), .ZN(new_n355));
  NAND2_X1  g0155(.A1(KEYINPUT69), .A2(G41), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI22_X1  g0157(.A1(new_n288), .A2(G232), .B1(new_n357), .B2(new_n284), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n351), .A2(new_n279), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n276), .A2(new_n287), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n282), .A2(new_n285), .B1(new_n360), .B2(new_n238), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n361), .B1(new_n277), .B2(new_n350), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n359), .B1(new_n362), .B2(G169), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n314), .B1(new_n346), .B2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(KEYINPUT82), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n351), .A2(new_n279), .A3(new_n358), .ZN(new_n366));
  AOI21_X1  g0166(.A(G169), .B1(new_n351), .B2(new_n358), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n344), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT16), .B1(new_n330), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n259), .B1(new_n343), .B2(new_n336), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n318), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n368), .A2(new_n372), .A3(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT82), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n375), .B(new_n314), .C1(new_n346), .C2(new_n363), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT81), .ZN(new_n377));
  NAND4_X1  g0177(.A1(new_n368), .A2(new_n372), .A3(new_n377), .A4(KEYINPUT18), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n365), .A2(new_n374), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n351), .A2(new_n358), .ZN(new_n380));
  OAI21_X1  g0180(.A(KEYINPUT83), .B1(new_n380), .B2(G190), .ZN(new_n381));
  INV_X1    g0181(.A(G200), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT83), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n351), .A2(new_n358), .A3(new_n384), .A4(new_n298), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AND3_X1   g0186(.A1(new_n386), .A2(KEYINPUT17), .A3(new_n346), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT17), .B1(new_n386), .B2(new_n346), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n379), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n313), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT73), .ZN(new_n392));
  INV_X1    g0192(.A(new_n256), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n253), .B1(G20), .B2(G77), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT15), .B(G87), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(new_n255), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n396), .A2(KEYINPUT71), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n394), .A2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT71), .B1(new_n396), .B2(new_n397), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n259), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT72), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n402), .B1(new_n262), .B2(G77), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n316), .A2(KEYINPUT72), .A3(new_n271), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n271), .B1(new_n207), .B2(G20), .ZN(new_n405));
  AOI22_X1  g0205(.A1(new_n403), .A2(new_n404), .B1(new_n317), .B2(new_n405), .ZN(new_n406));
  AND2_X1   g0206(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n268), .A2(G232), .A3(new_n269), .ZN(new_n408));
  INV_X1    g0208(.A(G107), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n409), .B2(new_n268), .C1(new_n272), .C2(new_n223), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n277), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n286), .B1(G244), .B2(new_n288), .ZN(new_n412));
  AOI21_X1  g0212(.A(G169), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n392), .B1(new_n407), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n401), .A2(new_n406), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n411), .A2(new_n412), .ZN(new_n416));
  OAI211_X1 g0216(.A(KEYINPUT73), .B(new_n415), .C1(new_n416), .C2(G169), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n279), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n414), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(G190), .ZN(new_n420));
  OAI211_X1 g0220(.A(new_n420), .B(new_n407), .C1(new_n382), .C2(new_n416), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  XNOR2_X1  g0222(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n238), .A2(G1698), .ZN(new_n425));
  OAI211_X1 g0225(.A(new_n268), .B(new_n425), .C1(G226), .C2(G1698), .ZN(new_n426));
  NAND2_X1  g0226(.A1(G33), .A2(G97), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n276), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n428), .ZN(new_n429));
  OAI22_X1  g0229(.A1(new_n282), .A2(new_n285), .B1(new_n360), .B2(new_n223), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n424), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n428), .A2(new_n430), .A3(new_n423), .ZN(new_n433));
  OAI21_X1  g0233(.A(G169), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(KEYINPUT14), .ZN(new_n435));
  OAI21_X1  g0235(.A(KEYINPUT13), .B1(new_n428), .B2(new_n430), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT77), .ZN(new_n437));
  INV_X1    g0237(.A(new_n433), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT77), .ZN(new_n439));
  OAI211_X1 g0239(.A(new_n439), .B(KEYINPUT13), .C1(new_n428), .C2(new_n430), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n437), .A2(new_n438), .A3(G179), .A4(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT14), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n442), .B(G169), .C1(new_n432), .C2(new_n433), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n435), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  AOI22_X1  g0244(.A1(new_n397), .A2(G77), .B1(G20), .B2(new_n222), .ZN(new_n445));
  INV_X1    g0245(.A(G50), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n445), .B1(new_n446), .B2(new_n254), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n447), .A2(new_n259), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT11), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n447), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT78), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n450), .A2(KEYINPUT78), .A3(new_n451), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT79), .B1(new_n262), .B2(G68), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT12), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n222), .B1(new_n207), .B2(G20), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n317), .B2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n454), .A2(new_n455), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n444), .A2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n460), .ZN(new_n462));
  NAND4_X1  g0262(.A1(new_n437), .A2(new_n438), .A3(G190), .A4(new_n440), .ZN(new_n463));
  OAI21_X1  g0263(.A(G200), .B1(new_n432), .B2(new_n433), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n461), .A2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT80), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n422), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(new_n467), .B2(new_n466), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n391), .A2(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n316), .A2(KEYINPUT25), .A3(new_n409), .ZN(new_n472));
  INV_X1    g0272(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(KEYINPUT25), .B1(new_n316), .B2(new_n409), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n261), .B(new_n262), .C1(G1), .C2(new_n325), .ZN(new_n475));
  OAI22_X1  g0275(.A1(new_n473), .A2(new_n474), .B1(new_n475), .B2(new_n409), .ZN(new_n476));
  INV_X1    g0276(.A(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT90), .ZN(new_n478));
  OAI211_X1 g0278(.A(new_n208), .B(G87), .C1(new_n320), .C2(new_n321), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT22), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT22), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n268), .A2(new_n481), .A3(new_n208), .A4(G87), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G116), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n484), .A2(G20), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT23), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n486), .B1(new_n208), .B2(G107), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n409), .A2(KEYINPUT23), .A3(G20), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n485), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n483), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT24), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT24), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n483), .A2(new_n492), .A3(new_n489), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n478), .B1(new_n494), .B2(new_n259), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n483), .A2(new_n492), .A3(new_n489), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n492), .B1(new_n483), .B2(new_n489), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n478), .B(new_n259), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(new_n498), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n477), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  OAI211_X1 g0300(.A(G250), .B(new_n269), .C1(new_n320), .C2(new_n321), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT92), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n268), .A2(KEYINPUT92), .A3(G250), .A4(new_n269), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT91), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n268), .A2(new_n505), .A3(G257), .A4(G1698), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  OAI211_X1 g0307(.A(G257), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n508));
  XNOR2_X1  g0308(.A(KEYINPUT93), .B(G294), .ZN(new_n509));
  AOI22_X1  g0309(.A1(new_n508), .A2(KEYINPUT91), .B1(G33), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n276), .B1(new_n507), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT5), .B1(new_n354), .B2(new_n356), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n355), .A2(G1), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g0314(.A(KEYINPUT86), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT5), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n280), .B2(new_n281), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT86), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(new_n518), .A3(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n353), .A2(KEYINPUT5), .ZN(new_n520));
  AND3_X1   g0320(.A1(new_n276), .A2(G274), .A3(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n515), .A2(new_n519), .A3(new_n521), .ZN(new_n522));
  NAND3_X1  g0322(.A1(new_n517), .A2(new_n513), .A3(new_n520), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G264), .A3(new_n276), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(G169), .B1(new_n511), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(KEYINPUT94), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT94), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n523), .A2(new_n528), .A3(G264), .A4(new_n276), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n510), .A2(new_n504), .A3(new_n506), .A4(new_n503), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n277), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n530), .A2(new_n532), .A3(G179), .A4(new_n522), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n500), .A2(KEYINPUT95), .A3(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT95), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n259), .B1(new_n496), .B2(new_n497), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(KEYINPUT90), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n476), .B1(new_n538), .B2(new_n498), .ZN(new_n539));
  AND2_X1   g0339(.A1(new_n526), .A2(new_n533), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n536), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n530), .A2(new_n532), .A3(new_n522), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n382), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n532), .A2(new_n522), .A3(new_n524), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n543), .B1(G190), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n539), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n535), .A2(new_n541), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(G33), .A2(G283), .ZN(new_n548));
  INV_X1    g0348(.A(G97), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n548), .B(new_n208), .C1(G33), .C2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(G116), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G20), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n259), .A3(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT20), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(KEYINPUT20), .A3(new_n259), .A4(new_n552), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NOR2_X1   g0357(.A1(new_n262), .A2(G116), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n325), .A2(G1), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n316), .A2(new_n259), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n558), .B1(new_n560), .B2(G116), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n557), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(new_n562), .ZN(new_n563));
  OAI211_X1 g0363(.A(G257), .B(new_n269), .C1(new_n320), .C2(new_n321), .ZN(new_n564));
  OAI211_X1 g0364(.A(G264), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n326), .A2(G303), .A3(new_n327), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n277), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n523), .A2(G270), .A3(new_n276), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n522), .A2(new_n568), .A3(G190), .A4(new_n569), .ZN(new_n570));
  AND3_X1   g0370(.A1(new_n522), .A2(new_n568), .A3(new_n569), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n563), .B(new_n570), .C1(new_n571), .C2(new_n382), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(G179), .A3(new_n562), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n292), .B1(new_n557), .B2(new_n561), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT21), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n522), .A2(new_n568), .A3(new_n569), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n575), .B1(new_n574), .B2(new_n576), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n572), .B(new_n573), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  INV_X1    g0380(.A(KEYINPUT89), .ZN(new_n581));
  OAI211_X1 g0381(.A(G244), .B(G1698), .C1(new_n320), .C2(new_n321), .ZN(new_n582));
  OAI211_X1 g0382(.A(G238), .B(new_n269), .C1(new_n320), .C2(new_n321), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n582), .A2(new_n583), .A3(new_n484), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n277), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n225), .B1(new_n355), .B2(G1), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n207), .A2(new_n283), .A3(G45), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n276), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n292), .B1(new_n585), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n279), .B(new_n588), .C1(new_n584), .C2(new_n277), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n581), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n585), .A2(G179), .A3(new_n589), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n588), .B1(new_n584), .B2(new_n277), .ZN(new_n594));
  OAI211_X1 g0394(.A(new_n593), .B(KEYINPUT89), .C1(new_n292), .C2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n268), .A2(new_n208), .A3(G68), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT19), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n208), .B1(new_n427), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n224), .A2(new_n549), .A3(new_n409), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n597), .B1(new_n255), .B2(new_n549), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n596), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  AOI22_X1  g0402(.A1(new_n602), .A2(new_n259), .B1(new_n316), .B2(new_n395), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n603), .B1(new_n475), .B2(new_n395), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n592), .A2(new_n595), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n560), .A2(G87), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n594), .A2(G190), .ZN(new_n608));
  OR2_X1    g0408(.A1(new_n594), .A2(new_n382), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n605), .A2(new_n610), .ZN(new_n611));
  NOR2_X1   g0411(.A1(new_n580), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT87), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n523), .A2(G257), .A3(new_n276), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n522), .A2(new_n614), .ZN(new_n615));
  OAI211_X1 g0415(.A(G244), .B(new_n269), .C1(new_n320), .C2(new_n321), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT4), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n548), .ZN(new_n619));
  NAND2_X1  g0419(.A1(G250), .A2(G1698), .ZN(new_n620));
  NAND2_X1  g0420(.A1(KEYINPUT4), .A2(G244), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n620), .B1(new_n621), .B2(G1698), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n619), .B1(new_n268), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n624), .A2(KEYINPUT85), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n618), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n625), .A2(new_n277), .A3(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n615), .A2(new_n628), .A3(G190), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n316), .A2(new_n549), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n630), .B1(new_n475), .B2(new_n549), .ZN(new_n631));
  OAI21_X1  g0431(.A(G107), .B1(new_n323), .B2(new_n329), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n253), .A2(G77), .ZN(new_n633));
  AND2_X1   g0433(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n634));
  NOR2_X1   g0434(.A1(KEYINPUT84), .A2(KEYINPUT6), .ZN(new_n635));
  OAI22_X1  g0435(.A1(new_n634), .A2(new_n635), .B1(new_n549), .B2(G107), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  XNOR2_X1  g0437(.A(G97), .B(G107), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n636), .B(G20), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n632), .A2(new_n633), .A3(new_n639), .ZN(new_n640));
  AOI21_X1  g0440(.A(new_n631), .B1(new_n640), .B2(new_n259), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n629), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n382), .B1(new_n615), .B2(new_n628), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n613), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n615), .A2(new_n628), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(G200), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n646), .A2(KEYINPUT87), .A3(new_n641), .A4(new_n629), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n641), .B1(new_n645), .B2(new_n292), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n522), .A2(new_n614), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n276), .B1(new_n624), .B2(KEYINPUT85), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n627), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(KEYINPUT88), .A3(new_n279), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n615), .A2(new_n628), .A3(new_n279), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT88), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n649), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g0457(.A1(new_n612), .A2(new_n648), .A3(new_n657), .ZN(new_n658));
  NOR3_X1   g0458(.A1(new_n471), .A2(new_n547), .A3(new_n658), .ZN(G372));
  NAND2_X1  g0459(.A1(new_n364), .A2(new_n373), .ZN(new_n660));
  INV_X1    g0460(.A(new_n419), .ZN(new_n661));
  AOI22_X1  g0461(.A1(new_n661), .A2(new_n465), .B1(new_n460), .B2(new_n444), .ZN(new_n662));
  INV_X1    g0462(.A(new_n389), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n660), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n308), .A2(new_n312), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n295), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  AND2_X1   g0466(.A1(new_n649), .A2(new_n656), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT26), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n593), .B1(new_n292), .B2(new_n594), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n604), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n610), .A2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n667), .A2(new_n668), .A3(new_n653), .A4(new_n672), .ZN(new_n673));
  OAI21_X1  g0473(.A(KEYINPUT26), .B1(new_n657), .B2(new_n611), .ZN(new_n674));
  AND3_X1   g0474(.A1(new_n673), .A2(new_n670), .A3(new_n674), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n671), .B1(new_n545), .B2(new_n539), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n563), .A2(new_n576), .A3(new_n279), .ZN(new_n677));
  INV_X1    g0477(.A(new_n579), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n577), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n539), .B2(new_n540), .ZN(new_n680));
  NAND4_X1  g0480(.A1(new_n676), .A2(new_n680), .A3(new_n648), .A4(new_n657), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n666), .B1(new_n471), .B2(new_n683), .ZN(G369));
  NOR2_X1   g0484(.A1(new_n539), .A2(new_n540), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(KEYINPUT27), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n687), .A2(G213), .A3(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(G343), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n685), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT96), .ZN(new_n693));
  AND3_X1   g0493(.A1(new_n535), .A2(new_n541), .A3(new_n546), .ZN(new_n694));
  INV_X1    g0494(.A(new_n691), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n694), .B1(new_n539), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n679), .A2(new_n691), .ZN(new_n698));
  AOI22_X1  g0498(.A1(new_n697), .A2(new_n698), .B1(new_n685), .B2(new_n695), .ZN(new_n699));
  INV_X1    g0499(.A(new_n679), .ZN(new_n700));
  NOR2_X1   g0500(.A1(new_n563), .A2(new_n695), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n580), .B2(new_n701), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G330), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n697), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n699), .A2(new_n706), .ZN(G399));
  NOR2_X1   g0507(.A1(new_n280), .A2(new_n281), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n211), .A2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n599), .A2(G116), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n711), .B1(new_n217), .B2(new_n709), .ZN(new_n712));
  XNOR2_X1  g0512(.A(new_n712), .B(KEYINPUT28), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n612), .A2(new_n648), .A3(new_n657), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n694), .A2(new_n714), .A3(new_n695), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT30), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n571), .A2(new_n530), .A3(new_n532), .A4(new_n591), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n645), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n576), .A2(new_n593), .ZN(new_n719));
  AOI22_X1  g0519(.A1(new_n527), .A2(new_n529), .B1(new_n531), .B2(new_n277), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n652), .A2(new_n719), .A3(new_n720), .A4(KEYINPUT30), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n594), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n542), .A2(new_n645), .A3(new_n576), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n718), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n691), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n724), .B2(new_n691), .ZN(new_n727));
  OAI21_X1  g0527(.A(KEYINPUT97), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n691), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT31), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g0531(.A(KEYINPUT97), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n725), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n715), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  AND3_X1   g0534(.A1(new_n734), .A2(KEYINPUT98), .A3(G330), .ZN(new_n735));
  AOI21_X1  g0535(.A(KEYINPUT98), .B1(new_n734), .B2(G330), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n691), .B1(new_n675), .B2(new_n681), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n648), .A2(new_n657), .ZN(new_n740));
  INV_X1    g0540(.A(KEYINPUT99), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n648), .A2(KEYINPUT99), .A3(new_n657), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n535), .A2(new_n541), .A3(new_n679), .ZN(new_n744));
  NAND4_X1  g0544(.A1(new_n742), .A2(new_n676), .A3(new_n743), .A4(new_n744), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n657), .A2(new_n611), .A3(KEYINPUT26), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT26), .B1(new_n657), .B2(new_n671), .ZN(new_n747));
  AND3_X1   g0547(.A1(new_n746), .A2(new_n670), .A3(new_n747), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n691), .B1(new_n745), .B2(new_n748), .ZN(new_n749));
  MUX2_X1   g0549(.A(new_n739), .B(new_n749), .S(KEYINPUT29), .Z(new_n750));
  AND2_X1   g0550(.A1(new_n737), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n713), .B1(new_n751), .B2(G1), .ZN(G364));
  INV_X1    g0552(.A(new_n709), .ZN(new_n753));
  INV_X1    g0553(.A(G13), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n207), .B1(new_n755), .B2(G45), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n705), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G330), .B2(new_n703), .ZN(new_n760));
  INV_X1    g0560(.A(new_n211), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n761), .A2(new_n322), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G355), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n763), .B1(G116), .B2(new_n211), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n211), .A2(new_n322), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT100), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n767), .B1(new_n355), .B2(new_n218), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n249), .A2(G45), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n764), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G13), .A2(G33), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n772), .A2(G20), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n215), .B1(G20), .B2(new_n292), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(new_n775), .B(KEYINPUT101), .Z(new_n776));
  OAI21_X1  g0576(.A(new_n758), .B1(new_n770), .B2(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n298), .A2(G179), .A3(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n208), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n208), .A2(new_n279), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(G200), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n782), .A2(new_n298), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G97), .A2(new_n780), .B1(new_n783), .B2(G50), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n268), .B1(new_n786), .B2(new_n271), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n781), .A2(G190), .A3(new_n382), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n787), .B1(G58), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n208), .A2(G179), .ZN(new_n791));
  NAND3_X1  g0591(.A1(new_n791), .A2(G190), .A3(G200), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G87), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n791), .A2(new_n785), .ZN(new_n795));
  INV_X1    g0595(.A(G159), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT32), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND4_X1  g0599(.A1(new_n784), .A2(new_n790), .A3(new_n794), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n782), .A2(G190), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n791), .A2(new_n298), .A3(G200), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n801), .A2(G68), .B1(new_n803), .B2(G107), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n798), .B2(new_n797), .ZN(new_n805));
  INV_X1    g0605(.A(G317), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(KEYINPUT33), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n801), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(G303), .ZN(new_n810));
  INV_X1    g0610(.A(new_n509), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n809), .B1(new_n810), .B2(new_n792), .C1(new_n811), .C2(new_n779), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n783), .A2(G326), .B1(new_n803), .B2(G283), .ZN(new_n813));
  INV_X1    g0613(.A(new_n795), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n789), .A2(G322), .B1(new_n814), .B2(G329), .ZN(new_n815));
  INV_X1    g0615(.A(new_n786), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n268), .B1(new_n816), .B2(G311), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n813), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n800), .A2(new_n805), .B1(new_n812), .B2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT102), .ZN(new_n820));
  OR2_X1    g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n774), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n822), .B1(new_n819), .B2(new_n820), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n777), .B1(new_n821), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n773), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n703), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n760), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  OAI211_X1 g0628(.A(new_n419), .B(new_n421), .C1(new_n407), .C2(new_n695), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n407), .A2(new_n695), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n414), .A2(new_n417), .A3(new_n830), .A4(new_n418), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n829), .A2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(new_n681), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n673), .A2(new_n670), .A3(new_n674), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n695), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n832), .A2(KEYINPUT104), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT104), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n829), .A2(new_n837), .A3(new_n831), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n835), .B1(new_n738), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n758), .B1(new_n737), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n841), .B1(new_n737), .B2(new_n840), .ZN(new_n842));
  INV_X1    g0642(.A(new_n758), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n789), .A2(G143), .B1(new_n816), .B2(G159), .ZN(new_n844));
  INV_X1    g0644(.A(new_n801), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(new_n783), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n844), .B1(new_n845), .B2(new_n252), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT34), .ZN(new_n849));
  AND2_X1   g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n803), .A2(G68), .ZN(new_n851));
  INV_X1    g0651(.A(G132), .ZN(new_n852));
  OAI211_X1 g0652(.A(new_n851), .B(new_n268), .C1(new_n852), .C2(new_n795), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n779), .A2(new_n331), .B1(new_n792), .B2(new_n446), .ZN(new_n854));
  NOR3_X1   g0654(.A1(new_n850), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n855), .B1(new_n849), .B2(new_n848), .ZN(new_n856));
  OAI22_X1  g0656(.A1(new_n847), .A2(new_n810), .B1(new_n792), .B2(new_n409), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n857), .B1(G87), .B2(new_n803), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n268), .B1(new_n789), .B2(G294), .ZN(new_n859));
  AOI22_X1  g0659(.A1(G116), .A2(new_n816), .B1(new_n814), .B2(G311), .ZN(new_n860));
  AOI22_X1  g0660(.A1(G97), .A2(new_n780), .B1(new_n801), .B2(G283), .ZN(new_n861));
  NAND4_X1  g0661(.A1(new_n858), .A2(new_n859), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n822), .B1(new_n856), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n774), .A2(new_n771), .ZN(new_n864));
  AOI211_X1 g0664(.A(new_n843), .B(new_n863), .C1(new_n271), .C2(new_n864), .ZN(new_n865));
  XOR2_X1   g0665(.A(new_n865), .B(KEYINPUT103), .Z(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n772), .B2(new_n832), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n842), .A2(new_n867), .ZN(G384));
  NOR2_X1   g0668(.A1(new_n755), .A2(new_n207), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT105), .ZN(new_n870));
  INV_X1    g0670(.A(new_n689), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n372), .A2(new_n871), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n870), .B1(new_n390), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n386), .A2(new_n346), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n372), .B1(new_n368), .B2(new_n871), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g0676(.A1(new_n876), .A2(KEYINPUT37), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT37), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n872), .B1(new_n379), .B2(new_n389), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n880), .B1(new_n881), .B2(KEYINPUT105), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n873), .A2(new_n882), .A3(KEYINPUT38), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT38), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n879), .A2(KEYINPUT106), .ZN(new_n885));
  XNOR2_X1  g0685(.A(new_n876), .B(KEYINPUT37), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(KEYINPUT106), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n872), .B1(new_n389), .B2(new_n660), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n887), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n461), .A2(new_n691), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n379), .A2(new_n389), .ZN(new_n894));
  INV_X1    g0694(.A(new_n872), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(KEYINPUT105), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n886), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n881), .A2(KEYINPUT105), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n884), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n899), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n892), .A2(new_n893), .A3(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT107), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n660), .A2(new_n871), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n899), .A2(new_n883), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n460), .A2(new_n691), .ZN(new_n905));
  AND3_X1   g0705(.A1(new_n461), .A2(new_n465), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n905), .B1(new_n461), .B2(new_n465), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g0708(.A1(new_n419), .A2(new_n691), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n908), .B1(new_n835), .B2(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n903), .B1(new_n904), .B2(new_n911), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n901), .A2(new_n902), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n902), .B1(new_n901), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n666), .B1(new_n750), .B2(new_n471), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n915), .B(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(G330), .ZN(new_n918));
  INV_X1    g0718(.A(new_n905), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n466), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n461), .A2(new_n465), .A3(new_n905), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n920), .A2(new_n921), .B1(new_n829), .B2(new_n831), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n652), .A2(new_n720), .A3(new_n719), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n722), .A2(new_n576), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n652), .A2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n716), .A2(new_n923), .B1(new_n925), .B2(new_n542), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n695), .B1(new_n926), .B2(new_n721), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT108), .B1(new_n927), .B2(KEYINPUT31), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT108), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n727), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n725), .A3(new_n930), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n547), .A2(new_n658), .A3(new_n691), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n922), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(new_n883), .B2(new_n899), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT109), .B1(new_n934), .B2(KEYINPUT40), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n832), .B1(new_n906), .B2(new_n907), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n727), .A2(new_n929), .ZN(new_n937));
  AOI211_X1 g0737(.A(KEYINPUT108), .B(KEYINPUT31), .C1(new_n724), .C2(new_n691), .ZN(new_n938));
  NOR3_X1   g0738(.A1(new_n937), .A2(new_n938), .A3(new_n726), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n936), .B1(new_n939), .B2(new_n715), .ZN(new_n940));
  NOR3_X1   g0740(.A1(new_n897), .A2(new_n884), .A3(new_n898), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT38), .B1(new_n873), .B2(new_n882), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT109), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT40), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI211_X1 g0746(.A(new_n922), .B(KEYINPUT40), .C1(new_n931), .C2(new_n932), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI22_X1  g0748(.A1(new_n935), .A2(new_n946), .B1(new_n890), .B2(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n931), .A2(new_n932), .ZN(new_n950));
  NOR2_X1   g0750(.A1(new_n471), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n918), .B1(new_n949), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n952), .B1(new_n949), .B2(new_n951), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n869), .B1(new_n917), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n953), .B2(new_n917), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT35), .ZN(new_n957));
  OAI211_X1 g0757(.A(G116), .B(new_n216), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n957), .B2(new_n956), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT36), .Z(new_n960));
  NOR3_X1   g0760(.A1(new_n332), .A2(new_n217), .A3(new_n271), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n222), .A2(G50), .ZN(new_n962));
  OAI211_X1 g0762(.A(G1), .B(new_n754), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n955), .A2(new_n960), .A3(new_n963), .ZN(G367));
  NAND2_X1  g0764(.A1(new_n697), .A2(new_n698), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT42), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n641), .A2(new_n695), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n742), .A2(new_n743), .A3(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n667), .A2(new_n653), .A3(new_n691), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  NOR3_X1   g0772(.A1(new_n965), .A2(new_n966), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n698), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n974), .B1(new_n693), .B2(new_n696), .ZN(new_n975));
  AOI21_X1  g0775(.A(KEYINPUT42), .B1(new_n975), .B2(new_n971), .ZN(new_n976));
  OR2_X1    g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n535), .A2(new_n541), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n742), .A2(new_n978), .A3(new_n743), .A4(new_n968), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n979), .A2(KEYINPUT110), .A3(new_n657), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n980), .A2(new_n695), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT110), .B1(new_n979), .B2(new_n657), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n607), .A2(new_n695), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n984), .A2(new_n669), .A3(new_n604), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n671), .B2(new_n984), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n987));
  NAND4_X1  g0787(.A1(new_n977), .A2(new_n983), .A3(KEYINPUT111), .A4(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT111), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n983), .B1(new_n973), .B2(new_n976), .ZN(new_n990));
  INV_X1    g0790(.A(new_n987), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n989), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n986), .A2(KEYINPUT43), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n990), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n706), .B2(new_n972), .ZN(new_n997));
  INV_X1    g0797(.A(new_n706), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n993), .A2(new_n998), .A3(new_n971), .A4(new_n995), .ZN(new_n999));
  XNOR2_X1  g0799(.A(new_n709), .B(KEYINPUT41), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n685), .A2(new_n695), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n965), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT44), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n971), .B1(KEYINPUT112), .B2(new_n1003), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1002), .A2(new_n1005), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1003), .A2(KEYINPUT112), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n972), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1004), .B1(new_n699), .B2(new_n1009), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT45), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1002), .B2(new_n972), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n699), .A2(KEYINPUT45), .A3(new_n971), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1011), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1016), .A2(new_n998), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n697), .A2(new_n698), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1018), .A2(new_n975), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(new_n704), .ZN(new_n1020));
  AND2_X1   g0820(.A1(new_n1020), .A2(new_n751), .ZN(new_n1021));
  NAND3_X1  g0821(.A1(new_n1011), .A2(new_n1015), .A3(new_n706), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1017), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1000), .B1(new_n1023), .B2(new_n751), .ZN(new_n1024));
  OAI211_X1 g0824(.A(new_n997), .B(new_n999), .C1(new_n1024), .C2(new_n757), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n776), .B1(new_n761), .B2(new_n396), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n766), .A2(new_n235), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n843), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n803), .A2(G77), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n268), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT113), .ZN(new_n1031));
  OAI22_X1  g0831(.A1(new_n788), .A2(new_n252), .B1(new_n786), .B2(new_n446), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1032), .B1(G137), .B2(new_n814), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n801), .A2(G159), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n780), .A2(G68), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n783), .A2(G143), .B1(new_n793), .B2(G58), .ZN(new_n1036));
  NAND4_X1  g0836(.A1(new_n1033), .A2(new_n1034), .A3(new_n1035), .A4(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n801), .A2(new_n509), .B1(new_n803), .B2(G97), .ZN(new_n1038));
  INV_X1    g0838(.A(G311), .ZN(new_n1039));
  OAI221_X1 g0839(.A(new_n1038), .B1(new_n409), .B2(new_n779), .C1(new_n1039), .C2(new_n847), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n789), .A2(G303), .B1(new_n814), .B2(G317), .ZN(new_n1041));
  INV_X1    g0841(.A(KEYINPUT46), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n792), .B2(new_n551), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n793), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n268), .B1(new_n816), .B2(G283), .ZN(new_n1045));
  NAND4_X1  g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .A4(new_n1045), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n1031), .A2(new_n1037), .B1(new_n1040), .B2(new_n1046), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT47), .Z(new_n1048));
  OAI221_X1 g0848(.A(new_n1028), .B1(new_n825), .B2(new_n986), .C1(new_n1048), .C2(new_n822), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1025), .A2(new_n1049), .ZN(G387));
  NAND2_X1  g0850(.A1(new_n1020), .A2(new_n757), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n393), .A2(new_n446), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT50), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n710), .ZN(new_n1055));
  AOI211_X1 g0855(.A(G45), .B(new_n1055), .C1(G68), .C2(G77), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n767), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OR2_X1    g0857(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1057), .A2(KEYINPUT114), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1058), .B(new_n1059), .C1(new_n355), .C2(new_n241), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n762), .A2(new_n1055), .B1(new_n409), .B2(new_n761), .ZN(new_n1061));
  AND2_X1   g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n776), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1062), .A2(KEYINPUT115), .ZN(new_n1065));
  NAND3_X1  g0865(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n786), .A2(new_n222), .B1(new_n795), .B2(new_n252), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n322), .B(new_n1067), .C1(G50), .C2(new_n789), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n793), .A2(G77), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(new_n396), .A2(new_n780), .B1(new_n801), .B2(new_n393), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n783), .A2(G159), .B1(new_n803), .B2(G97), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1068), .A2(new_n1069), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n268), .B1(new_n814), .B2(G326), .ZN(new_n1073));
  INV_X1    g0873(.A(G283), .ZN(new_n1074));
  OAI22_X1  g0874(.A1(new_n779), .A2(new_n1074), .B1(new_n811), .B2(new_n792), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n789), .A2(G317), .B1(new_n816), .B2(G303), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n783), .A2(G322), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n1076), .B(new_n1077), .C1(new_n1039), .C2(new_n845), .ZN(new_n1078));
  INV_X1    g0878(.A(KEYINPUT48), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1075), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1080), .B1(new_n1079), .B2(new_n1078), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT49), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1073), .B1(new_n551), .B2(new_n802), .C1(new_n1081), .C2(new_n1082), .ZN(new_n1083));
  AND2_X1   g0883(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1072), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n843), .B1(new_n1085), .B2(new_n774), .ZN(new_n1086));
  OAI211_X1 g0886(.A(new_n1066), .B(new_n1086), .C1(new_n697), .C2(new_n825), .ZN(new_n1087));
  OR2_X1    g0887(.A1(new_n1021), .A2(new_n709), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n1020), .A2(new_n751), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n1051), .B(new_n1087), .C1(new_n1088), .C2(new_n1089), .ZN(G393));
  AND3_X1   g0890(.A1(new_n1011), .A2(new_n706), .A3(new_n1015), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n706), .B1(new_n1011), .B2(new_n1015), .ZN(new_n1092));
  OAI21_X1  g0892(.A(KEYINPUT116), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  INV_X1    g0893(.A(KEYINPUT116), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1022), .A2(new_n1094), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1093), .A2(new_n757), .A3(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(G317), .A2(new_n783), .B1(new_n789), .B2(G311), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT52), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n268), .B1(new_n814), .B2(G322), .ZN(new_n1099));
  INV_X1    g0899(.A(G294), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1099), .B1(new_n1100), .B2(new_n786), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n409), .A2(new_n802), .B1(new_n792), .B2(new_n1074), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n845), .A2(new_n810), .B1(new_n551), .B2(new_n779), .ZN(new_n1103));
  OR4_X1    g0903(.A1(new_n1098), .A2(new_n1101), .A3(new_n1102), .A4(new_n1103), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n779), .A2(new_n271), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n845), .A2(new_n446), .B1(new_n802), .B2(new_n224), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n1105), .B(new_n1106), .C1(G68), .C2(new_n793), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n847), .A2(new_n252), .B1(new_n796), .B2(new_n788), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(new_n1108), .B(KEYINPUT51), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n816), .A2(new_n393), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n322), .B1(new_n814), .B2(G143), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n1107), .A2(new_n1109), .A3(new_n1110), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n822), .B1(new_n1104), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1064), .B1(new_n549), .B2(new_n211), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n246), .B2(new_n766), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n758), .B1(new_n1115), .B2(KEYINPUT117), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1113), .B(new_n1116), .C1(KEYINPUT117), .C2(new_n1115), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n1117), .B1(new_n971), .B2(new_n825), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1021), .B1(new_n1093), .B2(new_n1095), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1023), .A2(new_n753), .ZN(new_n1120));
  OAI211_X1 g0920(.A(new_n1096), .B(new_n1118), .C1(new_n1119), .C2(new_n1120), .ZN(G390));
  NAND2_X1  g0921(.A1(new_n892), .A2(new_n900), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n771), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n845), .A2(new_n409), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n1105), .B(new_n1124), .C1(G283), .C2(new_n783), .ZN(new_n1125));
  OAI22_X1  g0925(.A1(new_n786), .A2(new_n549), .B1(new_n795), .B2(new_n1100), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n268), .B(new_n1126), .C1(G116), .C2(new_n789), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1125), .A2(new_n794), .A3(new_n851), .A4(new_n1127), .ZN(new_n1128));
  XNOR2_X1  g0928(.A(KEYINPUT54), .B(G143), .ZN(new_n1129));
  OAI22_X1  g0929(.A1(new_n788), .A2(new_n852), .B1(new_n786), .B2(new_n1129), .ZN(new_n1130));
  AOI211_X1 g0930(.A(new_n322), .B(new_n1130), .C1(G125), .C2(new_n814), .ZN(new_n1131));
  NOR2_X1   g0931(.A1(new_n792), .A2(new_n252), .ZN(new_n1132));
  XNOR2_X1  g0932(.A(new_n1132), .B(KEYINPUT53), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n801), .A2(G137), .B1(new_n803), .B2(G50), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G159), .A2(new_n780), .B1(new_n783), .B2(G128), .ZN(new_n1135));
  NAND4_X1  g0935(.A1(new_n1131), .A2(new_n1133), .A3(new_n1134), .A4(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n822), .B1(new_n1128), .B2(new_n1136), .ZN(new_n1137));
  AOI211_X1 g0937(.A(new_n843), .B(new_n1137), .C1(new_n256), .C2(new_n864), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1123), .A2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n893), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n909), .B1(new_n738), .B2(new_n832), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1140), .B1(new_n1141), .B2(new_n908), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n908), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n832), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n691), .B(new_n1144), .C1(new_n745), .C2(new_n748), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1143), .B1(new_n1145), .B2(new_n909), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n893), .B1(new_n883), .B2(new_n889), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1122), .A2(new_n1142), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n939), .A2(new_n715), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1149), .A2(G330), .A3(new_n922), .ZN(new_n1150));
  OAI21_X1  g0950(.A(KEYINPUT118), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g0951(.A(new_n832), .B(new_n1143), .C1(new_n735), .C2(new_n736), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1148), .A2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT118), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1150), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n911), .A2(new_n893), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(new_n892), .B2(new_n900), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n890), .A2(new_n1140), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n749), .A2(new_n832), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(new_n910), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1158), .B1(new_n1160), .B2(new_n1143), .ZN(new_n1161));
  OAI211_X1 g0961(.A(new_n1154), .B(new_n1155), .C1(new_n1157), .C2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1151), .A2(new_n1153), .A3(new_n1162), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1139), .B1(new_n1163), .B2(new_n756), .ZN(new_n1164));
  AND3_X1   g0964(.A1(new_n899), .A2(KEYINPUT39), .A3(new_n883), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT39), .B1(new_n883), .B2(new_n889), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1142), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n909), .B1(new_n749), .B2(new_n832), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1147), .B1(new_n1168), .B2(new_n908), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1150), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1170), .A2(new_n1154), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n950), .A2(new_n918), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1172), .A2(new_n470), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n666), .B(new_n1173), .C1(new_n750), .C2(new_n471), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n839), .B(G330), .C1(new_n931), .C2(new_n932), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n908), .ZN(new_n1177));
  AND2_X1   g0977(.A1(new_n1177), .A2(new_n1168), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1152), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n832), .B1(new_n735), .B2(new_n736), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1155), .B1(new_n1180), .B2(new_n908), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1179), .B1(new_n1181), .B2(new_n1141), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1171), .A2(new_n1151), .A3(new_n1175), .A4(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1175), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n709), .B1(new_n1163), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1164), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G378));
  NAND2_X1  g0987(.A1(new_n665), .A2(new_n294), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n267), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n1189), .A2(new_n689), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1190), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n313), .B1(new_n1189), .B2(new_n689), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n771), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n446), .B1(G33), .B2(G41), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1201), .B1(new_n322), .B2(new_n708), .ZN(new_n1202));
  OAI22_X1  g1002(.A1(new_n847), .A2(new_n551), .B1(new_n802), .B2(new_n331), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1203), .B1(G97), .B2(new_n801), .ZN(new_n1204));
  OAI22_X1  g1004(.A1(new_n788), .A2(new_n409), .B1(new_n786), .B2(new_n395), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n708), .B(new_n322), .C1(new_n795), .C2(new_n1074), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND4_X1  g1007(.A1(new_n1204), .A2(new_n1035), .A3(new_n1069), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT58), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1202), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  AOI211_X1 g1010(.A(G33), .B(G41), .C1(new_n814), .C2(G124), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1129), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n789), .B1(new_n793), .B2(new_n1212), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT119), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n783), .A2(G125), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n846), .B2(new_n786), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n845), .A2(new_n852), .B1(new_n252), .B2(new_n779), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1214), .A2(new_n1216), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(KEYINPUT59), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1211), .B1(new_n796), .B2(new_n802), .C1(new_n1218), .C2(new_n1219), .ZN(new_n1220));
  AND2_X1   g1020(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n1210), .B1(new_n1209), .B2(new_n1208), .C1(new_n1220), .C2(new_n1221), .ZN(new_n1222));
  AND2_X1   g1022(.A1(new_n1222), .A2(new_n774), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n843), .B(new_n1223), .C1(new_n446), .C2(new_n864), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1200), .A2(new_n1224), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n914), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n901), .A2(new_n902), .A3(new_n912), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n935), .A2(new_n946), .ZN(new_n1230));
  AND2_X1   g1030(.A1(new_n883), .A2(new_n889), .ZN(new_n1231));
  OAI21_X1  g1031(.A(G330), .B1(new_n1231), .B2(new_n947), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1199), .B1(new_n1230), .B2(new_n1233), .ZN(new_n1234));
  AOI211_X1 g1034(.A(new_n1232), .B(new_n1198), .C1(new_n935), .C2(new_n946), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1229), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  AOI211_X1 g1036(.A(KEYINPUT109), .B(KEYINPUT40), .C1(new_n904), .C2(new_n940), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n944), .B1(new_n943), .B2(new_n945), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1233), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1198), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1230), .A2(new_n1233), .A3(new_n1199), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1240), .A2(new_n915), .A3(new_n1241), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1236), .A2(new_n1242), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1226), .B1(new_n1243), .B2(new_n757), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1182), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1175), .B1(new_n1163), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1246), .A2(KEYINPUT57), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT120), .ZN(new_n1248));
  AND3_X1   g1048(.A1(new_n1240), .A2(new_n915), .A3(new_n1241), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(new_n1240), .A2(new_n1241), .B1(new_n1228), .B2(new_n1227), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1248), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  OAI21_X1  g1051(.A(KEYINPUT120), .B1(new_n1242), .B2(new_n1229), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1247), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AOI22_X1  g1053(.A1(new_n1183), .A2(new_n1175), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n753), .B1(new_n1254), .B2(KEYINPUT57), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1244), .B1(new_n1253), .B2(new_n1255), .ZN(G375));
  OAI211_X1 g1056(.A(new_n1174), .B(new_n1179), .C1(new_n1181), .C2(new_n1141), .ZN(new_n1257));
  XOR2_X1   g1057(.A(new_n1000), .B(KEYINPUT121), .Z(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1184), .A2(new_n1257), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n908), .A2(new_n771), .ZN(new_n1261));
  OAI22_X1  g1061(.A1(new_n845), .A2(new_n551), .B1(new_n847), .B2(new_n1100), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(G97), .B2(new_n793), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n780), .A2(new_n396), .ZN(new_n1264));
  OAI22_X1  g1064(.A1(new_n788), .A2(new_n1074), .B1(new_n786), .B2(new_n409), .ZN(new_n1265));
  AOI211_X1 g1065(.A(new_n268), .B(new_n1265), .C1(G303), .C2(new_n814), .ZN(new_n1266));
  NAND4_X1  g1066(.A1(new_n1263), .A2(new_n1029), .A3(new_n1264), .A4(new_n1266), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n779), .A2(new_n446), .B1(new_n792), .B2(new_n796), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1268), .B1(G132), .B2(new_n783), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n322), .B1(new_n814), .B2(G128), .ZN(new_n1270));
  AOI22_X1  g1070(.A1(new_n789), .A2(G137), .B1(new_n816), .B2(G150), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(new_n801), .A2(new_n1212), .B1(new_n803), .B2(G58), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1269), .A2(new_n1270), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n822), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  AOI211_X1 g1074(.A(new_n843), .B(new_n1274), .C1(new_n222), .C2(new_n864), .ZN(new_n1275));
  AOI22_X1  g1075(.A1(new_n1182), .A2(new_n757), .B1(new_n1261), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1260), .A2(new_n1276), .ZN(G381));
  OR3_X1    g1077(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1278));
  NOR4_X1   g1078(.A1(G387), .A2(new_n1278), .A3(G390), .A4(G381), .ZN(new_n1279));
  XNOR2_X1  g1079(.A(new_n1279), .B(KEYINPUT122), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1244), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1243), .A2(new_n1246), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT57), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n709), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT120), .B1(new_n1236), .B2(new_n1242), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1248), .B1(new_n1286), .B2(new_n915), .ZN(new_n1287));
  OAI211_X1 g1087(.A(KEYINPUT57), .B(new_n1246), .C1(new_n1285), .C2(new_n1287), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1281), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1289), .A2(new_n1186), .ZN(new_n1290));
  OR2_X1    g1090(.A1(new_n1280), .A2(new_n1290), .ZN(G407));
  NAND2_X1  g1091(.A1(new_n690), .A2(G213), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1289), .A2(new_n1186), .A3(new_n1293), .ZN(new_n1294));
  OAI211_X1 g1094(.A(G213), .B(new_n1294), .C1(new_n1280), .C2(new_n1290), .ZN(G409));
  NAND2_X1  g1095(.A1(G375), .A2(G378), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n756), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1297));
  OAI21_X1  g1097(.A(KEYINPUT123), .B1(new_n1297), .B2(new_n1226), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n757), .B1(new_n1285), .B2(new_n1287), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1225), .ZN(new_n1301));
  NAND3_X1  g1101(.A1(new_n1243), .A2(new_n1246), .A3(new_n1259), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1186), .A2(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1298), .A2(new_n1301), .A3(new_n1303), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n709), .B1(new_n1182), .B2(new_n1175), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT60), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1257), .A2(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1141), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n734), .A2(G330), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT98), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1309), .A2(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n734), .A2(KEYINPUT98), .A3(G330), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1311), .A2(new_n1312), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1143), .B1(new_n1313), .B2(new_n832), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1308), .B1(new_n1314), .B2(new_n1155), .ZN(new_n1315));
  NAND4_X1  g1115(.A1(new_n1315), .A2(KEYINPUT60), .A3(new_n1174), .A4(new_n1179), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1305), .A2(new_n1307), .A3(new_n1316), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1317), .A2(new_n1276), .ZN(new_n1318));
  INV_X1    g1118(.A(G384), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1320), .A2(KEYINPUT125), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT125), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1318), .A2(new_n1322), .A3(new_n1319), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1317), .A2(G384), .A3(new_n1276), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1324), .A2(KEYINPUT124), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT124), .ZN(new_n1326));
  NAND4_X1  g1126(.A1(new_n1317), .A2(new_n1326), .A3(G384), .A4(new_n1276), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1321), .A2(new_n1323), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  NAND4_X1  g1128(.A1(new_n1296), .A2(new_n1304), .A3(new_n1292), .A4(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1329), .A2(KEYINPUT62), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1331));
  OR2_X1    g1131(.A1(new_n1292), .A2(KEYINPUT126), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1322), .B1(new_n1318), .B2(new_n1319), .ZN(new_n1333));
  AOI211_X1 g1133(.A(KEYINPUT125), .B(G384), .C1(new_n1317), .C2(new_n1276), .ZN(new_n1334));
  OAI211_X1 g1134(.A(new_n1331), .B(new_n1332), .C1(new_n1333), .C2(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1293), .A2(G2897), .ZN(new_n1336));
  INV_X1    g1136(.A(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1328), .A2(new_n1336), .A3(new_n1332), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1304), .ZN(new_n1340));
  OAI21_X1  g1140(.A(new_n1292), .B1(new_n1289), .B2(new_n1186), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1338), .B(new_n1339), .C1(new_n1340), .C2(new_n1341), .ZN(new_n1342));
  INV_X1    g1142(.A(KEYINPUT61), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1293), .B1(G375), .B2(G378), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT62), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1344), .A2(new_n1345), .A3(new_n1328), .A4(new_n1304), .ZN(new_n1346));
  NAND4_X1  g1146(.A1(new_n1330), .A2(new_n1342), .A3(new_n1343), .A4(new_n1346), .ZN(new_n1347));
  XNOR2_X1  g1147(.A(G393), .B(new_n827), .ZN(new_n1348));
  INV_X1    g1148(.A(new_n1348), .ZN(new_n1349));
  AND3_X1   g1149(.A1(G390), .A2(new_n1025), .A3(new_n1049), .ZN(new_n1350));
  AOI21_X1  g1150(.A(G390), .B1(new_n1025), .B2(new_n1049), .ZN(new_n1351));
  OAI21_X1  g1151(.A(new_n1349), .B1(new_n1350), .B2(new_n1351), .ZN(new_n1352));
  OR2_X1    g1152(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1353));
  AND2_X1   g1153(.A1(new_n1096), .A2(new_n1118), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(G387), .A2(new_n1353), .A3(new_n1354), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(G390), .A2(new_n1025), .A3(new_n1049), .ZN(new_n1356));
  NAND3_X1  g1156(.A1(new_n1355), .A2(new_n1348), .A3(new_n1356), .ZN(new_n1357));
  NAND2_X1  g1157(.A1(new_n1352), .A2(new_n1357), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1347), .A2(new_n1358), .ZN(new_n1359));
  INV_X1    g1159(.A(KEYINPUT63), .ZN(new_n1360));
  AOI21_X1  g1160(.A(new_n1358), .B1(new_n1360), .B2(new_n1329), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1344), .A2(KEYINPUT63), .A3(new_n1328), .A4(new_n1304), .ZN(new_n1362));
  NAND4_X1  g1162(.A1(new_n1361), .A2(new_n1343), .A3(new_n1342), .A4(new_n1362), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1359), .A2(new_n1363), .ZN(G405));
  NAND2_X1  g1164(.A1(new_n1328), .A2(KEYINPUT127), .ZN(new_n1365));
  OAI21_X1  g1165(.A(new_n1331), .B1(new_n1333), .B2(new_n1334), .ZN(new_n1366));
  INV_X1    g1166(.A(KEYINPUT127), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1366), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1365), .A2(new_n1368), .ZN(new_n1369));
  NAND3_X1  g1169(.A1(new_n1369), .A2(new_n1290), .A3(new_n1296), .ZN(new_n1370));
  INV_X1    g1170(.A(new_n1358), .ZN(new_n1371));
  NAND2_X1  g1171(.A1(new_n1296), .A2(new_n1290), .ZN(new_n1372));
  NAND3_X1  g1172(.A1(new_n1372), .A2(new_n1368), .A3(new_n1365), .ZN(new_n1373));
  AND3_X1   g1173(.A1(new_n1370), .A2(new_n1371), .A3(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1371), .B1(new_n1370), .B2(new_n1373), .ZN(new_n1375));
  NOR2_X1   g1175(.A1(new_n1374), .A2(new_n1375), .ZN(G402));
endmodule


