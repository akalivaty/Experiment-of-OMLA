//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 0 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 0 0 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:19 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n448, new_n450, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n540, new_n541, new_n542, new_n544, new_n545, new_n546, new_n547,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n559, new_n561, new_n562, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n577, new_n578, new_n579, new_n580, new_n581,
    new_n583, new_n584, new_n585, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n618, new_n621, new_n623, new_n624, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n858, new_n859, new_n860, new_n861, new_n862, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT67), .Z(G217));
  NOR4_X1   g026(.A1(G219), .A2(G220), .A3(G221), .A4(G218), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT68), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(KEYINPUT3), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  INV_X1    g043(.A(G2105), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n469), .A2(G101), .A3(G2104), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  NAND3_X1  g046(.A1(new_n471), .A2(G137), .A3(new_n469), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n468), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(G160));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n469), .ZN(new_n475));
  INV_X1    g050(.A(G136), .ZN(new_n476));
  OR3_X1    g051(.A1(new_n475), .A2(KEYINPUT69), .A3(new_n476), .ZN(new_n477));
  OAI21_X1  g052(.A(KEYINPUT69), .B1(new_n475), .B2(new_n476), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n469), .ZN(new_n483));
  NAND4_X1  g058(.A1(new_n477), .A2(new_n478), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  INV_X1    g060(.A(G138), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(KEYINPUT70), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n487), .A2(new_n462), .A3(new_n464), .A4(new_n469), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n471), .A2(KEYINPUT4), .A3(new_n469), .A4(new_n487), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n462), .A2(new_n464), .A3(G126), .A4(G2105), .ZN(new_n492));
  OR2_X1    g067(.A1(G102), .A2(G2105), .ZN(new_n493));
  OAI211_X1 g068(.A(new_n493), .B(G2104), .C1(G114), .C2(new_n469), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n490), .A2(new_n491), .A3(new_n492), .A4(new_n494), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  AND2_X1   g071(.A1(new_n494), .A2(new_n492), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT71), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n497), .A2(new_n498), .A3(new_n490), .A4(new_n491), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n496), .A2(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g080(.A(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  OAI21_X1  g082(.A(KEYINPUT72), .B1(new_n507), .B2(G651), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT72), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n509), .A2(new_n510), .A3(KEYINPUT6), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n508), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT73), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n513), .B1(new_n510), .B2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n507), .A2(KEYINPUT73), .A3(G651), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n506), .A2(new_n512), .A3(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G88), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n512), .A2(new_n516), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n520), .A2(new_n501), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(G50), .ZN(new_n522));
  NAND2_X1  g097(.A1(G75), .A2(G543), .ZN(new_n523));
  INV_X1    g098(.A(G62), .ZN(new_n524));
  OAI21_X1  g099(.A(new_n523), .B1(new_n505), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n525), .A2(G651), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n519), .A2(new_n522), .A3(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(G166));
  INV_X1    g103(.A(KEYINPUT75), .ZN(new_n529));
  NAND4_X1  g104(.A1(new_n506), .A2(new_n512), .A3(new_n516), .A4(G89), .ZN(new_n530));
  NAND4_X1  g105(.A1(new_n512), .A2(new_n516), .A3(G51), .A4(G543), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n506), .A2(G63), .A3(G651), .ZN(new_n532));
  AND3_X1   g107(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  XNOR2_X1  g109(.A(new_n534), .B(KEYINPUT74), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT7), .ZN(new_n536));
  AOI21_X1  g111(.A(new_n529), .B1(new_n533), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT7), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n535), .B(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n530), .A2(new_n531), .A3(new_n532), .ZN(new_n540));
  NOR3_X1   g115(.A1(new_n539), .A2(new_n540), .A3(KEYINPUT75), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n537), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(G168));
  AOI22_X1  g118(.A1(new_n506), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n544));
  OR2_X1    g119(.A1(new_n544), .A2(new_n510), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n518), .A2(G90), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n521), .A2(G52), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(new_n518), .A2(G81), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n521), .A2(G43), .ZN(new_n551));
  NAND2_X1  g126(.A1(G68), .A2(G543), .ZN(new_n552));
  INV_X1    g127(.A(G56), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n505), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n550), .A2(new_n551), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G860), .ZN(G153));
  AND3_X1   g133(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G36), .ZN(G176));
  NAND2_X1  g135(.A1(G1), .A2(G3), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n561), .B(KEYINPUT8), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n559), .A2(new_n562), .ZN(G188));
  NAND4_X1  g138(.A1(new_n512), .A2(new_n516), .A3(G53), .A4(G543), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT9), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(G78), .A2(G543), .ZN(new_n569));
  INV_X1    g144(.A(G65), .ZN(new_n570));
  OAI21_X1  g145(.A(new_n569), .B1(new_n505), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n571), .A2(G651), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n517), .B2(new_n573), .ZN(new_n574));
  NOR2_X1   g149(.A1(new_n568), .A2(new_n574), .ZN(new_n575));
  INV_X1    g150(.A(new_n575), .ZN(G299));
  INV_X1    g151(.A(KEYINPUT76), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n577), .B1(new_n537), .B2(new_n541), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n533), .A2(new_n529), .A3(new_n536), .ZN(new_n579));
  OAI21_X1  g154(.A(KEYINPUT75), .B1(new_n539), .B2(new_n540), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT76), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n578), .A2(new_n581), .ZN(G286));
  NAND2_X1  g157(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT77), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n519), .A2(new_n522), .A3(new_n584), .A4(new_n526), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G303));
  OAI21_X1  g161(.A(G651), .B1(new_n506), .B2(G74), .ZN(new_n587));
  XNOR2_X1  g162(.A(new_n587), .B(KEYINPUT78), .ZN(new_n588));
  AOI22_X1  g163(.A1(G87), .A2(new_n518), .B1(new_n521), .B2(G49), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(G288));
  NAND2_X1  g165(.A1(G73), .A2(G543), .ZN(new_n591));
  INV_X1    g166(.A(G61), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n591), .B1(new_n505), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(G651), .ZN(new_n594));
  NAND4_X1  g169(.A1(new_n512), .A2(new_n516), .A3(G48), .A4(G543), .ZN(new_n595));
  NAND4_X1  g170(.A1(new_n506), .A2(new_n512), .A3(new_n516), .A4(G86), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  AOI22_X1  g172(.A1(new_n506), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n598));
  OR2_X1    g173(.A1(new_n598), .A2(new_n510), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n521), .A2(G47), .ZN(new_n600));
  XNOR2_X1  g175(.A(KEYINPUT79), .B(G85), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n518), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g177(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(G290));
  NAND2_X1  g178(.A1(G301), .A2(G868), .ZN(new_n604));
  INV_X1    g179(.A(G92), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n517), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g181(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(G79), .A2(G543), .ZN(new_n609));
  INV_X1    g184(.A(G66), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n505), .B2(new_n610), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n521), .A2(G54), .B1(G651), .B2(new_n611), .ZN(new_n612));
  AND2_X1   g187(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n604), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n604), .B1(new_n613), .B2(G868), .ZN(G321));
  INV_X1    g190(.A(G868), .ZN(new_n616));
  NAND2_X1  g191(.A1(G299), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g192(.A1(new_n578), .A2(new_n581), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G297));
  OAI21_X1  g194(.A(new_n617), .B1(new_n618), .B2(new_n616), .ZN(G280));
  INV_X1    g195(.A(G559), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n613), .B1(new_n621), .B2(G860), .ZN(G148));
  NAND2_X1  g197(.A1(new_n613), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n623), .A2(G868), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n624), .B1(G868), .B2(new_n557), .ZN(G323));
  XNOR2_X1  g200(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g201(.A(new_n475), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G135), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT84), .ZN(new_n629));
  OR2_X1    g204(.A1(G99), .A2(G2105), .ZN(new_n630));
  OAI211_X1 g205(.A(new_n630), .B(G2104), .C1(G111), .C2(new_n469), .ZN(new_n631));
  INV_X1    g206(.A(G123), .ZN(new_n632));
  OAI21_X1  g207(.A(new_n631), .B1(new_n479), .B2(new_n632), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n629), .A2(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT85), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(G2096), .ZN(new_n636));
  NAND2_X1  g211(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT82), .B(KEYINPUT13), .Z(new_n638));
  NOR2_X1   g213(.A1(KEYINPUT83), .A2(G2100), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n641));
  NOR3_X1   g216(.A1(new_n463), .A2(new_n461), .A3(G2105), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n640), .B(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n636), .A2(new_n637), .A3(new_n644), .ZN(G156));
  XNOR2_X1  g220(.A(G2427), .B(G2438), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(G2430), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT15), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(G2435), .Z(new_n649));
  NAND2_X1  g224(.A1(new_n649), .A2(KEYINPUT14), .ZN(new_n650));
  XOR2_X1   g225(.A(G2443), .B(G2446), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XOR2_X1   g227(.A(G1341), .B(G1348), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT16), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G2451), .B(G2454), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n655), .B(new_n656), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  INV_X1    g233(.A(new_n658), .ZN(G401));
  XNOR2_X1  g234(.A(G2072), .B(G2078), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(KEYINPUT17), .ZN(new_n661));
  XOR2_X1   g236(.A(G2067), .B(G2678), .Z(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(G2084), .B(G2090), .Z(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n664), .B(new_n666), .C1(new_n663), .C2(new_n660), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT87), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n663), .A2(new_n665), .A3(new_n660), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(KEYINPUT86), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT18), .ZN(new_n671));
  OR3_X1    g246(.A1(new_n661), .A2(new_n666), .A3(new_n663), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n668), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(G2096), .B(G2100), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(G227));
  XOR2_X1   g251(.A(KEYINPUT89), .B(KEYINPUT20), .Z(new_n677));
  XNOR2_X1  g252(.A(G1956), .B(G2474), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT88), .ZN(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND2_X1  g255(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1971), .B(G1976), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT19), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n677), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n681), .A2(new_n683), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n681), .A2(new_n677), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n687), .A2(new_n685), .ZN(new_n688));
  OAI221_X1 g263(.A(new_n684), .B1(new_n685), .B2(new_n686), .C1(new_n688), .C2(new_n683), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1981), .ZN(new_n690));
  XOR2_X1   g265(.A(G1991), .B(G1996), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n693));
  INV_X1    g268(.A(G1986), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XOR2_X1   g270(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n692), .B(new_n697), .ZN(G229));
  NAND2_X1  g273(.A1(G171), .A2(G16), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G5), .B2(G16), .ZN(new_n700));
  INV_X1    g275(.A(G1961), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(KEYINPUT24), .A2(G34), .ZN(new_n703));
  INV_X1    g278(.A(G29), .ZN(new_n704));
  NAND2_X1  g279(.A1(KEYINPUT24), .A2(G34), .ZN(new_n705));
  AND3_X1   g280(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n473), .B2(G29), .ZN(new_n707));
  INV_X1    g282(.A(G2084), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n627), .A2(G141), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n480), .A2(G129), .ZN(new_n711));
  NAND3_X1  g286(.A1(new_n469), .A2(G105), .A3(G2104), .ZN(new_n712));
  NAND3_X1  g287(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT26), .Z(new_n714));
  NAND4_X1  g289(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G29), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G29), .B2(G32), .ZN(new_n718));
  XOR2_X1   g293(.A(KEYINPUT27), .B(G1996), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  OAI211_X1 g295(.A(new_n702), .B(new_n709), .C1(new_n718), .C2(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT103), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G16), .ZN(new_n724));
  AND2_X1   g299(.A1(new_n724), .A2(G19), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n725), .B1(new_n556), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(G1341), .ZN(new_n727));
  OR2_X1    g302(.A1(G4), .A2(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n608), .A2(new_n612), .ZN(new_n729));
  OAI211_X1 g304(.A(G1348), .B(new_n728), .C1(new_n729), .C2(new_n724), .ZN(new_n730));
  INV_X1    g305(.A(KEYINPUT28), .ZN(new_n731));
  INV_X1    g306(.A(G26), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n731), .B1(new_n732), .B2(G29), .ZN(new_n733));
  NOR2_X1   g308(.A1(new_n732), .A2(G29), .ZN(new_n734));
  AOI22_X1  g309(.A1(G128), .A2(new_n480), .B1(new_n627), .B2(G140), .ZN(new_n735));
  OAI21_X1  g310(.A(G2104), .B1(new_n469), .B2(G116), .ZN(new_n736));
  NOR2_X1   g311(.A1(G104), .A2(G2105), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT96), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n735), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  AOI21_X1  g314(.A(new_n734), .B1(new_n739), .B2(G29), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n733), .B1(new_n740), .B2(new_n731), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G2067), .ZN(new_n742));
  AND3_X1   g317(.A1(new_n727), .A2(new_n730), .A3(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n741), .A2(G2067), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n728), .B1(new_n729), .B2(new_n724), .ZN(new_n745));
  INV_X1    g320(.A(G1348), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n743), .A2(KEYINPUT97), .A3(new_n744), .A4(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT97), .ZN(new_n749));
  NAND4_X1  g324(.A1(new_n747), .A2(new_n727), .A3(new_n730), .A4(new_n742), .ZN(new_n750));
  INV_X1    g325(.A(new_n744), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n749), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n704), .A2(G27), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G164), .B2(new_n704), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n755), .A2(G2078), .ZN(new_n756));
  OR2_X1    g331(.A1(G29), .A2(G33), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n627), .A2(G139), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n469), .A2(G103), .A3(G2104), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT25), .Z(new_n760));
  AOI22_X1  g335(.A1(new_n471), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(KEYINPUT98), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n758), .B(new_n760), .C1(new_n762), .C2(new_n469), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT99), .Z(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(new_n704), .ZN(new_n765));
  INV_X1    g340(.A(G2072), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n723), .A2(new_n753), .A3(new_n756), .A4(new_n767), .ZN(new_n768));
  OR2_X1    g343(.A1(new_n700), .A2(new_n701), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n718), .A2(new_n720), .ZN(new_n770));
  INV_X1    g345(.A(KEYINPUT30), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n771), .A2(G28), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT102), .Z(new_n773));
  OAI211_X1 g348(.A(new_n773), .B(new_n704), .C1(new_n771), .C2(G28), .ZN(new_n774));
  AND3_X1   g349(.A1(new_n769), .A2(new_n770), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n704), .A2(G35), .ZN(new_n776));
  OAI21_X1  g351(.A(new_n776), .B1(G162), .B2(new_n704), .ZN(new_n777));
  XNOR2_X1  g352(.A(new_n777), .B(KEYINPUT29), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n778), .A2(G2090), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n775), .B(new_n779), .C1(new_n708), .C2(new_n707), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n724), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n724), .ZN(new_n782));
  NOR2_X1   g357(.A1(new_n782), .A2(G1966), .ZN(new_n783));
  NOR3_X1   g358(.A1(new_n768), .A2(new_n780), .A3(new_n783), .ZN(new_n784));
  XNOR2_X1  g359(.A(KEYINPUT31), .B(G11), .ZN(new_n785));
  OAI22_X1  g360(.A1(new_n778), .A2(G2090), .B1(new_n755), .B2(G2078), .ZN(new_n786));
  INV_X1    g361(.A(new_n786), .ZN(new_n787));
  NAND3_X1  g362(.A1(new_n724), .A2(KEYINPUT23), .A3(G20), .ZN(new_n788));
  INV_X1    g363(.A(KEYINPUT23), .ZN(new_n789));
  INV_X1    g364(.A(G20), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n789), .B1(new_n790), .B2(G16), .ZN(new_n791));
  OAI211_X1 g366(.A(new_n788), .B(new_n791), .C1(new_n575), .C2(new_n724), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(G1956), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  NAND4_X1  g369(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n794), .ZN(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n724), .A2(G24), .ZN(new_n797));
  INV_X1    g372(.A(G290), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(new_n724), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(new_n694), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OR2_X1    g376(.A1(G25), .A2(G29), .ZN(new_n802));
  AOI22_X1  g377(.A1(G119), .A2(new_n480), .B1(new_n627), .B2(G131), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(new_n469), .B2(G107), .ZN(new_n804));
  NOR2_X1   g379(.A1(G95), .A2(G2105), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT92), .Z(new_n806));
  OAI21_X1  g381(.A(new_n803), .B1(new_n804), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n802), .B1(new_n807), .B2(new_n704), .ZN(new_n808));
  XNOR2_X1  g383(.A(KEYINPUT35), .B(G1991), .ZN(new_n809));
  XOR2_X1   g384(.A(new_n809), .B(KEYINPUT93), .Z(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n811), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n808), .A2(new_n811), .ZN(new_n814));
  NOR3_X1   g389(.A1(new_n801), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  INV_X1    g390(.A(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(G288), .A2(G16), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n724), .A2(G23), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT33), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT33), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n817), .A2(new_n821), .A3(new_n818), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(G1976), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g400(.A(G22), .ZN(new_n826));
  OAI21_X1  g401(.A(KEYINPUT94), .B1(new_n826), .B2(G16), .ZN(new_n827));
  OR3_X1    g402(.A1(new_n826), .A2(KEYINPUT94), .A3(G16), .ZN(new_n828));
  OAI211_X1 g403(.A(new_n827), .B(new_n828), .C1(G166), .C2(new_n724), .ZN(new_n829));
  XOR2_X1   g404(.A(KEYINPUT95), .B(G1971), .Z(new_n830));
  XNOR2_X1  g405(.A(new_n829), .B(new_n830), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n820), .A2(G1976), .A3(new_n822), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n825), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  OR2_X1    g408(.A1(G305), .A2(new_n724), .ZN(new_n834));
  OR2_X1    g409(.A1(G6), .A2(G16), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT32), .ZN(new_n837));
  INV_X1    g412(.A(G1981), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n837), .B(new_n838), .ZN(new_n839));
  INV_X1    g414(.A(KEYINPUT34), .ZN(new_n840));
  OR3_X1    g415(.A1(new_n833), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n840), .B1(new_n833), .B2(new_n839), .ZN(new_n842));
  AOI21_X1  g417(.A(new_n816), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT36), .ZN(new_n844));
  NOR2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  AOI211_X1 g420(.A(KEYINPUT36), .B(new_n816), .C1(new_n841), .C2(new_n842), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  NOR3_X1   g423(.A1(new_n629), .A2(new_n633), .A3(new_n704), .ZN(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n765), .A2(new_n766), .ZN(new_n851));
  XOR2_X1   g426(.A(new_n851), .B(KEYINPUT100), .Z(new_n852));
  INV_X1    g427(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n796), .A2(new_n848), .A3(new_n850), .A4(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n782), .A2(G1966), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n855), .B(KEYINPUT101), .Z(new_n856));
  NOR2_X1   g431(.A1(new_n854), .A2(new_n856), .ZN(G311));
  INV_X1    g432(.A(KEYINPUT104), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n858), .B1(new_n854), .B2(new_n856), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n795), .A2(new_n847), .A3(new_n852), .ZN(new_n860));
  INV_X1    g435(.A(new_n856), .ZN(new_n861));
  NAND4_X1  g436(.A1(new_n860), .A2(KEYINPUT104), .A3(new_n861), .A4(new_n850), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n859), .A2(new_n862), .ZN(G150));
  NAND2_X1  g438(.A1(new_n518), .A2(G93), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n521), .A2(G55), .ZN(new_n865));
  NAND2_X1  g440(.A1(G80), .A2(G543), .ZN(new_n866));
  INV_X1    g441(.A(G67), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n866), .B1(new_n505), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(G651), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n864), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(G860), .ZN(new_n871));
  XOR2_X1   g446(.A(new_n871), .B(KEYINPUT37), .Z(new_n872));
  NAND2_X1  g447(.A1(new_n613), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n873), .B(KEYINPUT38), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT39), .ZN(new_n875));
  OR3_X1    g450(.A1(new_n556), .A2(new_n870), .A3(KEYINPUT105), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n870), .A2(KEYINPUT105), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT105), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n864), .A2(new_n865), .A3(new_n878), .A4(new_n869), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n877), .A2(new_n556), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n875), .B(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n872), .B1(new_n883), .B2(G860), .ZN(G145));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n495), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g461(.A1(new_n497), .A2(KEYINPUT106), .A3(new_n490), .A4(new_n491), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n484), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n634), .B(G160), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n764), .B(new_n715), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n627), .A2(G142), .ZN(new_n893));
  OAI21_X1  g468(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n469), .A2(G118), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n893), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n896), .B1(G130), .B2(new_n480), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n897), .B(new_n807), .Z(new_n898));
  OR2_X1    g473(.A1(new_n892), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n739), .B(new_n643), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n892), .A2(new_n898), .ZN(new_n901));
  NAND3_X1  g476(.A1(new_n899), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n900), .B1(new_n899), .B2(new_n901), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n891), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  INV_X1    g481(.A(new_n891), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n890), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  INV_X1    g485(.A(G37), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n905), .A2(new_n908), .A3(new_n890), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  XNOR2_X1  g488(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n913), .B(new_n914), .ZN(G395));
  NAND2_X1  g490(.A1(new_n870), .A2(new_n616), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n613), .A2(G299), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n729), .A2(new_n575), .ZN(new_n918));
  AND2_X1   g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n919), .A2(KEYINPUT41), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n917), .A2(KEYINPUT41), .A3(new_n918), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n922), .ZN(new_n923));
  XOR2_X1   g498(.A(new_n881), .B(new_n623), .Z(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n925), .B1(new_n919), .B2(new_n924), .ZN(new_n926));
  XNOR2_X1  g501(.A(G288), .B(new_n527), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n927), .B(G305), .ZN(new_n928));
  XNOR2_X1  g503(.A(new_n928), .B(G290), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT108), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n929), .B1(new_n930), .B2(KEYINPUT42), .ZN(new_n931));
  XNOR2_X1  g506(.A(new_n926), .B(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(KEYINPUT42), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n932), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n916), .B1(new_n934), .B2(new_n616), .ZN(G295));
  OAI21_X1  g510(.A(new_n916), .B1(new_n934), .B2(new_n616), .ZN(G331));
  INV_X1    g511(.A(KEYINPUT43), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT109), .ZN(new_n938));
  AOI21_X1  g513(.A(G301), .B1(new_n578), .B2(new_n581), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n542), .A2(G171), .ZN(new_n940));
  OAI211_X1 g515(.A(new_n882), .B(new_n938), .C1(new_n939), .C2(new_n940), .ZN(new_n941));
  OAI21_X1  g516(.A(new_n882), .B1(new_n939), .B2(new_n940), .ZN(new_n942));
  INV_X1    g517(.A(new_n940), .ZN(new_n943));
  OAI211_X1 g518(.A(new_n943), .B(new_n881), .C1(new_n618), .C2(G301), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n942), .A2(new_n944), .A3(KEYINPUT109), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n923), .A2(new_n941), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n917), .A2(new_n918), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n942), .A2(new_n944), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n946), .A2(new_n929), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n911), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT111), .ZN(new_n951));
  INV_X1    g526(.A(new_n929), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n945), .A2(new_n941), .ZN(new_n954));
  AOI21_X1  g529(.A(new_n953), .B1(new_n954), .B2(new_n947), .ZN(new_n955));
  AOI211_X1 g530(.A(KEYINPUT110), .B(new_n919), .C1(new_n945), .C2(new_n941), .ZN(new_n956));
  OR2_X1    g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n922), .B1(new_n942), .B2(new_n944), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n951), .B(new_n952), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n955), .A2(new_n956), .A3(new_n958), .ZN(new_n960));
  OAI21_X1  g535(.A(KEYINPUT111), .B1(new_n960), .B2(new_n929), .ZN(new_n961));
  AOI211_X1 g536(.A(new_n937), .B(new_n950), .C1(new_n959), .C2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n950), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n946), .A2(new_n948), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n952), .ZN(new_n965));
  AOI21_X1  g540(.A(KEYINPUT43), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  OAI21_X1  g541(.A(KEYINPUT44), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT44), .ZN(new_n968));
  AOI211_X1 g543(.A(KEYINPUT43), .B(new_n950), .C1(new_n959), .C2(new_n961), .ZN(new_n969));
  AOI21_X1  g544(.A(new_n937), .B1(new_n963), .B2(new_n965), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n968), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n971), .ZN(G397));
  INV_X1    g547(.A(G1384), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n496), .A2(new_n973), .A3(new_n499), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n888), .A2(KEYINPUT45), .A3(new_n973), .ZN(new_n977));
  NAND4_X1  g552(.A1(new_n468), .A2(G40), .A3(new_n470), .A4(new_n472), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(KEYINPUT56), .B(G2072), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n976), .A2(new_n977), .A3(new_n979), .A4(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT57), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(new_n568), .B2(new_n574), .ZN(new_n983));
  INV_X1    g558(.A(new_n574), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n984), .A2(KEYINPUT57), .A3(new_n567), .A4(new_n566), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n983), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n495), .A2(new_n973), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n978), .B1(new_n987), .B2(KEYINPUT50), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT50), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n496), .A2(new_n989), .A3(new_n973), .A4(new_n499), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G1956), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(new_n981), .A2(new_n986), .A3(new_n993), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n981), .A2(new_n993), .ZN(new_n995));
  INV_X1    g570(.A(new_n986), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT120), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g572(.A(KEYINPUT120), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n998), .B(new_n986), .C1(new_n981), .C2(new_n993), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n994), .B(KEYINPUT61), .C1(new_n997), .C2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n987), .A2(new_n978), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  XOR2_X1   g577(.A(KEYINPUT58), .B(G1341), .Z(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n976), .A2(new_n977), .A3(new_n979), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1004), .B1(new_n1005), .B2(G1996), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n557), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1007), .A2(KEYINPUT59), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT59), .ZN(new_n1009));
  NAND3_X1  g584(.A1(new_n1006), .A2(new_n1009), .A3(new_n557), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT61), .ZN(new_n1012));
  INV_X1    g587(.A(new_n994), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n986), .B1(new_n981), .B2(new_n993), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n1000), .A2(new_n1011), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n978), .B1(new_n974), .B2(KEYINPUT50), .ZN(new_n1017));
  AND3_X1   g592(.A1(new_n495), .A2(new_n989), .A3(new_n973), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g594(.A(G1348), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2067), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1001), .A2(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  OAI21_X1  g598(.A(KEYINPUT119), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT119), .ZN(new_n1025));
  AOI211_X1 g600(.A(new_n978), .B(new_n1018), .C1(new_n974), .C2(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1025), .B(new_n1022), .C1(new_n1026), .C2(G1348), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n729), .B1(new_n1028), .B2(KEYINPUT60), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT60), .ZN(new_n1030));
  AOI211_X1 g605(.A(new_n1030), .B(new_n613), .C1(new_n1024), .C2(new_n1027), .ZN(new_n1031));
  OAI22_X1  g606(.A1(new_n1029), .A2(new_n1031), .B1(KEYINPUT60), .B2(new_n1028), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1016), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1028), .A2(new_n729), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n997), .A2(new_n999), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n994), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT53), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n1005), .B2(G2078), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n701), .ZN(new_n1040));
  AOI21_X1  g615(.A(G1384), .B1(new_n886), .B2(new_n887), .ZN(new_n1041));
  OR2_X1    g616(.A1(new_n1041), .A2(KEYINPUT45), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n978), .B1(new_n1041), .B2(KEYINPUT45), .ZN(new_n1043));
  OR2_X1    g618(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1044));
  NAND2_X1  g619(.A1(KEYINPUT123), .A2(G2078), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1037), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1042), .A2(new_n1043), .A3(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1038), .A2(new_n1040), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT124), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1038), .A2(KEYINPUT124), .A3(new_n1040), .A4(new_n1047), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1050), .A2(G171), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n987), .A2(new_n975), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(KEYINPUT116), .A3(new_n979), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n973), .A4(new_n499), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT116), .ZN(new_n1056));
  AOI21_X1  g631(.A(KEYINPUT45), .B1(new_n495), .B2(new_n973), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(new_n978), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1054), .A2(new_n1055), .A3(new_n1058), .ZN(new_n1059));
  OR2_X1    g634(.A1(new_n1037), .A2(G2078), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1038), .B(new_n1040), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(G301), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1052), .A2(new_n1062), .A3(KEYINPUT54), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(G171), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT54), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1064), .B(new_n1065), .C1(G171), .C2(new_n1048), .ZN(new_n1066));
  AOI22_X1  g641(.A1(new_n1033), .A2(new_n1036), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(G8), .ZN(new_n1068));
  INV_X1    g643(.A(G1966), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1059), .A2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1017), .A2(new_n708), .A3(new_n1019), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1068), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(G168), .A2(new_n1068), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1072), .A2(KEYINPUT51), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT121), .ZN(new_n1076));
  AOI22_X1  g651(.A1(new_n1026), .A2(new_n708), .B1(new_n1059), .B2(new_n1069), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1076), .B1(new_n1077), .B2(new_n1068), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1073), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(KEYINPUT121), .A3(G8), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1078), .A2(new_n1079), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT122), .ZN(new_n1083));
  AND3_X1   g658(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT51), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1083), .B1(new_n1082), .B2(KEYINPUT51), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1075), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1079), .A2(new_n1077), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1086), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT55), .ZN(new_n1091));
  AOI211_X1 g666(.A(new_n1091), .B(new_n1068), .C1(new_n583), .C2(new_n585), .ZN(new_n1092));
  OR2_X1    g667(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(G1971), .B1(new_n1043), .B2(new_n976), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n1039), .A2(G2090), .ZN(new_n1095));
  OAI211_X1 g670(.A(new_n1093), .B(G8), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(G305), .A2(G1981), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n594), .A2(new_n596), .A3(new_n838), .A4(new_n595), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(KEYINPUT112), .B(KEYINPUT49), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1101), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT113), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n1105));
  AOI211_X1 g680(.A(new_n1105), .B(new_n1101), .C1(new_n1098), .C2(new_n1099), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(G8), .B1(new_n987), .B2(new_n978), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1108), .B1(new_n1109), .B2(KEYINPUT49), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1104), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT114), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1114));
  NAND3_X1  g689(.A1(new_n1114), .A2(KEYINPUT114), .A3(new_n1110), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n991), .A2(G2090), .ZN(new_n1117));
  OAI21_X1  g692(.A(G8), .B1(new_n1094), .B2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1090), .A2(new_n1092), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G288), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1108), .B1(new_n1121), .B2(G1976), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT52), .ZN(new_n1123));
  OR2_X1    g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1122), .B(new_n1123), .C1(G1976), .C2(new_n1121), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1116), .A2(new_n1120), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1126));
  NOR2_X1   g701(.A1(new_n1097), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1067), .A2(new_n1089), .A3(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT117), .ZN(new_n1130));
  NOR4_X1   g705(.A1(new_n1077), .A2(new_n1130), .A3(new_n1068), .A4(G286), .ZN(new_n1131));
  AOI21_X1  g706(.A(KEYINPUT117), .B1(new_n1072), .B2(new_n618), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n1096), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1129), .B1(new_n1133), .B2(new_n1126), .ZN(new_n1134));
  AND4_X1   g709(.A1(new_n1116), .A2(new_n1120), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1072), .A2(new_n618), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n1130), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1072), .A2(KEYINPUT117), .A3(new_n618), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1135), .A2(new_n1139), .A3(KEYINPUT118), .A4(new_n1096), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT63), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1134), .A2(new_n1140), .A3(new_n1141), .ZN(new_n1142));
  AOI211_X1 g717(.A(G1976), .B(G288), .C1(new_n1113), .C2(new_n1115), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1099), .ZN(new_n1144));
  OAI211_X1 g719(.A(G8), .B(new_n1002), .C1(new_n1143), .C2(new_n1144), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n1114), .A2(KEYINPUT114), .A3(new_n1110), .ZN(new_n1146));
  AOI21_X1  g721(.A(KEYINPUT114), .B1(new_n1114), .B2(new_n1110), .ZN(new_n1147));
  OAI211_X1 g722(.A(new_n1124), .B(new_n1125), .C1(new_n1146), .C2(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT115), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1148), .A2(new_n1149), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1116), .A2(KEYINPUT115), .A3(new_n1124), .A4(new_n1125), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(G8), .B1(new_n1095), .B2(new_n1094), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1153), .A2(new_n1119), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1096), .B(new_n1154), .C1(new_n1131), .C2(new_n1132), .ZN(new_n1155));
  OAI21_X1  g730(.A(KEYINPUT63), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1142), .A2(new_n1145), .A3(new_n1156), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1150), .A2(new_n1097), .A3(new_n1151), .ZN(new_n1158));
  AND3_X1   g733(.A1(new_n1128), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1081), .A2(new_n1079), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1072), .A2(KEYINPUT121), .ZN(new_n1161));
  OAI21_X1  g736(.A(KEYINPUT51), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1162), .A2(KEYINPUT122), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1082), .A2(new_n1083), .A3(KEYINPUT51), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1074), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  OAI21_X1  g740(.A(KEYINPUT62), .B1(new_n1165), .B2(new_n1087), .ZN(new_n1166));
  INV_X1    g741(.A(new_n1064), .ZN(new_n1167));
  INV_X1    g742(.A(KEYINPUT62), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1086), .A2(new_n1168), .A3(new_n1088), .ZN(new_n1169));
  NAND4_X1  g744(.A1(new_n1166), .A2(new_n1167), .A3(new_n1127), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT125), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n1064), .B1(new_n1089), .B2(KEYINPUT62), .ZN(new_n1173));
  NAND4_X1  g748(.A1(new_n1173), .A2(KEYINPUT125), .A3(new_n1127), .A4(new_n1169), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1159), .A2(new_n1172), .A3(new_n1174), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1042), .A2(new_n978), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n739), .B(new_n1021), .ZN(new_n1177));
  INV_X1    g752(.A(G1996), .ZN(new_n1178));
  XNOR2_X1  g753(.A(new_n715), .B(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1177), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g755(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n807), .A2(new_n810), .ZN(new_n1182));
  OR2_X1    g757(.A1(new_n807), .A2(new_n810), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1181), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g759(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1185), .B1(new_n694), .B2(new_n798), .ZN(new_n1186));
  NOR2_X1   g761(.A1(G290), .A2(G1986), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1176), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1175), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1177), .A2(new_n716), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT127), .ZN(new_n1191));
  AOI22_X1  g766(.A1(new_n1190), .A2(new_n1176), .B1(new_n1191), .B2(KEYINPUT46), .ZN(new_n1192));
  NOR2_X1   g767(.A1(new_n1191), .A2(KEYINPUT46), .ZN(new_n1193));
  AND3_X1   g768(.A1(new_n1176), .A2(new_n1178), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g769(.A(new_n1193), .B1(new_n1176), .B2(new_n1178), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1192), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  XOR2_X1   g771(.A(new_n1196), .B(KEYINPUT47), .Z(new_n1197));
  OAI22_X1  g772(.A1(new_n1180), .A2(new_n1183), .B1(G2067), .B2(new_n739), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1198), .A2(new_n1176), .ZN(new_n1199));
  XNOR2_X1  g774(.A(new_n1199), .B(KEYINPUT126), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1176), .A2(new_n1187), .ZN(new_n1201));
  XOR2_X1   g776(.A(new_n1201), .B(KEYINPUT48), .Z(new_n1202));
  AOI21_X1  g777(.A(new_n1202), .B1(new_n1176), .B2(new_n1184), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1197), .A2(new_n1200), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1189), .A2(new_n1204), .ZN(G329));
  assign    G231 = 1'b0;
  AOI21_X1  g780(.A(new_n950), .B1(new_n959), .B2(new_n961), .ZN(new_n1207));
  AOI21_X1  g781(.A(new_n970), .B1(new_n1207), .B2(new_n937), .ZN(new_n1208));
  AND3_X1   g782(.A1(new_n905), .A2(new_n908), .A3(new_n890), .ZN(new_n1209));
  NOR3_X1   g783(.A1(new_n1209), .A2(new_n909), .A3(G37), .ZN(new_n1210));
  INV_X1    g784(.A(G319), .ZN(new_n1211));
  NOR2_X1   g785(.A1(G229), .A2(new_n1211), .ZN(new_n1212));
  INV_X1    g786(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n658), .A2(new_n675), .ZN(new_n1214));
  NOR4_X1   g788(.A1(new_n1208), .A2(new_n1210), .A3(new_n1213), .A4(new_n1214), .ZN(G308));
  NAND2_X1  g789(.A1(new_n1207), .A2(new_n937), .ZN(new_n1216));
  INV_X1    g790(.A(new_n970), .ZN(new_n1217));
  NAND2_X1  g791(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g792(.A(new_n1214), .ZN(new_n1219));
  NAND4_X1  g793(.A1(new_n1218), .A2(new_n913), .A3(new_n1212), .A4(new_n1219), .ZN(G225));
endmodule


