//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:27 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n723, new_n724, new_n725, new_n726, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n754, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT69), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  INV_X1    g005(.A(G134), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(KEYINPUT66), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT66), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G134), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n191), .B1(new_n196), .B2(new_n190), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT11), .B1(new_n196), .B2(new_n190), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n197), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT11), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT66), .B(G134), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n200), .B1(new_n201), .B2(G137), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n201), .A2(G137), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n202), .A2(new_n203), .A3(new_n204), .A4(new_n191), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n199), .A2(new_n205), .ZN(new_n206));
  OR2_X1    g020(.A1(KEYINPUT64), .A2(G146), .ZN(new_n207));
  NAND2_X1  g021(.A1(KEYINPUT64), .A2(G146), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n207), .A2(KEYINPUT65), .A3(G143), .A4(new_n208), .ZN(new_n209));
  AND2_X1   g023(.A1(KEYINPUT0), .A2(G128), .ZN(new_n210));
  AND2_X1   g024(.A1(KEYINPUT64), .A2(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(KEYINPUT64), .A2(G146), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NOR3_X1   g027(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT65), .B1(new_n215), .B2(G143), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n209), .B(new_n210), .C1(new_n214), .C2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(KEYINPUT0), .A2(G128), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n210), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(G143), .B1(new_n207), .B2(new_n208), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n218), .A2(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n206), .A2(new_n226), .ZN(new_n227));
  XOR2_X1   g041(.A(G116), .B(G119), .Z(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT2), .B(G113), .ZN(new_n229));
  XNOR2_X1  g043(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g044(.A(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G128), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n207), .A2(G143), .A3(new_n208), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n232), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n207), .A2(new_n208), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n223), .B1(new_n235), .B2(new_n213), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT68), .B1(new_n234), .B2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT68), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n211), .A2(new_n212), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n222), .B1(new_n239), .B2(G143), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n241), .B1(new_n239), .B2(G143), .ZN(new_n242));
  OAI211_X1 g056(.A(new_n238), .B(new_n240), .C1(new_n242), .C2(new_n232), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n233), .A2(new_n216), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n244), .A2(new_n209), .A3(new_n245), .ZN(new_n246));
  AND3_X1   g060(.A1(new_n237), .A2(new_n243), .A3(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(G137), .B1(new_n193), .B2(new_n195), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT67), .ZN(new_n249));
  OAI22_X1  g063(.A1(new_n248), .A2(new_n249), .B1(G134), .B2(new_n190), .ZN(new_n250));
  NOR3_X1   g064(.A1(new_n201), .A2(KEYINPUT67), .A3(G137), .ZN(new_n251));
  OAI21_X1  g065(.A(G131), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n205), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n227), .B(new_n231), .C1(new_n247), .C2(new_n253), .ZN(new_n254));
  NOR2_X1   g068(.A1(G237), .A2(G953), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(G210), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT27), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT26), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT27), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n256), .B(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT26), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND3_X1   g076(.A1(new_n258), .A2(new_n262), .A3(G101), .ZN(new_n263));
  AOI21_X1  g077(.A(G101), .B1(new_n258), .B2(new_n262), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n254), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n237), .A2(new_n243), .A3(new_n246), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(new_n205), .A3(new_n252), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n268), .A2(new_n227), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n270), .B1(new_n206), .B2(new_n226), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n231), .B1(new_n268), .B2(new_n272), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n266), .B1(new_n271), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT31), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n189), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AND2_X1   g090(.A1(new_n252), .A2(new_n205), .ZN(new_n277));
  AOI22_X1  g091(.A1(new_n277), .A2(new_n267), .B1(new_n206), .B2(new_n226), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n273), .B1(KEYINPUT30), .B2(new_n278), .ZN(new_n279));
  AND2_X1   g093(.A1(new_n254), .A2(new_n265), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT69), .A3(KEYINPUT31), .ZN(new_n282));
  INV_X1    g096(.A(new_n254), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n231), .B1(new_n268), .B2(new_n227), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT28), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n254), .A2(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n265), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT71), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n276), .A2(new_n282), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n265), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n269), .A2(new_n230), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n286), .B1(new_n292), .B2(new_n254), .ZN(new_n293));
  INV_X1    g107(.A(new_n287), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XOR2_X1   g109(.A(KEYINPUT70), .B(KEYINPUT31), .Z(new_n296));
  AOI22_X1  g110(.A1(new_n295), .A2(KEYINPUT71), .B1(new_n274), .B2(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n188), .B1(new_n290), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT73), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n287), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n254), .A2(KEYINPUT73), .A3(new_n286), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT29), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n291), .A2(new_n302), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n285), .A2(new_n300), .A3(new_n301), .A4(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G902), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT74), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n279), .A2(new_n254), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n291), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n285), .A2(new_n287), .A3(new_n265), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n310), .A2(new_n302), .A3(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n304), .A2(KEYINPUT74), .A3(new_n305), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n308), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  AOI22_X1  g128(.A1(new_n298), .A2(KEYINPUT32), .B1(new_n314), .B2(G472), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n298), .B2(KEYINPUT32), .ZN(new_n316));
  AOI21_X1  g130(.A(KEYINPUT69), .B1(new_n281), .B2(KEYINPUT31), .ZN(new_n317));
  AOI211_X1 g131(.A(new_n189), .B(new_n275), .C1(new_n279), .C2(new_n280), .ZN(new_n318));
  OAI22_X1  g132(.A1(new_n317), .A2(new_n318), .B1(new_n295), .B2(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n274), .A2(new_n296), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n320), .B1(new_n288), .B2(new_n289), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n187), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT32), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n315), .A2(new_n316), .A3(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G214), .B1(G237), .B2(G902), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT83), .ZN(new_n328));
  INV_X1    g142(.A(G125), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n237), .A2(new_n243), .A3(new_n329), .A4(new_n246), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n225), .A2(G125), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n328), .B1(new_n330), .B2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n328), .ZN(new_n333));
  INV_X1    g147(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n332), .A2(new_n334), .A3(KEYINPUT86), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT86), .B1(new_n332), .B2(new_n334), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G224), .ZN(new_n339));
  XOR2_X1   g153(.A(new_n339), .B(KEYINPUT85), .Z(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(KEYINPUT84), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n336), .A2(new_n337), .A3(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n341), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n330), .A2(new_n331), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(KEYINPUT83), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n344), .B1(new_n346), .B2(new_n333), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n343), .B1(new_n347), .B2(new_n335), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT3), .ZN(new_n351));
  INV_X1    g165(.A(G107), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n352), .A3(G104), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n349), .A2(G107), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n350), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(G101), .ZN(new_n356));
  INV_X1    g170(.A(G101), .ZN(new_n357));
  NAND4_X1  g171(.A1(new_n350), .A2(new_n353), .A3(new_n357), .A4(new_n354), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(KEYINPUT4), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n355), .A2(new_n360), .A3(G101), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n230), .A2(new_n359), .A3(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n354), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n349), .A2(G107), .ZN(new_n364));
  OAI21_X1  g178(.A(G101), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n365), .A2(new_n358), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n228), .A2(new_n229), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT5), .ZN(new_n368));
  INV_X1    g182(.A(G119), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G116), .ZN(new_n370));
  OAI211_X1 g184(.A(G113), .B(new_n370), .C1(new_n228), .C2(new_n368), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n366), .A2(new_n367), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n362), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(KEYINPUT81), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT6), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n362), .A2(new_n376), .A3(new_n372), .ZN(new_n377));
  XNOR2_X1  g191(.A(G110), .B(G122), .ZN(new_n378));
  INV_X1    g192(.A(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n374), .A2(new_n375), .A3(new_n377), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(KEYINPUT82), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n378), .B1(new_n373), .B2(KEYINPUT81), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n383));
  NAND4_X1  g197(.A1(new_n382), .A2(new_n383), .A3(new_n375), .A4(new_n377), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n377), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n362), .A2(new_n372), .A3(new_n378), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n386), .A2(KEYINPUT6), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n342), .A2(new_n348), .A3(new_n385), .A4(new_n388), .ZN(new_n389));
  OAI21_X1  g203(.A(G210), .B1(G237), .B2(G902), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n371), .A2(new_n367), .ZN(new_n391));
  XNOR2_X1  g205(.A(new_n391), .B(new_n366), .ZN(new_n392));
  XOR2_X1   g206(.A(new_n378), .B(KEYINPUT8), .Z(new_n393));
  OAI21_X1  g207(.A(new_n387), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n340), .A2(KEYINPUT7), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n345), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n333), .A4(new_n340), .ZN(new_n397));
  AOI21_X1  g211(.A(G902), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n389), .A2(new_n390), .A3(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n399), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n390), .B1(new_n389), .B2(new_n398), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n327), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G475), .ZN(new_n403));
  OR2_X1    g217(.A1(new_n329), .A2(G140), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT16), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n329), .A2(G140), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(KEYINPUT79), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT79), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(new_n329), .A3(G140), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(KEYINPUT77), .A2(G140), .ZN(new_n412));
  NOR2_X1   g226(.A1(KEYINPUT77), .A2(G140), .ZN(new_n413));
  OAI21_X1  g227(.A(G125), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT78), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT78), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n416), .B(G125), .C1(new_n412), .C2(new_n413), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n411), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n406), .B1(new_n418), .B2(new_n405), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n419), .A2(G146), .ZN(new_n420));
  OAI211_X1 g234(.A(new_n215), .B(new_n406), .C1(new_n418), .C2(new_n405), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n255), .A2(G214), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT87), .A3(G143), .ZN(new_n423));
  OR2_X1    g237(.A1(KEYINPUT87), .A2(G143), .ZN(new_n424));
  NAND2_X1  g238(.A1(KEYINPUT87), .A2(G143), .ZN(new_n425));
  NAND4_X1  g239(.A1(new_n424), .A2(G214), .A3(new_n255), .A4(new_n425), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n423), .A2(G131), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(KEYINPUT17), .ZN(new_n428));
  AOI21_X1  g242(.A(G131), .B1(new_n423), .B2(new_n426), .ZN(new_n429));
  OR3_X1    g243(.A1(new_n427), .A2(new_n429), .A3(KEYINPUT17), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n420), .A2(new_n421), .A3(new_n428), .A4(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n239), .A2(new_n404), .A3(new_n407), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n432), .B1(new_n418), .B2(new_n215), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n423), .A2(new_n426), .ZN(new_n434));
  NAND2_X1  g248(.A1(KEYINPUT88), .A2(KEYINPUT18), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n427), .A2(new_n429), .ZN(new_n437));
  OAI211_X1 g251(.A(new_n433), .B(new_n436), .C1(new_n435), .C2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g253(.A(G113), .B(G122), .ZN(new_n440));
  XNOR2_X1  g254(.A(new_n440), .B(new_n349), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT89), .ZN(new_n443));
  AOI21_X1  g257(.A(G902), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n431), .A2(KEYINPUT89), .A3(new_n442), .A4(new_n438), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n403), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n439), .A2(new_n441), .ZN(new_n447));
  AND2_X1   g261(.A1(new_n433), .A2(new_n436), .ZN(new_n448));
  OR2_X1    g262(.A1(new_n437), .A2(new_n435), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n441), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n437), .B1(new_n419), .B2(G146), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT19), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n404), .A2(new_n407), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n418), .B2(new_n452), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n451), .B1(new_n235), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n450), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n447), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(G475), .A2(G902), .ZN(new_n458));
  INV_X1    g272(.A(new_n458), .ZN(new_n459));
  OAI21_X1  g273(.A(KEYINPUT20), .B1(new_n457), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n439), .A2(new_n441), .B1(new_n450), .B2(new_n455), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT20), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n461), .A2(new_n462), .A3(new_n458), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n446), .B1(new_n460), .B2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(G116), .ZN(new_n465));
  OAI21_X1  g279(.A(KEYINPUT90), .B1(new_n465), .B2(G122), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT90), .ZN(new_n467));
  INV_X1    g281(.A(G122), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n467), .A2(new_n468), .A3(G116), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n465), .A2(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(KEYINPUT14), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n472), .A2(new_n473), .A3(G107), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n470), .B(new_n471), .C1(KEYINPUT14), .C2(new_n352), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n213), .A2(G128), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n232), .A2(G143), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT91), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT91), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n480), .B1(new_n476), .B2(new_n477), .ZN(new_n481));
  NOR3_X1   g295(.A1(new_n479), .A2(new_n201), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n478), .A2(KEYINPUT91), .ZN(new_n483));
  XNOR2_X1  g297(.A(G128), .B(G143), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n480), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n196), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g300(.A(new_n474), .B(new_n475), .C1(new_n482), .C2(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n201), .B1(new_n479), .B2(new_n481), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n484), .A2(KEYINPUT13), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n489), .B(G134), .C1(KEYINPUT13), .C2(new_n476), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n352), .B1(new_n470), .B2(new_n471), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n470), .A2(new_n352), .A3(new_n471), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n488), .B(new_n490), .C1(new_n491), .C2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT9), .B(G234), .ZN(new_n495));
  INV_X1    g309(.A(G217), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(G953), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n487), .A2(new_n493), .A3(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n499), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n487), .A2(new_n493), .A3(KEYINPUT92), .A4(new_n497), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n305), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n505), .A3(G478), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(G478), .ZN(new_n507));
  NAND4_X1  g321(.A1(new_n502), .A2(new_n305), .A3(new_n503), .A4(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(G234), .A2(G237), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(G952), .A3(new_n338), .ZN(new_n512));
  INV_X1    g326(.A(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n511), .A2(G902), .A3(G953), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g329(.A(KEYINPUT21), .B(G898), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n513), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n464), .A2(new_n510), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT93), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND4_X1  g335(.A1(new_n464), .A2(KEYINPUT93), .A3(new_n510), .A4(new_n518), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n402), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(G234), .ZN(new_n524));
  OAI21_X1  g338(.A(G217), .B1(new_n524), .B2(G902), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT75), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n420), .A2(new_n421), .ZN(new_n528));
  OAI21_X1  g342(.A(KEYINPUT23), .B1(new_n232), .B2(G119), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n529), .B(KEYINPUT76), .C1(new_n369), .C2(G128), .ZN(new_n530));
  NOR2_X1   g344(.A1(new_n369), .A2(G128), .ZN(new_n531));
  INV_X1    g345(.A(KEYINPUT76), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n531), .B1(new_n532), .B2(KEYINPUT23), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G110), .ZN(new_n536));
  XOR2_X1   g350(.A(G119), .B(G128), .Z(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT24), .B(G110), .ZN(new_n538));
  OAI22_X1  g352(.A1(new_n535), .A2(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n528), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n432), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n536), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n537), .A2(new_n538), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n420), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n338), .A2(G221), .A3(G234), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n547), .B(KEYINPUT22), .ZN(new_n548));
  XNOR2_X1  g362(.A(new_n548), .B(new_n190), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n541), .A2(new_n546), .A3(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n545), .A2(new_n420), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n539), .B1(new_n420), .B2(new_n421), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n549), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n551), .A2(new_n554), .A3(new_n305), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n527), .B1(new_n555), .B2(KEYINPUT25), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n551), .A2(new_n554), .A3(new_n557), .A4(new_n305), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n551), .A2(new_n554), .ZN(new_n559));
  NOR2_X1   g373(.A1(new_n526), .A2(G902), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n556), .A2(new_n558), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G221), .B1(new_n495), .B2(G902), .ZN(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(G469), .ZN(new_n564));
  NOR2_X1   g378(.A1(new_n564), .A2(new_n305), .ZN(new_n565));
  XNOR2_X1  g379(.A(G110), .B(G140), .ZN(new_n566));
  INV_X1    g380(.A(G227), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(G953), .ZN(new_n568));
  XNOR2_X1  g382(.A(new_n566), .B(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n206), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n267), .A2(KEYINPUT10), .A3(new_n366), .ZN(new_n571));
  INV_X1    g385(.A(new_n246), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n232), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n244), .B2(new_n209), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n366), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT80), .B(KEYINPUT10), .Z(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AND2_X1   g391(.A1(new_n359), .A2(new_n361), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n226), .ZN(new_n579));
  AND4_X1   g393(.A1(new_n570), .A2(new_n571), .A3(new_n577), .A4(new_n579), .ZN(new_n580));
  AOI22_X1  g394(.A1(new_n575), .A2(new_n576), .B1(new_n578), .B2(new_n226), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n570), .B1(new_n581), .B2(new_n571), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n569), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n569), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n571), .A2(new_n577), .A3(new_n570), .A4(new_n579), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n575), .B1(new_n267), .B2(new_n366), .ZN(new_n586));
  AND3_X1   g400(.A1(new_n586), .A2(KEYINPUT12), .A3(new_n206), .ZN(new_n587));
  AOI21_X1  g401(.A(KEYINPUT12), .B1(new_n586), .B2(new_n206), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n584), .B(new_n585), .C1(new_n587), .C2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(G902), .B1(new_n583), .B2(new_n589), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n565), .B1(new_n590), .B2(new_n564), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n581), .A2(new_n571), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n206), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n593), .A2(new_n584), .A3(new_n585), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(KEYINPUT12), .A3(new_n206), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n586), .A2(new_n206), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT12), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n580), .B1(new_n595), .B2(new_n598), .ZN(new_n599));
  OAI211_X1 g413(.A(new_n594), .B(G469), .C1(new_n599), .C2(new_n584), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n563), .B1(new_n591), .B2(new_n600), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n326), .A2(new_n523), .A3(new_n561), .A4(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  INV_X1    g417(.A(new_n327), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT94), .ZN(new_n605));
  AOI21_X1  g419(.A(new_n604), .B1(new_n400), .B2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n389), .A2(new_n398), .ZN(new_n607));
  INV_X1    g421(.A(new_n390), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n609), .A2(KEYINPUT94), .A3(new_n399), .ZN(new_n610));
  INV_X1    g424(.A(G478), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n504), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(KEYINPUT95), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n504), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n502), .A2(new_n616), .A3(new_n503), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n499), .A2(KEYINPUT33), .A3(new_n501), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n611), .A2(G902), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n613), .A2(new_n615), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n621), .A2(new_n464), .ZN(new_n622));
  AND4_X1   g436(.A1(new_n518), .A2(new_n606), .A3(new_n610), .A4(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n290), .A2(new_n297), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n305), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n585), .A2(new_n584), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n627), .B1(new_n595), .B2(new_n598), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n584), .B1(new_n593), .B2(new_n585), .ZN(new_n629));
  OAI211_X1 g443(.A(new_n564), .B(new_n305), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n565), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n630), .A2(new_n600), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n632), .A2(new_n561), .A3(new_n562), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n626), .A2(new_n298), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n623), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT96), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT34), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n637), .B(G104), .ZN(G6));
  NAND2_X1  g452(.A1(new_n606), .A2(new_n610), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n464), .A2(new_n509), .A3(new_n518), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n634), .ZN(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  AOI21_X1  g458(.A(G902), .B1(new_n290), .B2(new_n297), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n322), .B1(new_n645), .B2(new_n624), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n541), .A2(new_n546), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n549), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n556), .A2(new_n558), .B1(new_n649), .B2(new_n560), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n651), .A2(new_n562), .A3(new_n632), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n646), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n523), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT37), .B(G110), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  INV_X1    g470(.A(new_n639), .ZN(new_n657));
  INV_X1    g471(.A(new_n652), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n444), .A2(new_n445), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(G475), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n461), .A2(new_n462), .A3(new_n458), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n462), .B1(new_n461), .B2(new_n458), .ZN(new_n662));
  OAI211_X1 g476(.A(new_n509), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  INV_X1    g477(.A(G900), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n515), .A2(new_n664), .ZN(new_n665));
  AOI21_X1  g479(.A(new_n513), .B1(new_n665), .B2(KEYINPUT97), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(KEYINPUT97), .B2(new_n665), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT98), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n663), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n326), .A2(new_n657), .A3(new_n658), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(G128), .ZN(G30));
  NAND3_X1  g485(.A1(new_n609), .A2(KEYINPUT38), .A3(new_n399), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n650), .A2(new_n327), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n509), .ZN(new_n675));
  OR3_X1    g489(.A1(new_n673), .A2(new_n675), .A3(KEYINPUT99), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n609), .A2(new_n399), .ZN(new_n677));
  INV_X1    g491(.A(KEYINPUT38), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g493(.A(KEYINPUT99), .B1(new_n673), .B2(new_n675), .ZN(new_n680));
  AND4_X1   g494(.A1(new_n672), .A2(new_n676), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n632), .A2(new_n562), .ZN(new_n682));
  XOR2_X1   g496(.A(new_n668), .B(KEYINPUT39), .Z(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT40), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n291), .B1(new_n283), .B2(new_n284), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n281), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n624), .B1(new_n688), .B2(new_n305), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n689), .B1(new_n298), .B2(KEYINPUT32), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n316), .A2(new_n690), .A3(new_n325), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n681), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT100), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n681), .A2(new_n686), .A3(KEYINPUT100), .A4(new_n691), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n213), .ZN(G45));
  NAND3_X1  g511(.A1(new_n617), .A2(new_n618), .A3(new_n620), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n504), .A2(new_n614), .A3(new_n611), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n614), .B1(new_n504), .B2(new_n611), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n698), .B1(new_n699), .B2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n668), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n674), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n601), .A3(new_n651), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n326), .A2(new_n657), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT101), .B(G146), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n706), .B(new_n707), .ZN(G48));
  NOR2_X1   g522(.A1(new_n590), .A2(new_n564), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n710), .A2(new_n562), .A3(new_n630), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT102), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g527(.A(new_n630), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n714), .A2(new_n709), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n715), .A2(KEYINPUT102), .A3(new_n562), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n623), .A2(new_n326), .A3(new_n717), .A4(new_n561), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND4_X1  g534(.A1(new_n641), .A2(new_n326), .A3(new_n717), .A4(new_n561), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G116), .ZN(G18));
  NOR3_X1   g536(.A1(new_n714), .A2(new_n709), .A3(new_n563), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n606), .A2(new_n610), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n650), .B1(new_n521), .B2(new_n522), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n326), .A2(new_n724), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G119), .ZN(G21));
  AND3_X1   g541(.A1(new_n713), .A2(new_n518), .A3(new_n716), .ZN(new_n728));
  INV_X1    g542(.A(new_n675), .ZN(new_n729));
  AND3_X1   g543(.A1(new_n606), .A2(new_n610), .A3(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n285), .A2(new_n301), .A3(new_n300), .ZN(new_n731));
  OAI221_X1 g545(.A(new_n320), .B1(new_n275), .B2(new_n274), .C1(new_n731), .C2(new_n265), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n187), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n733), .B1(new_n645), .B2(new_n624), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n561), .B(KEYINPUT103), .Z(new_n736));
  NAND4_X1  g550(.A1(new_n728), .A2(new_n730), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G122), .ZN(G24));
  NOR2_X1   g552(.A1(new_n734), .A2(new_n650), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n739), .A2(new_n724), .A3(new_n703), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND2_X1  g555(.A1(new_n322), .A2(new_n324), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n315), .A2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n609), .A2(new_n327), .A3(new_n399), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n674), .A2(new_n701), .A3(new_n702), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n744), .A2(new_n682), .A3(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n743), .A2(new_n736), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT42), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n744), .A2(new_n682), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n745), .A2(KEYINPUT42), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n326), .A2(new_n561), .A3(new_n749), .A4(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n203), .ZN(G33));
  NAND4_X1  g567(.A1(new_n326), .A2(new_n561), .A3(new_n669), .A4(new_n749), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G134), .ZN(G36));
  INV_X1    g569(.A(new_n744), .ZN(new_n756));
  OAI21_X1  g570(.A(KEYINPUT43), .B1(new_n621), .B2(new_n674), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT43), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n464), .A2(new_n701), .A3(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n757), .A2(KEYINPUT105), .A3(new_n759), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n646), .A3(new_n651), .A4(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT44), .ZN(new_n765));
  OAI21_X1  g579(.A(new_n756), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(KEYINPUT106), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  OAI211_X1 g582(.A(new_n768), .B(new_n756), .C1(new_n764), .C2(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n767), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT104), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n594), .B1(new_n599), .B2(new_n584), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n564), .B1(new_n772), .B2(new_n773), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n565), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n630), .B1(new_n776), .B2(KEYINPUT46), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n772), .A2(new_n773), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(G469), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n772), .A2(new_n773), .ZN(new_n780));
  OAI211_X1 g594(.A(KEYINPUT46), .B(new_n631), .C1(new_n779), .C2(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n562), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n771), .B1(new_n783), .B2(new_n684), .ZN(new_n784));
  OR2_X1    g598(.A1(new_n776), .A2(KEYINPUT46), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n785), .A2(new_n630), .A3(new_n781), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT104), .A3(new_n562), .A4(new_n683), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n764), .A2(new_n765), .ZN(new_n788));
  AND3_X1   g602(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n770), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G137), .ZN(G39));
  INV_X1    g605(.A(KEYINPUT47), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n786), .A2(new_n792), .A3(new_n562), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n794));
  OR3_X1    g608(.A1(new_n744), .A2(new_n561), .A3(new_n745), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n326), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n794), .A3(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G140), .ZN(G42));
  NOR2_X1   g612(.A1(new_n744), .A2(new_n711), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(new_n561), .A3(new_n513), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n691), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n464), .A3(new_n621), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n757), .A2(new_n513), .A3(new_n759), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(KEYINPUT111), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n739), .A3(new_n799), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n715), .A2(new_n563), .ZN(new_n808));
  AOI21_X1  g622(.A(new_n792), .B1(new_n786), .B2(new_n562), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n783), .A2(KEYINPUT47), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n808), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n735), .A2(new_n736), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n804), .A2(new_n812), .A3(new_n756), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  AOI211_X1 g628(.A(new_n327), .B(new_n711), .C1(new_n679), .C2(new_n672), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n804), .A2(new_n812), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NOR2_X1   g632(.A1(KEYINPUT113), .A2(KEYINPUT50), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n804), .A2(new_n812), .A3(new_n815), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n818), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n807), .A2(new_n814), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(KEYINPUT51), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT114), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n818), .A2(KEYINPUT114), .A3(new_n821), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n806), .A2(KEYINPUT51), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n826), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n811), .A2(new_n830), .A3(new_n813), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n830), .B1(new_n811), .B2(new_n813), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n824), .B1(new_n829), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n804), .A2(new_n812), .A3(new_n724), .ZN(new_n835));
  INV_X1    g649(.A(G952), .ZN(new_n836));
  AOI211_X1 g650(.A(new_n836), .B(G953), .C1(new_n801), .C2(new_n622), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n804), .A2(new_n736), .A3(new_n743), .A4(new_n799), .ZN(new_n838));
  NAND2_X1  g652(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  XOR2_X1   g654(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n834), .A2(new_n835), .A3(new_n837), .A4(new_n842), .ZN(new_n843));
  XNOR2_X1  g657(.A(new_n843), .B(KEYINPUT116), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n663), .B1(new_n621), .B2(new_n464), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(new_n518), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n402), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n523), .A2(new_n653), .B1(new_n634), .B2(new_n848), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n652), .A2(new_n509), .A3(new_n674), .A4(new_n668), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n326), .A2(new_n850), .B1(new_n705), .B2(new_n735), .ZN(new_n851));
  OAI211_X1 g665(.A(new_n602), .B(new_n849), .C1(new_n851), .C2(new_n744), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n748), .A2(new_n751), .A3(new_n754), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT108), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n601), .A2(new_n855), .A3(new_n650), .A4(new_n702), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n650), .A2(new_n702), .ZN(new_n857));
  OAI21_X1  g671(.A(KEYINPUT108), .B1(new_n682), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n691), .A2(new_n730), .A3(new_n859), .ZN(new_n860));
  NAND4_X1  g674(.A1(new_n670), .A2(new_n706), .A3(new_n860), .A4(new_n740), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT52), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n854), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n737), .A2(new_n726), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(KEYINPUT107), .A3(new_n718), .A4(new_n721), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n718), .A2(new_n721), .A3(new_n737), .A4(new_n726), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT107), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n845), .B1(new_n865), .B2(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n861), .B(new_n862), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT109), .ZN(new_n875));
  OR2_X1    g689(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n845), .B1(new_n868), .B2(new_n875), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n874), .A2(new_n854), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n872), .A2(new_n873), .A3(new_n878), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT110), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n872), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n865), .A2(new_n871), .A3(new_n845), .ZN(new_n883));
  OAI21_X1  g697(.A(KEYINPUT54), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n872), .A2(new_n878), .ZN(new_n885));
  OAI21_X1  g699(.A(KEYINPUT110), .B1(new_n885), .B2(KEYINPUT54), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n881), .A2(new_n884), .A3(new_n886), .ZN(new_n887));
  OAI22_X1  g701(.A1(new_n844), .A2(new_n887), .B1(G952), .B2(G953), .ZN(new_n888));
  INV_X1    g702(.A(new_n691), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n621), .A2(new_n674), .A3(new_n563), .A4(new_n604), .ZN(new_n890));
  AND2_X1   g704(.A1(new_n736), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n679), .A2(new_n672), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n715), .B(KEYINPUT49), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n889), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n888), .A2(new_n894), .ZN(G75));
  NAND2_X1  g709(.A1(new_n836), .A2(G953), .ZN(new_n896));
  XOR2_X1   g710(.A(new_n896), .B(KEYINPUT118), .Z(new_n897));
  NAND2_X1  g711(.A1(new_n885), .A2(G902), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  AOI21_X1  g713(.A(KEYINPUT56), .B1(new_n899), .B2(G210), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n342), .A2(new_n348), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n385), .A2(new_n388), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n389), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT55), .Z(new_n905));
  OAI21_X1  g719(.A(new_n897), .B1(new_n900), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT56), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n899), .A2(KEYINPUT117), .A3(G210), .ZN(new_n909));
  INV_X1    g723(.A(KEYINPUT117), .ZN(new_n910));
  INV_X1    g724(.A(G210), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n910), .B1(new_n898), .B2(new_n911), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n908), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n906), .A2(new_n913), .ZN(G51));
  INV_X1    g728(.A(new_n897), .ZN(new_n915));
  NOR3_X1   g729(.A1(new_n898), .A2(new_n780), .A3(new_n779), .ZN(new_n916));
  XNOR2_X1  g730(.A(new_n565), .B(KEYINPUT119), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT57), .Z(new_n918));
  AOI21_X1  g732(.A(new_n873), .B1(new_n872), .B2(new_n878), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n918), .B1(new_n879), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n583), .A2(new_n589), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT120), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n916), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n920), .A2(KEYINPUT120), .A3(new_n921), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(G54));
  NAND3_X1  g740(.A1(new_n899), .A2(KEYINPUT58), .A3(G475), .ZN(new_n927));
  AND2_X1   g741(.A1(new_n927), .A2(new_n457), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n927), .A2(new_n457), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n928), .A2(new_n929), .A3(new_n915), .ZN(G60));
  NAND2_X1  g744(.A1(G478), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT59), .Z(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n619), .B1(new_n887), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n879), .A2(new_n919), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n619), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n897), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n934), .A2(new_n937), .ZN(G63));
  NAND2_X1  g752(.A1(G217), .A2(G902), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT60), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n872), .B2(new_n878), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n941), .A2(new_n649), .ZN(new_n942));
  XOR2_X1   g756(.A(new_n559), .B(KEYINPUT121), .Z(new_n943));
  OAI211_X1 g757(.A(new_n942), .B(new_n897), .C1(new_n941), .C2(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n944), .B(new_n945), .ZN(G66));
  NAND4_X1  g760(.A1(new_n867), .A2(new_n870), .A3(new_n602), .A4(new_n849), .ZN(new_n947));
  NAND2_X1  g761(.A1(G224), .A2(G953), .ZN(new_n948));
  OAI22_X1  g762(.A1(new_n947), .A2(G953), .B1(new_n516), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g763(.A(new_n949), .B(KEYINPUT122), .Z(new_n950));
  OAI21_X1  g764(.A(new_n902), .B1(G898), .B2(new_n338), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(G69));
  NOR2_X1   g766(.A1(new_n338), .A2(G900), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n748), .A2(new_n751), .A3(new_n754), .ZN(new_n954));
  AND3_X1   g768(.A1(new_n670), .A2(new_n706), .A3(new_n740), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n955), .A2(new_n797), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n730), .A2(new_n743), .A3(new_n736), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n784), .A2(new_n787), .A3(new_n957), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n790), .A2(new_n954), .A3(new_n956), .A4(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n953), .B1(new_n959), .B2(new_n338), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT126), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n797), .A2(new_n954), .A3(new_n955), .A4(new_n958), .ZN(new_n963));
  AOI21_X1  g777(.A(G953), .B1(new_n963), .B2(new_n790), .ZN(new_n964));
  OAI21_X1  g778(.A(KEYINPUT126), .B1(new_n964), .B2(new_n953), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n268), .A2(new_n272), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n271), .A2(new_n966), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(new_n454), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n962), .A2(new_n965), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n694), .A2(new_n955), .A3(new_n695), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(KEYINPUT62), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n685), .A2(new_n846), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n326), .A2(new_n973), .A3(new_n561), .A4(new_n756), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n797), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT62), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n694), .A2(new_n955), .A3(new_n976), .A4(new_n695), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n972), .A2(new_n790), .A3(new_n975), .A4(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n338), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n968), .B(KEYINPUT123), .Z(new_n980));
  AOI21_X1  g794(.A(new_n970), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n969), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n567), .B2(new_n664), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT124), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n968), .B1(new_n960), .B2(new_n961), .ZN(new_n986));
  NOR3_X1   g800(.A1(new_n964), .A2(KEYINPUT126), .A3(new_n953), .ZN(new_n987));
  OAI211_X1 g801(.A(new_n981), .B(new_n985), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n983), .A2(new_n984), .A3(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n984), .ZN(new_n990));
  INV_X1    g804(.A(new_n988), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n985), .B1(new_n969), .B2(new_n981), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(new_n993), .ZN(G72));
  NAND2_X1  g808(.A1(G472), .A2(G902), .ZN(new_n995));
  XOR2_X1   g809(.A(new_n995), .B(KEYINPUT63), .Z(new_n996));
  OAI21_X1  g810(.A(new_n996), .B1(new_n978), .B2(new_n947), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n309), .B(KEYINPUT127), .Z(new_n998));
  NOR2_X1   g812(.A1(new_n998), .A2(new_n291), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n915), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n310), .A2(new_n281), .ZN(new_n1001));
  OAI211_X1 g815(.A(new_n996), .B(new_n1001), .C1(new_n882), .C2(new_n883), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n996), .B1(new_n959), .B2(new_n947), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1003), .A2(new_n291), .A3(new_n998), .ZN(new_n1004));
  AND3_X1   g818(.A1(new_n1000), .A2(new_n1002), .A3(new_n1004), .ZN(G57));
endmodule


