//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 1 0 1 1 1 1 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:46 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n600, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n609, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044;
  INV_X1    g000(.A(KEYINPUT65), .ZN(new_n187));
  INV_X1    g001(.A(G119), .ZN(new_n188));
  OAI21_X1  g002(.A(KEYINPUT64), .B1(new_n188), .B2(G116), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  INV_X1    g004(.A(G116), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n189), .A2(new_n192), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n191), .A2(G119), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G113), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(KEYINPUT2), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT2), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G113), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  AND3_X1   g014(.A1(new_n193), .A2(new_n195), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n200), .B1(new_n193), .B2(new_n195), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n187), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n190), .B1(new_n191), .B2(G119), .ZN(new_n204));
  NOR3_X1   g018(.A1(new_n188), .A2(KEYINPUT64), .A3(G116), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n195), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(new_n200), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n194), .B1(new_n189), .B2(new_n192), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(new_n200), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(KEYINPUT65), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n203), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT11), .ZN(new_n213));
  INV_X1    g027(.A(G134), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(G137), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(G137), .ZN(new_n216));
  INV_X1    g030(.A(G137), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n217), .A2(KEYINPUT11), .A3(G134), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G131), .ZN(new_n220));
  INV_X1    g034(.A(G131), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n215), .A2(new_n218), .A3(new_n221), .A4(new_n216), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(G146), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G143), .ZN(new_n225));
  INV_X1    g039(.A(G143), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT0), .ZN(new_n229));
  INV_X1    g043(.A(G128), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NOR2_X1   g045(.A1(KEYINPUT0), .A2(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n228), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  XNOR2_X1  g047(.A(G143), .B(G146), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n234), .B1(new_n229), .B2(new_n230), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n233), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(new_n217), .A2(G134), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n214), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n222), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n230), .A2(KEYINPUT1), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n241), .A2(new_n225), .A3(new_n227), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n226), .A2(KEYINPUT1), .A3(G146), .ZN(new_n243));
  OAI211_X1 g057(.A(new_n242), .B(new_n243), .C1(G128), .C2(new_n234), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n223), .A2(new_n236), .B1(new_n240), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n212), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n222), .A2(new_n239), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n241), .A2(new_n225), .A3(new_n227), .ZN(new_n248));
  AOI21_X1  g062(.A(G128), .B1(new_n225), .B2(new_n227), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n247), .B1(new_n250), .B2(new_n243), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n220), .A2(new_n222), .B1(new_n233), .B2(new_n235), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n211), .B(new_n203), .C1(new_n251), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(KEYINPUT28), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT67), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT28), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n258), .B1(new_n246), .B2(new_n253), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT28), .B1(new_n212), .B2(new_n245), .ZN(new_n260));
  OAI21_X1  g074(.A(KEYINPUT67), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(G237), .A2(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G210), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(G101), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n257), .A2(new_n261), .A3(new_n266), .ZN(new_n267));
  AND2_X1   g081(.A1(new_n203), .A2(new_n211), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n251), .A2(new_n252), .A3(KEYINPUT30), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT30), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n223), .A2(new_n236), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n240), .A2(new_n244), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n268), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n246), .ZN(new_n275));
  INV_X1    g089(.A(new_n266), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(KEYINPUT68), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n267), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT29), .ZN(new_n280));
  NAND4_X1  g094(.A1(new_n257), .A2(new_n261), .A3(KEYINPUT68), .A4(new_n266), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n255), .A2(KEYINPUT69), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n284), .B1(new_n259), .B2(new_n260), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT29), .A4(new_n266), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  AND2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n282), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n289), .A2(G472), .ZN(new_n290));
  NOR2_X1   g104(.A1(G472), .A2(G902), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n266), .B1(new_n257), .B2(new_n261), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT66), .B(KEYINPUT31), .Z(new_n293));
  NAND4_X1  g107(.A1(new_n274), .A2(new_n266), .A3(new_n246), .A4(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT30), .B1(new_n251), .B2(new_n252), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n271), .A2(new_n272), .A3(new_n270), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n212), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n246), .ZN(new_n298));
  NOR3_X1   g112(.A1(new_n297), .A2(new_n298), .A3(new_n276), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT66), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n300), .A2(KEYINPUT31), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n294), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n291), .B1(new_n292), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(KEYINPUT32), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT32), .ZN(new_n305));
  OAI211_X1 g119(.A(new_n305), .B(new_n291), .C1(new_n292), .C2(new_n302), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(G234), .ZN(new_n308));
  OAI21_X1  g122(.A(G217), .B1(new_n308), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT23), .ZN(new_n310));
  OAI21_X1  g124(.A(new_n310), .B1(new_n188), .B2(G128), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n188), .A2(G128), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n230), .A2(KEYINPUT23), .A3(G119), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(G110), .ZN(new_n315));
  XOR2_X1   g129(.A(KEYINPUT24), .B(G110), .Z(new_n316));
  XNOR2_X1  g130(.A(G119), .B(G128), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AND2_X1   g132(.A1(G125), .A2(G140), .ZN(new_n319));
  NOR2_X1   g133(.A1(G125), .A2(G140), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT16), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  INV_X1    g135(.A(G125), .ZN(new_n322));
  OR3_X1    g136(.A1(new_n322), .A2(KEYINPUT16), .A3(G140), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n321), .A2(G146), .A3(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(G146), .B1(new_n321), .B2(new_n323), .ZN(new_n325));
  OAI211_X1 g139(.A(new_n315), .B(new_n318), .C1(new_n324), .C2(new_n325), .ZN(new_n326));
  OAI22_X1  g140(.A1(new_n314), .A2(G110), .B1(new_n316), .B2(new_n317), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n321), .A2(new_n323), .A3(G146), .ZN(new_n328));
  INV_X1    g142(.A(new_n320), .ZN(new_n329));
  NAND2_X1  g143(.A1(G125), .A2(G140), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n224), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n327), .A2(new_n328), .A3(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT22), .B(G137), .ZN(new_n334));
  INV_X1    g148(.A(G953), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n335), .A2(G221), .A3(G234), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n334), .B(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n326), .A2(new_n333), .A3(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n337), .B1(new_n326), .B2(new_n333), .ZN(new_n339));
  NOR3_X1   g153(.A1(new_n338), .A2(new_n339), .A3(G902), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT71), .B1(new_n340), .B2(KEYINPUT25), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT70), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT71), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT25), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n341), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n344), .B1(new_n342), .B2(new_n343), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n340), .A2(new_n347), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n309), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n326), .A2(new_n333), .ZN(new_n350));
  INV_X1    g164(.A(new_n337), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n326), .A2(new_n333), .A3(new_n337), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n309), .A2(new_n287), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT72), .B1(new_n349), .B2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT72), .ZN(new_n358));
  INV_X1    g172(.A(new_n356), .ZN(new_n359));
  INV_X1    g173(.A(new_n348), .ZN(new_n360));
  OAI21_X1  g174(.A(new_n344), .B1(new_n354), .B2(G902), .ZN(new_n361));
  AOI21_X1  g175(.A(KEYINPUT70), .B1(new_n361), .B2(KEYINPUT71), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n362), .B2(new_n345), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n358), .B(new_n359), .C1(new_n363), .C2(new_n309), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n290), .A2(new_n307), .B1(new_n357), .B2(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT81), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n366), .B1(new_n230), .B2(G143), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n226), .A2(KEYINPUT81), .A3(G128), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(KEYINPUT13), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(KEYINPUT82), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n367), .A2(new_n368), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT13), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n230), .A2(G143), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n367), .A2(new_n368), .A3(new_n375), .A4(KEYINPUT13), .ZN(new_n376));
  NAND4_X1  g190(.A1(new_n370), .A2(new_n373), .A3(new_n374), .A4(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G134), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n214), .A3(new_n374), .ZN(new_n379));
  NOR2_X1   g193(.A1(KEYINPUT73), .A2(G107), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(KEYINPUT73), .A2(G107), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(G116), .B(G122), .ZN(new_n384));
  XNOR2_X1  g198(.A(new_n383), .B(new_n384), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n378), .A2(new_n379), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n384), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(KEYINPUT83), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n371), .A2(new_n374), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G134), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n379), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n191), .A2(KEYINPUT14), .A3(G122), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n393), .A2(G107), .A3(new_n394), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n391), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n386), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g211(.A(KEYINPUT9), .B(G234), .ZN(new_n398));
  INV_X1    g212(.A(new_n398), .ZN(new_n399));
  AND3_X1   g213(.A1(new_n399), .A2(G217), .A3(new_n335), .ZN(new_n400));
  INV_X1    g214(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(KEYINPUT85), .B1(new_n397), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT85), .ZN(new_n403));
  AOI211_X1 g217(.A(new_n403), .B(new_n400), .C1(new_n386), .C2(new_n396), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n386), .A2(new_n396), .A3(new_n400), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT84), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n386), .A2(new_n396), .A3(KEYINPUT84), .A4(new_n400), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n287), .B1(new_n405), .B2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(G478), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT86), .ZN(new_n413));
  OR2_X1    g227(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(KEYINPUT15), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n411), .A2(new_n416), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G475), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n331), .B(new_n224), .ZN(new_n421));
  AOI21_X1  g235(.A(G143), .B1(new_n262), .B2(G214), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n262), .A2(G143), .A3(G214), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(new_n221), .ZN(new_n427));
  INV_X1    g241(.A(new_n424), .ZN(new_n428));
  OAI21_X1  g242(.A(G131), .B1(new_n428), .B2(new_n422), .ZN(new_n429));
  OAI221_X1 g243(.A(new_n421), .B1(new_n425), .B2(new_n427), .C1(new_n426), .C2(new_n429), .ZN(new_n430));
  NOR2_X1   g244(.A1(new_n324), .A2(new_n325), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n425), .A2(KEYINPUT17), .A3(G131), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n423), .A2(new_n221), .A3(new_n424), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n431), .B(new_n432), .C1(new_n434), .C2(KEYINPUT17), .ZN(new_n435));
  XNOR2_X1  g249(.A(G113), .B(G122), .ZN(new_n436));
  INV_X1    g250(.A(G104), .ZN(new_n437));
  XNOR2_X1  g251(.A(new_n436), .B(new_n437), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n430), .A2(new_n435), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n438), .B1(new_n430), .B2(new_n435), .ZN(new_n440));
  OR2_X1    g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n420), .B1(new_n441), .B2(new_n287), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT19), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT80), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n443), .A2(KEYINPUT80), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n331), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n329), .A2(KEYINPUT80), .A3(new_n443), .A4(new_n330), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n224), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n328), .A3(new_n434), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n438), .B1(new_n430), .B2(new_n450), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n420), .B(new_n287), .C1(new_n439), .C2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(KEYINPUT20), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n439), .A2(new_n451), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(new_n420), .A4(new_n287), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n442), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(G234), .A2(G237), .ZN(new_n458));
  AND3_X1   g272(.A1(new_n458), .A2(G952), .A3(new_n335), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(G902), .A3(G953), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT87), .ZN(new_n461));
  XNOR2_X1  g275(.A(KEYINPUT21), .B(G898), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n419), .A2(new_n457), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G214), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n236), .A2(G125), .ZN(new_n469));
  INV_X1    g283(.A(new_n243), .ZN(new_n470));
  NOR3_X1   g284(.A1(new_n248), .A2(new_n249), .A3(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n469), .B1(G125), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n335), .A2(G224), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(G110), .B(G122), .Z(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n477), .A2(G104), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n478), .B1(new_n381), .B2(new_n382), .ZN(new_n479));
  AOI21_X1  g293(.A(G107), .B1(new_n437), .B2(KEYINPUT3), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n437), .A2(KEYINPUT3), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(G101), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  AND2_X1   g297(.A1(KEYINPUT73), .A2(G107), .ZN(new_n484));
  OAI21_X1  g298(.A(new_n481), .B1(new_n484), .B2(new_n380), .ZN(new_n485));
  INV_X1    g299(.A(G107), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n486), .B1(new_n477), .B2(G104), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n478), .ZN(new_n488));
  INV_X1    g302(.A(G101), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n485), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n483), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n492));
  OAI211_X1 g306(.A(new_n492), .B(G101), .C1(new_n479), .C2(new_n482), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n203), .A2(new_n491), .A3(new_n211), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n209), .A2(KEYINPUT5), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT5), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n196), .B1(new_n194), .B2(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n201), .B1(new_n495), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n437), .B1(new_n484), .B2(new_n380), .ZN(new_n499));
  NAND2_X1  g313(.A1(G104), .A2(G107), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(G101), .A3(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n490), .A2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n498), .A2(new_n503), .ZN(new_n504));
  AOI21_X1  g318(.A(new_n476), .B1(new_n494), .B2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT6), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(KEYINPUT77), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n494), .A2(new_n476), .A3(new_n504), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT75), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g325(.A1(new_n494), .A2(KEYINPUT75), .A3(new_n504), .A4(new_n476), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n505), .A2(new_n506), .ZN(new_n514));
  AND3_X1   g328(.A1(new_n513), .A2(KEYINPUT76), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT76), .B1(new_n513), .B2(new_n514), .ZN(new_n516));
  OAI211_X1 g330(.A(new_n474), .B(new_n508), .C1(new_n515), .C2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n473), .A2(KEYINPUT7), .ZN(new_n518));
  XOR2_X1   g332(.A(new_n472), .B(new_n518), .Z(new_n519));
  AOI21_X1  g333(.A(new_n519), .B1(new_n511), .B2(new_n512), .ZN(new_n520));
  XNOR2_X1  g334(.A(new_n497), .B(KEYINPUT79), .ZN(new_n521));
  INV_X1    g335(.A(new_n495), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n503), .B(new_n210), .C1(new_n521), .C2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n498), .B2(new_n503), .ZN(new_n524));
  XNOR2_X1  g338(.A(new_n475), .B(KEYINPUT78), .ZN(new_n525));
  XOR2_X1   g339(.A(new_n525), .B(KEYINPUT8), .Z(new_n526));
  NAND2_X1  g340(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g341(.A(G902), .B1(new_n520), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n517), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G210), .B1(G237), .B2(G902), .ZN(new_n530));
  INV_X1    g344(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n529), .A2(new_n531), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n517), .A2(new_n528), .A3(new_n530), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n468), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(G469), .ZN(new_n535));
  XNOR2_X1  g349(.A(G110), .B(G140), .ZN(new_n536));
  AND2_X1   g350(.A1(new_n335), .A2(G227), .ZN(new_n537));
  XOR2_X1   g351(.A(new_n536), .B(new_n537), .Z(new_n538));
  NAND3_X1  g352(.A1(new_n244), .A2(new_n490), .A3(new_n501), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT74), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n540), .A2(KEYINPUT10), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n491), .A2(new_n236), .A3(new_n493), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT10), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(KEYINPUT74), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n541), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n545), .A2(new_n223), .ZN(new_n546));
  AND2_X1   g360(.A1(new_n220), .A2(new_n222), .ZN(new_n547));
  NAND4_X1  g361(.A1(new_n541), .A2(new_n547), .A3(new_n542), .A4(new_n544), .ZN(new_n548));
  AOI21_X1  g362(.A(new_n538), .B1(new_n546), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n538), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n502), .A2(new_n471), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n539), .ZN(new_n552));
  AOI21_X1  g366(.A(KEYINPUT12), .B1(new_n552), .B2(new_n223), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT12), .ZN(new_n554));
  AOI211_X1 g368(.A(new_n554), .B(new_n547), .C1(new_n551), .C2(new_n539), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n550), .A2(new_n556), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n535), .B(new_n287), .C1(new_n549), .C2(new_n557), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n548), .B1(new_n555), .B2(new_n553), .ZN(new_n559));
  INV_X1    g373(.A(new_n538), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n546), .A2(new_n548), .A3(new_n538), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n561), .A2(G469), .A3(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n535), .A2(new_n287), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G221), .B1(new_n398), .B2(G902), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g382(.A1(new_n365), .A2(new_n466), .A3(new_n534), .A4(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(new_n569), .B(G101), .ZN(G3));
  NAND2_X1  g384(.A1(new_n357), .A2(new_n364), .ZN(new_n571));
  OAI21_X1  g385(.A(new_n287), .B1(new_n292), .B2(new_n302), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT88), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n303), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n572), .A2(new_n574), .A3(G472), .ZN(new_n577));
  NAND4_X1  g391(.A1(new_n571), .A2(new_n576), .A3(new_n568), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT89), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT33), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n580), .B1(new_n405), .B2(new_n410), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n412), .A2(G902), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n397), .A2(new_n401), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT33), .A3(new_n406), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n411), .A2(new_n412), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n457), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n534), .A2(new_n464), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(KEYINPUT34), .B(G104), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n589), .B(new_n590), .ZN(G6));
  INV_X1    g405(.A(new_n453), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n452), .A2(KEYINPUT20), .ZN(new_n593));
  OAI21_X1  g407(.A(KEYINPUT90), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT90), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n456), .A2(new_n595), .A3(new_n453), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n442), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n597), .B1(new_n418), .B2(new_n417), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT92), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n463), .B(KEYINPUT91), .ZN(new_n601));
  NAND4_X1  g415(.A1(new_n534), .A2(new_n599), .A3(new_n600), .A4(new_n601), .ZN(new_n602));
  AND3_X1   g416(.A1(new_n517), .A2(new_n528), .A3(new_n530), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n530), .B1(new_n517), .B2(new_n528), .ZN(new_n604));
  OAI211_X1 g418(.A(new_n467), .B(new_n601), .C1(new_n603), .C2(new_n604), .ZN(new_n605));
  OAI21_X1  g419(.A(KEYINPUT92), .B1(new_n605), .B2(new_n598), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n579), .B1(new_n602), .B2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G107), .ZN(new_n608));
  XNOR2_X1  g422(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n608), .B(new_n609), .ZN(G9));
  OAI211_X1 g424(.A(new_n467), .B(new_n568), .C1(new_n603), .C2(new_n604), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n351), .A2(KEYINPUT36), .ZN(new_n613));
  XNOR2_X1  g427(.A(new_n350), .B(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n355), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(new_n616), .B1(new_n363), .B2(new_n309), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n576), .A2(new_n577), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(KEYINPUT94), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT94), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n576), .A2(new_n620), .A3(new_n577), .A4(new_n617), .ZN(new_n621));
  NAND4_X1  g435(.A1(new_n612), .A2(new_n619), .A3(new_n466), .A4(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT37), .B(G110), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G12));
  AOI22_X1  g438(.A1(new_n289), .A2(G472), .B1(new_n304), .B2(new_n306), .ZN(new_n625));
  INV_X1    g439(.A(new_n568), .ZN(new_n626));
  INV_X1    g440(.A(new_n617), .ZN(new_n627));
  NOR3_X1   g441(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(G900), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n459), .B1(new_n461), .B2(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  OAI211_X1 g445(.A(new_n597), .B(new_n631), .C1(new_n418), .C2(new_n417), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n628), .A2(new_n534), .A3(new_n633), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n634), .B(G128), .ZN(G30));
  NOR2_X1   g449(.A1(new_n603), .A2(new_n604), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n532), .A2(new_n533), .ZN(new_n639));
  INV_X1    g453(.A(new_n637), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND2_X1   g455(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n643));
  INV_X1    g457(.A(G472), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n275), .A2(new_n266), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n287), .B1(new_n254), .B2(new_n266), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n644), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n304), .B2(new_n306), .ZN(new_n649));
  INV_X1    g463(.A(new_n457), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(new_n417), .B2(new_n418), .ZN(new_n651));
  NOR3_X1   g465(.A1(new_n649), .A2(new_n651), .A3(new_n617), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n642), .A2(new_n643), .A3(new_n467), .A4(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n638), .A2(new_n641), .A3(new_n467), .ZN(new_n654));
  INV_X1    g468(.A(new_n652), .ZN(new_n655));
  OAI21_X1  g469(.A(KEYINPUT96), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n630), .B(KEYINPUT39), .Z(new_n657));
  NAND2_X1  g471(.A1(new_n568), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT40), .Z(new_n659));
  NAND3_X1  g473(.A1(new_n653), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT97), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n653), .A2(new_n656), .A3(KEYINPUT97), .A4(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(new_n226), .ZN(G45));
  OAI21_X1  g479(.A(new_n467), .B1(new_n603), .B2(new_n604), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n587), .A2(new_n631), .ZN(new_n667));
  OAI21_X1  g481(.A(KEYINPUT98), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  AOI211_X1 g482(.A(new_n630), .B(new_n457), .C1(new_n586), .C2(new_n585), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT98), .ZN(new_n670));
  NAND4_X1  g484(.A1(new_n639), .A2(new_n669), .A3(new_n670), .A4(new_n467), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n668), .A2(new_n628), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G146), .ZN(G48));
  NAND2_X1  g487(.A1(new_n290), .A2(new_n307), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n549), .A2(new_n557), .ZN(new_n675));
  OAI21_X1  g489(.A(G469), .B1(new_n675), .B2(G902), .ZN(new_n676));
  AND3_X1   g490(.A1(new_n676), .A2(new_n567), .A3(new_n558), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n571), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  INV_X1    g493(.A(new_n587), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n666), .A2(new_n463), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n679), .A2(new_n681), .A3(KEYINPUT99), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT99), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n683), .B1(new_n588), .B2(new_n678), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(KEYINPUT41), .B(G113), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G15));
  NAND2_X1  g501(.A1(new_n606), .A2(new_n602), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n679), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  OAI211_X1 g504(.A(new_n467), .B(new_n677), .C1(new_n603), .C2(new_n604), .ZN(new_n691));
  NOR4_X1   g505(.A1(new_n691), .A2(new_n625), .A3(new_n465), .A4(new_n627), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n188), .ZN(G21));
  AND3_X1   g507(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT100), .ZN(new_n694));
  AOI21_X1  g508(.A(KEYINPUT100), .B1(new_n283), .B2(new_n285), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n694), .A2(new_n695), .A3(new_n266), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n291), .B1(new_n696), .B2(new_n302), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n359), .B1(new_n363), .B2(new_n309), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n699), .A3(new_n573), .ZN(new_n700));
  INV_X1    g514(.A(new_n677), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n605), .A2(new_n700), .A3(new_n651), .A4(new_n701), .ZN(new_n702));
  XOR2_X1   g516(.A(new_n702), .B(G122), .Z(G24));
  NAND2_X1  g517(.A1(new_n283), .A2(new_n285), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT100), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n266), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n283), .A2(new_n285), .A3(KEYINPUT100), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n302), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n291), .ZN(new_n709));
  OAI211_X1 g523(.A(new_n573), .B(new_n617), .C1(new_n708), .C2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n710), .A2(KEYINPUT101), .ZN(new_n711));
  INV_X1    g525(.A(KEYINPUT101), .ZN(new_n712));
  NAND4_X1  g526(.A1(new_n697), .A2(new_n712), .A3(new_n573), .A4(new_n617), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n691), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n714), .A2(new_n715), .A3(new_n669), .ZN(new_n716));
  XNOR2_X1  g530(.A(KEYINPUT102), .B(G125), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(G27));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n307), .A2(new_n719), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n304), .A2(KEYINPUT104), .A3(new_n306), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n720), .A2(new_n290), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n699), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  INV_X1    g538(.A(new_n567), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n563), .B(KEYINPUT103), .ZN(new_n726));
  AND2_X1   g540(.A1(new_n558), .A2(new_n565), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n725), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n467), .A3(new_n532), .A4(new_n533), .ZN(new_n729));
  NOR4_X1   g543(.A1(new_n723), .A2(new_n724), .A3(new_n667), .A4(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n304), .A2(new_n306), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n644), .B1(new_n282), .B2(new_n288), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n571), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n733), .A2(new_n729), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT42), .B1(new_n734), .B2(new_n669), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT105), .B1(new_n730), .B2(new_n735), .ZN(new_n736));
  AND2_X1   g550(.A1(new_n722), .A2(new_n699), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n729), .A2(new_n667), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n737), .A2(KEYINPUT42), .A3(new_n738), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n603), .A2(new_n604), .A3(new_n468), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n365), .A2(new_n740), .A3(new_n728), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n724), .B1(new_n741), .B2(new_n667), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT105), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n739), .A2(new_n742), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  XOR2_X1   g559(.A(KEYINPUT106), .B(G131), .Z(new_n746));
  XNOR2_X1  g560(.A(new_n745), .B(new_n746), .ZN(G33));
  NAND4_X1  g561(.A1(new_n365), .A2(new_n633), .A3(new_n740), .A4(new_n728), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT107), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G134), .ZN(G36));
  NAND2_X1  g565(.A1(new_n561), .A2(new_n562), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n561), .A2(KEYINPUT45), .A3(new_n562), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n565), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n757), .A2(new_n558), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(KEYINPUT108), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT108), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n757), .A2(new_n760), .A3(new_n558), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n756), .A2(new_n565), .ZN(new_n762));
  OAI211_X1 g576(.A(new_n759), .B(new_n761), .C1(new_n762), .C2(KEYINPUT46), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n763), .A2(new_n567), .A3(new_n657), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n576), .A2(new_n577), .ZN(new_n765));
  AND3_X1   g579(.A1(new_n581), .A2(new_n582), .A3(new_n584), .ZN(new_n766));
  AND2_X1   g580(.A1(new_n411), .A2(new_n412), .ZN(new_n767));
  OAI21_X1  g581(.A(new_n457), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT43), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT43), .ZN(new_n770));
  OAI211_X1 g584(.A(new_n770), .B(new_n457), .C1(new_n766), .C2(new_n767), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n765), .A2(new_n769), .A3(new_n617), .A4(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  AND2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n764), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n740), .B1(new_n772), .B2(new_n773), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n217), .ZN(G39));
  INV_X1    g592(.A(new_n740), .ZN(new_n779));
  NOR4_X1   g593(.A1(new_n779), .A2(new_n674), .A3(new_n571), .A4(new_n667), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n763), .A2(KEYINPUT47), .A3(new_n567), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  AOI21_X1  g596(.A(KEYINPUT47), .B1(new_n763), .B2(new_n567), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n780), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT109), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n763), .A2(new_n567), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n781), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n790), .A2(KEYINPUT109), .A3(new_n780), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n786), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  AND2_X1   g607(.A1(new_n676), .A2(new_n558), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OR2_X1    g609(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n698), .A2(new_n468), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(KEYINPUT49), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n567), .A4(new_n798), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n768), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n638), .A2(new_n641), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n801), .A3(new_n649), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n419), .A2(new_n631), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n740), .A2(KEYINPUT111), .A3(new_n597), .A4(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(KEYINPUT111), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n532), .A2(new_n467), .A3(new_n533), .A4(new_n597), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n807), .B1(new_n808), .B2(new_n804), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n806), .A2(new_n809), .A3(new_n628), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n738), .A2(new_n714), .ZN(new_n811));
  AOI21_X1  g625(.A(KEYINPUT107), .B1(new_n734), .B2(new_n633), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n733), .A2(new_n729), .A3(new_n749), .A4(new_n632), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n810), .B(new_n811), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  AND4_X1   g629(.A1(new_n571), .A2(new_n576), .A3(new_n568), .A4(new_n577), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n816), .A2(new_n534), .A3(new_n587), .A4(new_n601), .ZN(new_n817));
  AND3_X1   g631(.A1(new_n817), .A2(KEYINPUT110), .A3(new_n569), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT110), .B1(new_n817), .B2(new_n569), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n419), .A2(new_n650), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(new_n534), .A3(new_n601), .A4(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n622), .A2(new_n821), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n818), .A2(new_n819), .A3(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n652), .A2(new_n534), .A3(new_n631), .A4(new_n728), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n672), .A2(new_n634), .A3(new_n716), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n568), .B(new_n617), .C1(new_n731), .C2(new_n732), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n666), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n667), .B1(new_n711), .B2(new_n713), .ZN(new_n829));
  AOI22_X1  g643(.A1(new_n828), .A2(new_n633), .B1(new_n829), .B2(new_n715), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT52), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n830), .A2(new_n831), .A3(new_n672), .A4(new_n824), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n815), .A2(new_n823), .A3(new_n826), .A4(new_n832), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n702), .B1(new_n682), .B2(new_n684), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n692), .B1(new_n688), .B2(new_n679), .ZN(new_n835));
  INV_X1    g649(.A(new_n744), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n743), .B1(new_n739), .B2(new_n742), .ZN(new_n837));
  OAI211_X1 g651(.A(new_n834), .B(new_n835), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n803), .B1(new_n833), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n840));
  AND2_X1   g654(.A1(new_n826), .A2(new_n832), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n622), .A2(new_n821), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT110), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n733), .A2(new_n611), .A3(new_n465), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n605), .A2(new_n578), .A3(new_n680), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n817), .A2(new_n569), .A3(KEYINPUT110), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(new_n814), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n834), .A2(new_n835), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT53), .B1(new_n730), .B2(new_n735), .ZN(new_n852));
  INV_X1    g666(.A(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n841), .A2(new_n849), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n839), .A2(new_n840), .A3(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n850), .B1(new_n736), .B2(new_n744), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(KEYINPUT53), .A3(new_n849), .A4(new_n841), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n840), .B1(new_n839), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n855), .A2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT115), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n801), .A2(new_n468), .A3(new_n677), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(KEYINPUT113), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n769), .A2(new_n459), .A3(new_n771), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT112), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n769), .A2(KEYINPUT112), .A3(new_n459), .A4(new_n771), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n700), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT113), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n801), .A2(new_n868), .A3(new_n468), .A4(new_n677), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n862), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n862), .A2(new_n867), .A3(new_n869), .A4(KEYINPUT50), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n865), .A2(new_n866), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n779), .A2(new_n701), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n875), .A2(new_n714), .A3(new_n876), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT114), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n876), .A2(new_n571), .A3(new_n459), .A4(new_n649), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n585), .A2(new_n457), .A3(new_n586), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n881), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n860), .A2(new_n874), .A3(new_n878), .A4(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n881), .B1(new_n872), .B2(new_n873), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n860), .B1(new_n884), .B2(new_n878), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n795), .A2(new_n567), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n740), .B(new_n867), .C1(new_n790), .C2(new_n887), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n888), .A2(KEYINPUT51), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n875), .A2(new_n737), .A3(new_n876), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT116), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT48), .B1(new_n891), .B2(new_n892), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT48), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n335), .A2(G952), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n898), .B1(new_n867), .B2(new_n715), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n895), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n879), .A2(new_n680), .ZN(new_n901));
  OAI21_X1  g715(.A(KEYINPUT117), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  AND2_X1   g716(.A1(new_n897), .A2(new_n899), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT117), .ZN(new_n904));
  INV_X1    g718(.A(new_n901), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .A4(new_n895), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n902), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n884), .A2(new_n878), .A3(new_n888), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT51), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  AND4_X1   g724(.A1(new_n859), .A2(new_n890), .A3(new_n907), .A4(new_n910), .ZN(new_n911));
  NOR2_X1   g725(.A1(G952), .A2(G953), .ZN(new_n912));
  OAI21_X1  g726(.A(new_n802), .B1(new_n911), .B2(new_n912), .ZN(G75));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n839), .A2(new_n854), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n915), .A2(G902), .ZN(new_n916));
  INV_X1    g730(.A(G210), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n508), .B1(new_n515), .B2(new_n516), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(new_n474), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT55), .Z(new_n921));
  NAND2_X1  g735(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n335), .A2(G952), .ZN(new_n923));
  INV_X1    g737(.A(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(new_n921), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n914), .B(new_n925), .C1(new_n916), .C2(new_n917), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n922), .A2(new_n924), .A3(new_n926), .ZN(G51));
  XNOR2_X1  g741(.A(new_n675), .B(KEYINPUT118), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n840), .B1(new_n839), .B2(new_n854), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n855), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n564), .B(KEYINPUT57), .Z(new_n931));
  OAI21_X1  g745(.A(new_n928), .B1(new_n930), .B2(new_n931), .ZN(new_n932));
  OR2_X1    g746(.A1(new_n916), .A2(new_n756), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n923), .B1(new_n932), .B2(new_n933), .ZN(G54));
  NAND4_X1  g748(.A1(new_n915), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n935));
  INV_X1    g749(.A(new_n454), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n924), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n935), .A2(new_n936), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT119), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT119), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n935), .A2(new_n940), .A3(new_n936), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n937), .B1(new_n939), .B2(new_n941), .ZN(G60));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT59), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n944), .B1(new_n855), .B2(new_n858), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n581), .A2(new_n584), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n923), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n946), .B(new_n944), .C1(new_n855), .C2(new_n929), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT120), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n915), .A2(KEYINPUT54), .ZN(new_n952));
  NAND3_X1  g766(.A1(new_n839), .A2(new_n840), .A3(new_n854), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT120), .A3(new_n946), .A4(new_n944), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n948), .A2(new_n951), .A3(new_n955), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT121), .Z(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT60), .Z(new_n959));
  NAND2_X1  g773(.A1(new_n826), .A2(new_n832), .ZN(new_n960));
  NOR3_X1   g774(.A1(new_n960), .A2(new_n848), .A3(new_n814), .ZN(new_n961));
  AOI21_X1  g775(.A(KEYINPUT53), .B1(new_n961), .B2(new_n856), .ZN(new_n962));
  INV_X1    g776(.A(new_n854), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n614), .B(new_n959), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NOR4_X1   g780(.A1(new_n960), .A2(new_n848), .A3(new_n852), .A4(new_n814), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n841), .A2(new_n849), .A3(new_n745), .A4(new_n851), .ZN(new_n968));
  AOI22_X1  g782(.A1(new_n851), .A2(new_n967), .B1(new_n968), .B2(new_n803), .ZN(new_n969));
  INV_X1    g783(.A(new_n959), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n354), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n915), .A2(KEYINPUT122), .A3(new_n614), .A4(new_n959), .ZN(new_n972));
  NAND4_X1  g786(.A1(new_n966), .A2(new_n924), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n915), .A2(new_n959), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n923), .B1(new_n976), .B2(new_n354), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n977), .A2(new_n966), .A3(KEYINPUT61), .A4(new_n972), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n975), .A2(new_n978), .ZN(G66));
  NAND2_X1  g793(.A1(new_n851), .A2(new_n823), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(new_n335), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT123), .Z(new_n982));
  INV_X1    g796(.A(G224), .ZN(new_n983));
  OAI21_X1  g797(.A(G953), .B1(new_n462), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n919), .B1(G898), .B2(new_n335), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G69));
  AOI21_X1  g801(.A(new_n335), .B1(G227), .B2(G900), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n988), .B(KEYINPUT124), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n269), .A2(new_n273), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n991), .B(new_n448), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n335), .A2(G900), .ZN(new_n994));
  OAI21_X1  g808(.A(new_n993), .B1(KEYINPUT125), .B2(new_n994), .ZN(new_n995));
  OR2_X1    g809(.A1(new_n775), .A2(new_n776), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n792), .A2(new_n996), .ZN(new_n997));
  AND3_X1   g811(.A1(new_n672), .A2(new_n634), .A3(new_n716), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n723), .A2(new_n666), .A3(new_n651), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n999), .A2(new_n567), .A3(new_n657), .A4(new_n763), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n745), .A2(new_n750), .A3(new_n998), .A4(new_n1000), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n335), .B1(new_n997), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n994), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g818(.A(new_n995), .B1(new_n1004), .B2(KEYINPUT125), .ZN(new_n1005));
  NAND3_X1  g819(.A1(new_n662), .A2(new_n663), .A3(new_n998), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n662), .A2(KEYINPUT62), .A3(new_n663), .A4(new_n998), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n779), .A2(new_n658), .ZN(new_n1011));
  OAI211_X1 g825(.A(new_n1011), .B(new_n365), .C1(new_n587), .C2(new_n820), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n777), .B1(new_n786), .B2(new_n791), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n993), .A2(G953), .ZN(new_n1015));
  AND2_X1   g829(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI211_X1 g830(.A(KEYINPUT126), .B(new_n990), .C1(new_n1005), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(KEYINPUT126), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1000), .A2(new_n750), .A3(new_n998), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n1019), .B1(new_n736), .B2(new_n744), .ZN(new_n1020));
  AOI21_X1  g834(.A(G953), .B1(new_n1020), .B2(new_n1013), .ZN(new_n1021));
  OAI21_X1  g835(.A(KEYINPUT125), .B1(new_n1021), .B2(new_n994), .ZN(new_n1022));
  INV_X1    g836(.A(new_n995), .ZN(new_n1023));
  AOI22_X1  g837(.A1(new_n1022), .A2(new_n1023), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1024));
  OAI21_X1  g838(.A(new_n1018), .B1(new_n1024), .B2(new_n989), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1024), .A2(new_n988), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1017), .A2(new_n1025), .A3(new_n1026), .ZN(G72));
  NAND2_X1  g841(.A1(G472), .A2(G902), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT63), .Z(new_n1029));
  OAI21_X1  g843(.A(new_n1029), .B1(new_n1014), .B2(new_n980), .ZN(new_n1030));
  INV_X1    g844(.A(new_n645), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n923), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n839), .A2(new_n857), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n275), .A2(new_n266), .ZN(new_n1034));
  INV_X1    g848(.A(new_n1029), .ZN(new_n1035));
  NOR2_X1   g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1033), .A2(new_n645), .A3(new_n1036), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1037), .A2(KEYINPUT127), .ZN(new_n1038));
  INV_X1    g852(.A(KEYINPUT127), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n1033), .A2(new_n1039), .A3(new_n645), .A4(new_n1036), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1020), .A2(new_n1013), .ZN(new_n1042));
  OAI21_X1  g856(.A(new_n1029), .B1(new_n1042), .B2(new_n980), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1043), .A2(new_n1034), .ZN(new_n1044));
  AND3_X1   g858(.A1(new_n1032), .A2(new_n1041), .A3(new_n1044), .ZN(G57));
endmodule


