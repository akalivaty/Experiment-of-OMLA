

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584;

  INV_X1 U325 ( .A(KEYINPUT93), .ZN(n395) );
  NOR2_X1 U326 ( .A1(n413), .A2(n518), .ZN(n567) );
  XNOR2_X1 U327 ( .A(KEYINPUT98), .B(n468), .ZN(n518) );
  AND2_X1 U328 ( .A1(G232GAT), .A2(G233GAT), .ZN(n293) );
  AND2_X1 U329 ( .A1(G230GAT), .A2(G233GAT), .ZN(n294) );
  NOR2_X1 U330 ( .A1(n540), .A2(n365), .ZN(n366) );
  XNOR2_X1 U331 ( .A(n299), .B(n293), .ZN(n300) );
  XNOR2_X1 U332 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U333 ( .A(n425), .B(n294), .ZN(n347) );
  XNOR2_X1 U334 ( .A(n301), .B(n300), .ZN(n303) );
  XNOR2_X1 U335 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U336 ( .A(n347), .B(n378), .ZN(n348) );
  INV_X1 U337 ( .A(n406), .ZN(n407) );
  XNOR2_X1 U338 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U339 ( .A(n382), .B(n343), .ZN(n310) );
  XNOR2_X1 U340 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U341 ( .A(n355), .B(n354), .ZN(n359) );
  XNOR2_X1 U342 ( .A(n311), .B(n310), .ZN(n368) );
  XNOR2_X1 U343 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U344 ( .A(n557), .B(KEYINPUT76), .ZN(n545) );
  XNOR2_X1 U345 ( .A(n452), .B(n451), .ZN(n528) );
  XNOR2_X1 U346 ( .A(n454), .B(G190GAT), .ZN(n455) );
  XNOR2_X1 U347 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U348 ( .A(n456), .B(n455), .ZN(G1351GAT) );
  XNOR2_X1 U349 ( .A(n481), .B(n480), .ZN(G1330GAT) );
  XOR2_X1 U350 ( .A(KEYINPUT72), .B(KEYINPUT65), .Z(n296) );
  XOR2_X1 U351 ( .A(G50GAT), .B(G162GAT), .Z(n428) );
  XOR2_X1 U352 ( .A(G29GAT), .B(G134GAT), .Z(n405) );
  XNOR2_X1 U353 ( .A(n428), .B(n405), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n301) );
  XOR2_X1 U355 ( .A(KEYINPUT73), .B(KEYINPUT10), .Z(n298) );
  XNOR2_X1 U356 ( .A(KEYINPUT11), .B(KEYINPUT74), .ZN(n297) );
  XNOR2_X1 U357 ( .A(n298), .B(n297), .ZN(n299) );
  INV_X1 U358 ( .A(KEYINPUT9), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U360 ( .A(G92GAT), .B(G85GAT), .Z(n305) );
  XNOR2_X1 U361 ( .A(G99GAT), .B(G106GAT), .ZN(n304) );
  XNOR2_X1 U362 ( .A(n305), .B(n304), .ZN(n357) );
  XNOR2_X1 U363 ( .A(n357), .B(KEYINPUT75), .ZN(n306) );
  XNOR2_X1 U364 ( .A(n307), .B(n306), .ZN(n311) );
  XOR2_X1 U365 ( .A(G36GAT), .B(G190GAT), .Z(n308) );
  XOR2_X1 U366 ( .A(G218GAT), .B(n308), .Z(n382) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n309), .B(KEYINPUT7), .ZN(n343) );
  INV_X1 U369 ( .A(n368), .ZN(n557) );
  XNOR2_X1 U370 ( .A(KEYINPUT36), .B(n545), .ZN(n581) );
  XOR2_X1 U371 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n313) );
  XNOR2_X1 U372 ( .A(G57GAT), .B(KEYINPUT79), .ZN(n312) );
  XNOR2_X1 U373 ( .A(n313), .B(n312), .ZN(n328) );
  XOR2_X1 U374 ( .A(G1GAT), .B(G127GAT), .Z(n390) );
  XOR2_X1 U375 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n315) );
  NAND2_X1 U376 ( .A1(G231GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U377 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U378 ( .A(n390), .B(n316), .ZN(n326) );
  XOR2_X1 U379 ( .A(G71GAT), .B(KEYINPUT13), .Z(n349) );
  XOR2_X1 U380 ( .A(n349), .B(G211GAT), .Z(n318) );
  XOR2_X1 U381 ( .A(G22GAT), .B(G15GAT), .Z(n342) );
  XNOR2_X1 U382 ( .A(n342), .B(G155GAT), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U384 ( .A(KEYINPUT12), .B(G64GAT), .Z(n320) );
  XNOR2_X1 U385 ( .A(G8GAT), .B(KEYINPUT80), .ZN(n319) );
  XNOR2_X1 U386 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U387 ( .A(n322), .B(n321), .Z(n324) );
  XNOR2_X1 U388 ( .A(G183GAT), .B(G78GAT), .ZN(n323) );
  XNOR2_X1 U389 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n577) );
  NOR2_X1 U392 ( .A1(n581), .A2(n577), .ZN(n329) );
  XNOR2_X1 U393 ( .A(n329), .B(KEYINPUT45), .ZN(n361) );
  XOR2_X1 U394 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n331) );
  NAND2_X1 U395 ( .A1(G229GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U396 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U397 ( .A(n332), .B(KEYINPUT66), .Z(n340) );
  XOR2_X1 U398 ( .A(G197GAT), .B(G36GAT), .Z(n334) );
  XNOR2_X1 U399 ( .A(G50GAT), .B(G29GAT), .ZN(n333) );
  XNOR2_X1 U400 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U401 ( .A(KEYINPUT30), .B(G1GAT), .Z(n336) );
  XNOR2_X1 U402 ( .A(G141GAT), .B(G113GAT), .ZN(n335) );
  XNOR2_X1 U403 ( .A(n336), .B(n335), .ZN(n337) );
  XNOR2_X1 U404 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U406 ( .A(G169GAT), .B(G8GAT), .Z(n375) );
  XOR2_X1 U407 ( .A(n341), .B(n375), .Z(n345) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U409 ( .A(n345), .B(n344), .ZN(n568) );
  XOR2_X1 U410 ( .A(KEYINPUT69), .B(G78GAT), .Z(n425) );
  XNOR2_X1 U411 ( .A(G176GAT), .B(G204GAT), .ZN(n346) );
  XNOR2_X1 U412 ( .A(n346), .B(G64GAT), .ZN(n378) );
  XNOR2_X1 U413 ( .A(n348), .B(KEYINPUT33), .ZN(n355) );
  XOR2_X1 U414 ( .A(n349), .B(KEYINPUT71), .Z(n353) );
  XOR2_X1 U415 ( .A(KEYINPUT70), .B(KEYINPUT68), .Z(n351) );
  XNOR2_X1 U416 ( .A(KEYINPUT32), .B(KEYINPUT31), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U418 ( .A(G120GAT), .B(G148GAT), .ZN(n356) );
  XNOR2_X1 U419 ( .A(n356), .B(G57GAT), .ZN(n406) );
  XOR2_X1 U420 ( .A(n406), .B(n357), .Z(n358) );
  XNOR2_X1 U421 ( .A(n359), .B(n358), .ZN(n573) );
  AND2_X1 U422 ( .A1(n568), .A2(n573), .ZN(n360) );
  AND2_X1 U423 ( .A1(n361), .A2(n360), .ZN(n362) );
  XOR2_X1 U424 ( .A(n362), .B(KEYINPUT113), .Z(n371) );
  INV_X1 U425 ( .A(n577), .ZN(n540) );
  XOR2_X1 U426 ( .A(KEYINPUT64), .B(KEYINPUT41), .Z(n363) );
  XNOR2_X1 U427 ( .A(n573), .B(n363), .ZN(n551) );
  NOR2_X1 U428 ( .A1(n568), .A2(n551), .ZN(n364) );
  XNOR2_X1 U429 ( .A(n364), .B(KEYINPUT46), .ZN(n365) );
  XOR2_X1 U430 ( .A(KEYINPUT112), .B(n366), .Z(n367) );
  NOR2_X1 U431 ( .A1(n368), .A2(n367), .ZN(n369) );
  XOR2_X1 U432 ( .A(KEYINPUT47), .B(n369), .Z(n370) );
  NOR2_X1 U433 ( .A1(n371), .A2(n370), .ZN(n372) );
  XNOR2_X1 U434 ( .A(KEYINPUT48), .B(n372), .ZN(n526) );
  XOR2_X1 U435 ( .A(G183GAT), .B(KEYINPUT17), .Z(n374) );
  XNOR2_X1 U436 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n373) );
  XNOR2_X1 U437 ( .A(n374), .B(n373), .ZN(n434) );
  XOR2_X1 U438 ( .A(G92GAT), .B(n375), .Z(n377) );
  NAND2_X1 U439 ( .A1(G226GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U440 ( .A(n377), .B(n376), .ZN(n379) );
  XOR2_X1 U441 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U442 ( .A(G211GAT), .B(KEYINPUT21), .Z(n381) );
  XNOR2_X1 U443 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n380) );
  XNOR2_X1 U444 ( .A(n381), .B(n380), .ZN(n427) );
  XNOR2_X1 U445 ( .A(n427), .B(n382), .ZN(n383) );
  XNOR2_X1 U446 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U447 ( .A(n434), .B(n385), .ZN(n457) );
  NOR2_X1 U448 ( .A1(n526), .A2(n457), .ZN(n386) );
  XOR2_X1 U449 ( .A(n386), .B(KEYINPUT54), .Z(n413) );
  XOR2_X1 U450 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n388) );
  XNOR2_X1 U451 ( .A(KEYINPUT4), .B(KEYINPUT95), .ZN(n387) );
  XNOR2_X1 U452 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U453 ( .A(n389), .B(G85GAT), .Z(n392) );
  XNOR2_X1 U454 ( .A(G162GAT), .B(n390), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n412) );
  XOR2_X1 U456 ( .A(KEYINPUT92), .B(KEYINPUT1), .Z(n394) );
  XNOR2_X1 U457 ( .A(KEYINPUT6), .B(KEYINPUT94), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n398) );
  NAND2_X1 U459 ( .A1(G225GAT), .A2(G233GAT), .ZN(n396) );
  XOR2_X1 U460 ( .A(n399), .B(KEYINPUT97), .Z(n404) );
  XOR2_X1 U461 ( .A(KEYINPUT89), .B(KEYINPUT3), .Z(n401) );
  XNOR2_X1 U462 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U464 ( .A(G141GAT), .B(n402), .Z(n432) );
  XNOR2_X1 U465 ( .A(n432), .B(KEYINPUT91), .ZN(n403) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n410) );
  XOR2_X1 U467 ( .A(G113GAT), .B(KEYINPUT0), .Z(n446) );
  XNOR2_X1 U468 ( .A(n405), .B(n446), .ZN(n408) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n468) );
  XOR2_X1 U470 ( .A(G148GAT), .B(G204GAT), .Z(n415) );
  XNOR2_X1 U471 ( .A(G218GAT), .B(G106GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U473 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n417) );
  XNOR2_X1 U474 ( .A(G22GAT), .B(KEYINPUT22), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n418) );
  XOR2_X1 U476 ( .A(n419), .B(n418), .Z(n424) );
  XOR2_X1 U477 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n421) );
  NAND2_X1 U478 ( .A1(G228GAT), .A2(G233GAT), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U480 ( .A(KEYINPUT90), .B(n422), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n426) );
  XOR2_X1 U482 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U485 ( .A(n432), .B(n431), .ZN(n463) );
  NAND2_X1 U486 ( .A1(n567), .A2(n463), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n433), .B(KEYINPUT55), .ZN(n453) );
  XOR2_X1 U488 ( .A(G169GAT), .B(n434), .Z(n436) );
  NAND2_X1 U489 ( .A1(G227GAT), .A2(G233GAT), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n452) );
  XOR2_X1 U491 ( .A(G71GAT), .B(G176GAT), .Z(n438) );
  XNOR2_X1 U492 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n437) );
  XNOR2_X1 U493 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U494 ( .A(G127GAT), .B(G120GAT), .Z(n440) );
  XNOR2_X1 U495 ( .A(G15GAT), .B(KEYINPUT82), .ZN(n439) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U497 ( .A(n442), .B(n441), .ZN(n450) );
  XOR2_X1 U498 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n444) );
  XNOR2_X1 U499 ( .A(G99GAT), .B(G134GAT), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U501 ( .A(n445), .B(G190GAT), .Z(n448) );
  XNOR2_X1 U502 ( .A(G43GAT), .B(n446), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n451) );
  NAND2_X1 U505 ( .A1(n453), .A2(n528), .ZN(n562) );
  NOR2_X1 U506 ( .A1(n545), .A2(n562), .ZN(n456) );
  XNOR2_X1 U507 ( .A(KEYINPUT121), .B(KEYINPUT58), .ZN(n454) );
  INV_X1 U508 ( .A(n457), .ZN(n520) );
  XOR2_X1 U509 ( .A(KEYINPUT27), .B(KEYINPUT99), .Z(n458) );
  XNOR2_X1 U510 ( .A(n520), .B(n458), .ZN(n465) );
  NAND2_X1 U511 ( .A1(n465), .A2(n518), .ZN(n459) );
  XNOR2_X1 U512 ( .A(n459), .B(KEYINPUT100), .ZN(n527) );
  NOR2_X1 U513 ( .A1(n528), .A2(n527), .ZN(n460) );
  XNOR2_X1 U514 ( .A(KEYINPUT28), .B(n463), .ZN(n497) );
  NAND2_X1 U515 ( .A1(n460), .A2(n497), .ZN(n472) );
  NAND2_X1 U516 ( .A1(n520), .A2(n528), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n463), .A2(n461), .ZN(n462) );
  XNOR2_X1 U518 ( .A(n462), .B(KEYINPUT25), .ZN(n467) );
  NOR2_X1 U519 ( .A1(n528), .A2(n463), .ZN(n464) );
  XNOR2_X1 U520 ( .A(KEYINPUT26), .B(n464), .ZN(n566) );
  AND2_X1 U521 ( .A1(n465), .A2(n566), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n469) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n470) );
  XNOR2_X1 U524 ( .A(KEYINPUT101), .B(n470), .ZN(n471) );
  NAND2_X1 U525 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U526 ( .A(KEYINPUT102), .B(n473), .Z(n487) );
  NOR2_X1 U527 ( .A1(n540), .A2(n487), .ZN(n474) );
  XNOR2_X1 U528 ( .A(n474), .B(KEYINPUT105), .ZN(n475) );
  NOR2_X1 U529 ( .A1(n581), .A2(n475), .ZN(n476) );
  XNOR2_X1 U530 ( .A(KEYINPUT37), .B(n476), .ZN(n517) );
  INV_X1 U531 ( .A(n568), .ZN(n532) );
  NAND2_X1 U532 ( .A1(n573), .A2(n532), .ZN(n489) );
  NOR2_X1 U533 ( .A1(n517), .A2(n489), .ZN(n477) );
  XNOR2_X1 U534 ( .A(KEYINPUT38), .B(n477), .ZN(n503) );
  NAND2_X1 U535 ( .A1(n503), .A2(n528), .ZN(n481) );
  XOR2_X1 U536 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n479) );
  XNOR2_X1 U537 ( .A(G43GAT), .B(KEYINPUT106), .ZN(n478) );
  XNOR2_X1 U538 ( .A(KEYINPUT108), .B(n551), .ZN(n535) );
  NOR2_X1 U539 ( .A1(n535), .A2(n562), .ZN(n484) );
  XNOR2_X1 U540 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n482), .B(G176GAT), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT81), .B(KEYINPUT16), .Z(n486) );
  NAND2_X1 U544 ( .A1(n545), .A2(n540), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n488) );
  OR2_X1 U546 ( .A1(n488), .A2(n487), .ZN(n505) );
  NOR2_X1 U547 ( .A1(n489), .A2(n505), .ZN(n490) );
  XOR2_X1 U548 ( .A(KEYINPUT103), .B(n490), .Z(n498) );
  NAND2_X1 U549 ( .A1(n498), .A2(n518), .ZN(n493) );
  XNOR2_X1 U550 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n491) );
  XNOR2_X1 U551 ( .A(n491), .B(KEYINPUT104), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(G1324GAT) );
  NAND2_X1 U553 ( .A1(n498), .A2(n520), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n494), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(G15GAT), .B(KEYINPUT35), .Z(n496) );
  NAND2_X1 U556 ( .A1(n498), .A2(n528), .ZN(n495) );
  XNOR2_X1 U557 ( .A(n496), .B(n495), .ZN(G1326GAT) );
  INV_X1 U558 ( .A(n497), .ZN(n531) );
  NAND2_X1 U559 ( .A1(n531), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U561 ( .A(G29GAT), .B(KEYINPUT39), .Z(n501) );
  NAND2_X1 U562 ( .A1(n503), .A2(n518), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(G1328GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n520), .ZN(n502) );
  XNOR2_X1 U565 ( .A(n502), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U566 ( .A1(n531), .A2(n503), .ZN(n504) );
  XNOR2_X1 U567 ( .A(G50GAT), .B(n504), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n508) );
  OR2_X1 U569 ( .A1(n532), .A2(n535), .ZN(n516) );
  NOR2_X1 U570 ( .A1(n516), .A2(n505), .ZN(n506) );
  XOR2_X1 U571 ( .A(KEYINPUT109), .B(n506), .Z(n512) );
  NAND2_X1 U572 ( .A1(n512), .A2(n518), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U574 ( .A(G57GAT), .B(n509), .Z(G1332GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n520), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n528), .A2(n512), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT111), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U580 ( .A1(n512), .A2(n531), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(n515) );
  XOR2_X1 U582 ( .A(G78GAT), .B(n515), .Z(G1335GAT) );
  NOR2_X1 U583 ( .A1(n517), .A2(n516), .ZN(n523) );
  NAND2_X1 U584 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U585 ( .A(n519), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n523), .A2(n520), .ZN(n521) );
  XNOR2_X1 U587 ( .A(n521), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n528), .A2(n523), .ZN(n522) );
  XNOR2_X1 U589 ( .A(n522), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n531), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n524), .B(KEYINPUT44), .ZN(n525) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n525), .ZN(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT115), .Z(n534) );
  NOR2_X1 U594 ( .A1(n527), .A2(n526), .ZN(n548) );
  NAND2_X1 U595 ( .A1(n548), .A2(n528), .ZN(n529) );
  XNOR2_X1 U596 ( .A(KEYINPUT114), .B(n529), .ZN(n530) );
  NOR2_X1 U597 ( .A1(n531), .A2(n530), .ZN(n541) );
  NAND2_X1 U598 ( .A1(n541), .A2(n532), .ZN(n533) );
  XNOR2_X1 U599 ( .A(n534), .B(n533), .ZN(G1340GAT) );
  INV_X1 U600 ( .A(n541), .ZN(n544) );
  NOR2_X1 U601 ( .A1(n544), .A2(n535), .ZN(n539) );
  XOR2_X1 U602 ( .A(KEYINPUT116), .B(KEYINPUT117), .Z(n537) );
  XNOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1341GAT) );
  NAND2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U607 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U608 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  NOR2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n547) );
  XNOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U611 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U612 ( .A1(n548), .A2(n566), .ZN(n558) );
  NOR2_X1 U613 ( .A1(n568), .A2(n558), .ZN(n549) );
  XOR2_X1 U614 ( .A(G141GAT), .B(n549), .Z(n550) );
  XNOR2_X1 U615 ( .A(KEYINPUT118), .B(n550), .ZN(G1344GAT) );
  NOR2_X1 U616 ( .A1(n551), .A2(n558), .ZN(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NOR2_X1 U620 ( .A1(n577), .A2(n558), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1346GAT) );
  NOR2_X1 U623 ( .A1(n557), .A2(n558), .ZN(n559) );
  XOR2_X1 U624 ( .A(KEYINPUT120), .B(n559), .Z(n560) );
  XNOR2_X1 U625 ( .A(G162GAT), .B(n560), .ZN(G1347GAT) );
  NOR2_X1 U626 ( .A1(n568), .A2(n562), .ZN(n561) );
  XOR2_X1 U627 ( .A(G169GAT), .B(n561), .Z(G1348GAT) );
  NOR2_X1 U628 ( .A1(n577), .A2(n562), .ZN(n563) );
  XOR2_X1 U629 ( .A(G183GAT), .B(n563), .Z(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U631 ( .A(KEYINPUT59), .B(KEYINPUT60), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n580) );
  NOR2_X1 U634 ( .A1(n568), .A2(n580), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT122), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n580), .ZN(n575) );
  XNOR2_X1 U639 ( .A(KEYINPUT125), .B(KEYINPUT61), .ZN(n574) );
  XNOR2_X1 U640 ( .A(n575), .B(n574), .ZN(n576) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n576), .Z(G1353GAT) );
  NOR2_X1 U642 ( .A1(n577), .A2(n580), .ZN(n578) );
  XOR2_X1 U643 ( .A(KEYINPUT126), .B(n578), .Z(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

