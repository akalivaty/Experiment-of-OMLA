//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 0 0 1 0 0 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:15 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n771, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n866, new_n867, new_n868, new_n870,
    new_n871, new_n872, new_n874, new_n875, new_n876, new_n877, new_n878,
    new_n879, new_n880, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n995,
    new_n996;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  XOR2_X1   g001(.A(G127gat), .B(G134gat), .Z(new_n203));
  XNOR2_X1  g002(.A(G113gat), .B(G120gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(KEYINPUT1), .B2(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G113gat), .B(G120gat), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT1), .ZN(new_n207));
  XNOR2_X1  g006(.A(G127gat), .B(G134gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n206), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n205), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT69), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n212), .A2(new_n213), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n215), .A2(KEYINPUT23), .A3(new_n216), .ZN(new_n217));
  NAND2_X1  g016(.A1(G169gat), .A2(G176gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(KEYINPUT25), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(G169gat), .A2(G176gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT23), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n217), .B(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  NAND3_X1  g022(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(G183gat), .B2(G190gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(G183gat), .A2(G190gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT24), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT68), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n232));
  AOI21_X1  g031(.A(new_n225), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n223), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT23), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT66), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT66), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT23), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n221), .B1(new_n236), .B2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n218), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NOR2_X1   g041(.A1(G183gat), .A2(G190gat), .ZN(new_n243));
  AND2_X1   g042(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n243), .B1(new_n244), .B2(G190gat), .ZN(new_n245));
  AND3_X1   g044(.A1(new_n226), .A2(KEYINPUT65), .A3(new_n227), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT65), .B1(new_n226), .B2(new_n227), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  AOI21_X1  g047(.A(KEYINPUT25), .B1(new_n242), .B2(new_n248), .ZN(new_n249));
  OAI21_X1  g048(.A(new_n211), .B1(new_n234), .B2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT25), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n231), .A2(KEYINPUT65), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n225), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n218), .B(new_n240), .C1(new_n222), .C2(new_n221), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n251), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n228), .A2(new_n229), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n231), .A2(KEYINPUT68), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n245), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n239), .A2(new_n219), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n260), .A2(new_n261), .A3(new_n217), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT69), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n250), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT26), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n218), .B1(new_n221), .B2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n215), .A2(new_n265), .A3(new_n216), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(KEYINPUT70), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT70), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n215), .A2(new_n269), .A3(new_n265), .A4(new_n216), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n266), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(KEYINPUT27), .B(G183gat), .ZN(new_n272));
  INV_X1    g071(.A(G190gat), .ZN(new_n273));
  AOI21_X1  g072(.A(KEYINPUT28), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G183gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(KEYINPUT27), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT27), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(G183gat), .ZN(new_n278));
  AND4_X1   g077(.A1(KEYINPUT28), .A2(new_n276), .A3(new_n278), .A4(new_n273), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n226), .B1(new_n274), .B2(new_n279), .ZN(new_n280));
  OR2_X1    g079(.A1(new_n271), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n210), .B1(new_n264), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n205), .A2(new_n209), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n271), .A2(new_n280), .ZN(new_n284));
  AOI211_X1 g083(.A(new_n283), .B(new_n284), .C1(new_n250), .C2(new_n263), .ZN(new_n285));
  NOR2_X1   g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT34), .ZN(new_n287));
  NAND2_X1  g086(.A1(G227gat), .A2(G233gat), .ZN(new_n288));
  XNOR2_X1  g087(.A(new_n288), .B(KEYINPUT64), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n286), .A2(KEYINPUT72), .A3(new_n287), .A4(new_n290), .ZN(new_n291));
  AND3_X1   g090(.A1(new_n257), .A2(KEYINPUT69), .A3(new_n262), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT69), .B1(new_n257), .B2(new_n262), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n281), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(new_n283), .ZN(new_n295));
  NAND3_X1  g094(.A1(new_n264), .A2(new_n210), .A3(new_n281), .ZN(new_n296));
  NAND4_X1  g095(.A1(new_n295), .A2(new_n287), .A3(new_n290), .A4(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n290), .A3(new_n296), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT71), .A3(KEYINPUT34), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g102(.A(KEYINPUT71), .B1(new_n301), .B2(KEYINPUT34), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n300), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n289), .B1(new_n282), .B2(new_n285), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n306), .A2(KEYINPUT32), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT33), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  XOR2_X1   g108(.A(G15gat), .B(G43gat), .Z(new_n310));
  XNOR2_X1  g109(.A(G71gat), .B(G99gat), .ZN(new_n311));
  XNOR2_X1  g110(.A(new_n310), .B(new_n311), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n307), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(new_n312), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n306), .B(KEYINPUT32), .C1(new_n308), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n305), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n301), .A2(KEYINPUT34), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n302), .ZN(new_n321));
  AOI22_X1  g120(.A1(new_n321), .A2(new_n300), .B1(new_n313), .B2(new_n315), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n202), .B1(new_n317), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(G228gat), .A2(G233gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(G197gat), .B(G204gat), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT22), .ZN(new_n326));
  INV_X1    g125(.A(G211gat), .ZN(new_n327));
  INV_X1    g126(.A(G218gat), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G211gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n331), .A2(new_n325), .A3(new_n329), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT29), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT3), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(G141gat), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(G148gat), .ZN(new_n341));
  INV_X1    g140(.A(G148gat), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(G141gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT2), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G155gat), .ZN(new_n347));
  INV_X1    g146(.A(G162gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G155gat), .A2(G162gat), .ZN(new_n350));
  AND2_X1   g149(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n341), .A2(KEYINPUT75), .ZN(new_n353));
  XNOR2_X1  g152(.A(KEYINPUT74), .B(G148gat), .ZN(new_n354));
  AOI21_X1  g153(.A(new_n353), .B1(new_n354), .B2(G141gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n342), .A2(KEYINPUT74), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT74), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(G148gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT75), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n356), .A2(new_n358), .A3(new_n359), .A4(G141gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n350), .B1(new_n349), .B2(KEYINPUT2), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n352), .B1(new_n355), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n324), .B1(new_n339), .B2(new_n363), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n352), .B(new_n338), .C1(new_n355), .C2(new_n362), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n336), .ZN(new_n366));
  INV_X1    g165(.A(new_n335), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT3), .B1(new_n335), .B2(new_n336), .ZN(new_n369));
  INV_X1    g168(.A(new_n363), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT81), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(KEYINPUT81), .ZN(new_n372));
  AOI21_X1  g171(.A(KEYINPUT29), .B1(new_n333), .B2(new_n334), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n372), .B(new_n363), .C1(new_n373), .C2(KEYINPUT3), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n371), .A2(new_n368), .A3(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n324), .B(KEYINPUT80), .Z(new_n376));
  AOI221_X4 g175(.A(G22gat), .B1(new_n364), .B2(new_n368), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G22gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n376), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n368), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n378), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  XNOR2_X1  g180(.A(G78gat), .B(G106gat), .ZN(new_n382));
  INV_X1    g181(.A(G50gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(new_n382), .B(new_n383), .ZN(new_n384));
  XOR2_X1   g183(.A(KEYINPUT79), .B(KEYINPUT31), .Z(new_n385));
  XNOR2_X1  g184(.A(new_n384), .B(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n386), .ZN(new_n387));
  NOR4_X1   g186(.A1(new_n377), .A2(new_n381), .A3(KEYINPUT82), .A4(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n377), .A2(new_n381), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT82), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n386), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  OAI21_X1  g190(.A(KEYINPUT82), .B1(new_n377), .B2(new_n381), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n388), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n305), .A2(new_n316), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n321), .A2(new_n313), .A3(new_n315), .A4(new_n300), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT85), .ZN(new_n396));
  INV_X1    g195(.A(G226gat), .ZN(new_n397));
  INV_X1    g196(.A(G233gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n257), .A2(new_n262), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n281), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n284), .B1(new_n250), .B2(new_n263), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n399), .A2(KEYINPUT29), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n367), .B(new_n401), .C1(new_n402), .C2(new_n404), .ZN(new_n405));
  XNOR2_X1  g204(.A(G8gat), .B(G36gat), .ZN(new_n406));
  XNOR2_X1  g205(.A(G64gat), .B(G92gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  AOI21_X1  g207(.A(new_n404), .B1(new_n281), .B2(new_n400), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n409), .B1(new_n402), .B2(new_n399), .ZN(new_n410));
  OAI211_X1 g209(.A(new_n405), .B(new_n408), .C1(new_n410), .C2(new_n367), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT30), .ZN(new_n412));
  INV_X1    g211(.A(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(new_n399), .ZN(new_n414));
  AOI211_X1 g213(.A(new_n414), .B(new_n284), .C1(new_n250), .C2(new_n263), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n335), .B1(new_n415), .B2(new_n409), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT73), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n416), .A2(new_n417), .A3(new_n405), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n416), .B2(new_n405), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n413), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  XOR2_X1   g220(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n422));
  NAND3_X1  g221(.A1(new_n412), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n363), .A2(KEYINPUT3), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n424), .A2(new_n365), .A3(new_n283), .ZN(new_n425));
  NAND2_X1  g224(.A1(G225gat), .A2(G233gat), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT4), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n427), .B1(new_n363), .B2(new_n283), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n356), .A2(new_n358), .A3(G141gat), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n429), .A2(KEYINPUT75), .A3(new_n341), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n430), .A2(new_n360), .A3(new_n361), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n210), .A2(KEYINPUT4), .A3(new_n431), .A4(new_n352), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n425), .A2(new_n426), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT5), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n363), .A2(new_n283), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n431), .A2(new_n352), .A3(new_n209), .A4(new_n205), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n426), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n433), .A2(new_n439), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n428), .A2(new_n432), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n441), .A2(new_n434), .A3(new_n426), .A4(new_n425), .ZN(new_n442));
  XOR2_X1   g241(.A(G1gat), .B(G29gat), .Z(new_n443));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  XNOR2_X1  g244(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n445), .B(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n440), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT77), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n440), .A2(new_n442), .ZN(new_n451));
  INV_X1    g250(.A(new_n447), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n440), .A2(new_n442), .A3(KEYINPUT77), .A4(new_n447), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n450), .A2(new_n453), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n447), .B1(new_n440), .B2(new_n442), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT6), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(KEYINPUT84), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT84), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n457), .A2(new_n460), .A3(KEYINPUT6), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n456), .A2(new_n459), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n423), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g262(.A1(new_n323), .A2(new_n393), .A3(new_n396), .A4(new_n463), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n393), .A2(new_n395), .A3(new_n394), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT30), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n411), .B(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n416), .A2(new_n405), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n468), .A2(KEYINPUT73), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n408), .B1(new_n469), .B2(new_n418), .ZN(new_n470));
  NOR2_X1   g269(.A1(new_n467), .A2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT78), .ZN(new_n472));
  XNOR2_X1  g271(.A(new_n457), .B(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n450), .A2(new_n454), .A3(new_n455), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n458), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n471), .A2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(KEYINPUT35), .B1(new_n465), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n464), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT36), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n479), .B1(new_n317), .B2(new_n322), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n394), .A2(new_n395), .A3(KEYINPUT36), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n441), .A2(new_n425), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n483), .A2(new_n438), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n484), .B(KEYINPUT39), .C1(new_n438), .C2(new_n437), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT39), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n486), .A3(new_n438), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n485), .A2(new_n447), .A3(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(KEYINPUT83), .A2(KEYINPUT40), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n457), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(new_n489), .ZN(new_n491));
  NAND4_X1  g290(.A1(new_n485), .A2(new_n447), .A3(new_n491), .A4(new_n487), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n490), .B(new_n492), .C1(new_n470), .C2(new_n467), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT37), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n416), .A2(new_n494), .A3(new_n405), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n335), .B(new_n401), .C1(new_n402), .C2(new_n404), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(KEYINPUT37), .C1(new_n410), .C2(new_n335), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT38), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n495), .A2(new_n497), .A3(new_n498), .A4(new_n413), .ZN(new_n499));
  AND2_X1   g298(.A1(new_n499), .A2(new_n411), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n462), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT37), .B1(new_n419), .B2(new_n420), .ZN(new_n502));
  AND2_X1   g301(.A1(new_n495), .A2(new_n413), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI211_X1 g303(.A(new_n493), .B(new_n393), .C1(new_n501), .C2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n391), .A2(new_n392), .ZN(new_n506));
  INV_X1    g305(.A(new_n388), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n476), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n482), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n478), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  OR2_X1    g311(.A1(new_n512), .A2(G1gat), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT16), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n514), .B2(G1gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n513), .A2(KEYINPUT88), .ZN(new_n517));
  INV_X1    g316(.A(G8gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n513), .B(new_n515), .C1(KEYINPUT88), .C2(G8gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT89), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(KEYINPUT89), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(G71gat), .A2(G78gat), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n526), .A2(KEYINPUT9), .ZN(new_n527));
  NAND2_X1  g326(.A1(G71gat), .A2(G78gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  XOR2_X1   g328(.A(G57gat), .B(G64gat), .Z(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT92), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT92), .ZN(new_n534));
  XNOR2_X1  g333(.A(G57gat), .B(G64gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT91), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(G57gat), .A2(G64gat), .ZN(new_n538));
  NAND2_X1  g337(.A1(G57gat), .A2(G64gat), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n538), .A2(KEYINPUT91), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n537), .A2(KEYINPUT9), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(new_n528), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n542), .A2(new_n526), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n533), .A2(new_n534), .B1(new_n541), .B2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT21), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n525), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT95), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n525), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  AND3_X1   g350(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n551), .B1(new_n547), .B2(new_n549), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n533), .A2(new_n534), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n541), .A2(new_n543), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g356(.A(KEYINPUT93), .B(KEYINPUT21), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(G231gat), .A2(G233gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n557), .A2(new_n560), .A3(new_n558), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G127gat), .B(G155gat), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n565), .B(KEYINPUT94), .Z(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n562), .A2(new_n568), .A3(new_n563), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  XOR2_X1   g369(.A(G183gat), .B(G211gat), .Z(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n571), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n567), .A2(new_n573), .A3(new_n569), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n554), .A2(new_n572), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n572), .A2(new_n574), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n576), .B1(new_n552), .B2(new_n553), .ZN(new_n577));
  AND2_X1   g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G43gat), .B(G50gat), .Z(new_n579));
  INV_X1    g378(.A(G36gat), .ZN(new_n580));
  AND2_X1   g379(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n581));
  NOR2_X1   g380(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G29gat), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n584), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n579), .B1(new_n586), .B2(KEYINPUT15), .ZN(new_n587));
  INV_X1    g386(.A(KEYINPUT15), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n583), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n586), .A2(KEYINPUT15), .A3(new_n579), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n590), .A2(KEYINPUT17), .A3(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(G99gat), .A2(G106gat), .ZN(new_n593));
  NAND2_X1  g392(.A1(G99gat), .A2(G106gat), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(G85gat), .A2(G92gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n596), .B(KEYINPUT7), .ZN(new_n597));
  INV_X1    g396(.A(G85gat), .ZN(new_n598));
  INV_X1    g397(.A(G92gat), .ZN(new_n599));
  AOI22_X1  g398(.A1(KEYINPUT8), .A2(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n595), .B1(new_n597), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n597), .A2(new_n595), .A3(new_n600), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n590), .A2(new_n591), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT87), .B(KEYINPUT17), .ZN(new_n606));
  OAI211_X1 g405(.A(new_n592), .B(new_n604), .C1(new_n605), .C2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n591), .ZN(new_n608));
  AND3_X1   g407(.A1(new_n597), .A2(new_n595), .A3(new_n600), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n601), .ZN(new_n610));
  AND2_X1   g409(.A1(G232gat), .A2(G233gat), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n608), .A2(new_n610), .B1(KEYINPUT41), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(G190gat), .B(G218gat), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n614), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n607), .A2(new_n616), .A3(new_n612), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n611), .A2(KEYINPUT41), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n615), .A2(new_n617), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n624), .B(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n615), .A2(new_n627), .A3(new_n617), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n607), .A2(KEYINPUT98), .A3(new_n616), .A4(new_n612), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n626), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT105), .ZN(new_n633));
  XOR2_X1   g432(.A(G120gat), .B(G148gat), .Z(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT103), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT100), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n557), .A2(new_n639), .A3(new_n604), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT100), .B1(new_n544), .B2(new_n610), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n609), .B1(new_n642), .B2(new_n601), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n602), .A2(KEYINPUT101), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n643), .A2(new_n544), .A3(new_n644), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n640), .A2(new_n641), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT102), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n646), .A2(KEYINPUT102), .A3(new_n648), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  XOR2_X1   g452(.A(new_n647), .B(KEYINPUT104), .Z(new_n654));
  INV_X1    g453(.A(KEYINPUT10), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n640), .A2(new_n641), .A3(new_n645), .A4(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n544), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n654), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n638), .B1(new_n653), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n648), .B1(new_n656), .B2(new_n657), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND4_X1  g460(.A1(new_n661), .A2(new_n652), .A3(new_n651), .A4(new_n637), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n578), .A2(new_n632), .A3(new_n633), .A4(new_n664), .ZN(new_n665));
  NAND4_X1  g464(.A1(new_n575), .A2(new_n577), .A3(new_n630), .A4(new_n626), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT105), .B1(new_n666), .B2(new_n663), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n523), .A2(new_n608), .A3(new_n524), .ZN(new_n668));
  OAI211_X1 g467(.A(new_n521), .B(new_n592), .C1(new_n605), .C2(new_n606), .ZN(new_n669));
  NAND2_X1  g468(.A1(G229gat), .A2(G233gat), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n668), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT18), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(KEYINPUT90), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g472(.A(new_n670), .B(KEYINPUT13), .Z(new_n674));
  INV_X1    g473(.A(new_n668), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n608), .B1(new_n523), .B2(new_n524), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n672), .A2(KEYINPUT90), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n668), .A2(new_n669), .A3(new_n670), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n673), .A2(new_n677), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g479(.A(G113gat), .B(G141gat), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G197gat), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT11), .B(G169gat), .Z(new_n683));
  XNOR2_X1  g482(.A(new_n682), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(KEYINPUT12), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n680), .A2(new_n686), .ZN(new_n687));
  NAND4_X1  g486(.A1(new_n673), .A2(new_n677), .A3(new_n685), .A4(new_n679), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AND3_X1   g488(.A1(new_n665), .A2(new_n667), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n511), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n475), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(G1gat), .ZN(G1324gat));
  INV_X1    g494(.A(new_n471), .ZN(new_n696));
  XOR2_X1   g495(.A(KEYINPUT16), .B(G8gat), .Z(new_n697));
  AND3_X1   g496(.A1(new_n692), .A2(new_n696), .A3(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n518), .B1(new_n692), .B2(new_n696), .ZN(new_n699));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT106), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n692), .A2(new_n696), .A3(new_n697), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT42), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  AND3_X1   g503(.A1(new_n700), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n701), .B1(new_n700), .B2(new_n704), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(G1325gat));
  INV_X1    g506(.A(new_n323), .ZN(new_n708));
  INV_X1    g507(.A(new_n396), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  OR3_X1    g510(.A1(new_n691), .A2(G15gat), .A3(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(G15gat), .B1(new_n691), .B2(new_n482), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(G1326gat));
  NOR2_X1   g513(.A1(new_n691), .A2(new_n393), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT107), .ZN(new_n716));
  XNOR2_X1  g515(.A(KEYINPUT43), .B(G22gat), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n716), .B(new_n717), .ZN(G1327gat));
  AOI21_X1  g517(.A(new_n632), .B1(new_n478), .B2(new_n510), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n687), .A2(new_n688), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n578), .A2(new_n720), .A3(new_n663), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n719), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n584), .A3(new_n693), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT45), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n726), .B1(new_n511), .B2(new_n631), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n631), .A2(new_n726), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n509), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n476), .A2(KEYINPUT108), .A3(new_n508), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n730), .A2(new_n482), .A3(new_n505), .A4(new_n731), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n728), .B1(new_n732), .B2(new_n478), .ZN(new_n733));
  OR2_X1    g532(.A1(new_n727), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n721), .ZN(new_n735));
  OAI21_X1  g534(.A(G29gat), .B1(new_n735), .B2(new_n475), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n725), .A2(new_n736), .ZN(G1328gat));
  NOR3_X1   g536(.A1(new_n722), .A2(G36gat), .A3(new_n471), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT46), .ZN(new_n739));
  OAI21_X1  g538(.A(G36gat), .B1(new_n735), .B2(new_n471), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n739), .A2(new_n740), .ZN(G1329gat));
  INV_X1    g540(.A(new_n482), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n734), .A2(G43gat), .A3(new_n742), .A4(new_n721), .ZN(new_n743));
  INV_X1    g542(.A(G43gat), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n722), .B2(new_n711), .ZN(new_n745));
  XNOR2_X1  g544(.A(KEYINPUT109), .B(KEYINPUT47), .ZN(new_n746));
  AND3_X1   g545(.A1(new_n743), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n746), .B1(new_n743), .B2(new_n745), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(new_n748), .ZN(G1330gat));
  NAND2_X1  g548(.A1(new_n723), .A2(new_n508), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n751));
  AOI22_X1  g550(.A1(new_n750), .A2(new_n383), .B1(new_n751), .B2(KEYINPUT48), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n751), .A2(KEYINPUT48), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n734), .A2(G50gat), .A3(new_n508), .A4(new_n721), .ZN(new_n754));
  AND3_X1   g553(.A1(new_n752), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n752), .B2(new_n754), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(G1331gat));
  INV_X1    g556(.A(new_n666), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n720), .A3(new_n663), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n759), .B1(new_n732), .B2(new_n478), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(new_n693), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n696), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n763), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n764));
  XOR2_X1   g563(.A(KEYINPUT49), .B(G64gat), .Z(new_n765));
  OAI21_X1  g564(.A(new_n764), .B1(new_n763), .B2(new_n765), .ZN(G1333gat));
  NAND2_X1  g565(.A1(new_n760), .A2(new_n742), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n711), .A2(G71gat), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n767), .A2(G71gat), .B1(new_n760), .B2(new_n768), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g569(.A1(new_n760), .A2(new_n508), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g571(.A1(new_n475), .A2(new_n664), .A3(G85gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n732), .A2(new_n478), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n578), .A2(new_n689), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n774), .A2(new_n631), .A3(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT51), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g577(.A1(new_n774), .A2(KEYINPUT51), .A3(new_n631), .A4(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n778), .A2(KEYINPUT112), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n782), .A3(new_n777), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n780), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n781), .B1(new_n780), .B2(new_n783), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n773), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n775), .A2(new_n663), .ZN(new_n787));
  XOR2_X1   g586(.A(new_n787), .B(KEYINPUT111), .Z(new_n788));
  AND2_X1   g587(.A1(new_n734), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n693), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n790), .A2(G85gat), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n786), .A2(new_n791), .ZN(G1336gat));
  NAND3_X1  g591(.A1(new_n734), .A2(new_n696), .A3(new_n788), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n793), .A2(G92gat), .ZN(new_n794));
  XNOR2_X1  g593(.A(KEYINPUT115), .B(KEYINPUT52), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n471), .A2(new_n664), .A3(G92gat), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT114), .ZN(new_n798));
  AND3_X1   g597(.A1(new_n780), .A2(new_n783), .A3(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n778), .A2(new_n779), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n793), .A2(G92gat), .B1(new_n800), .B2(new_n798), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  OAI22_X1  g601(.A1(new_n796), .A2(new_n799), .B1(new_n801), .B2(new_n802), .ZN(G1337gat));
  NOR3_X1   g602(.A1(new_n711), .A2(G99gat), .A3(new_n664), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n804), .B1(new_n784), .B2(new_n785), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n742), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(G99gat), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1338gat));
  NOR3_X1   g607(.A1(new_n393), .A2(G106gat), .A3(new_n664), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n780), .A2(new_n783), .A3(new_n809), .ZN(new_n810));
  OAI211_X1 g609(.A(new_n508), .B(new_n788), .C1(new_n727), .C2(new_n733), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT53), .B1(new_n811), .B2(G106gat), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n811), .A2(KEYINPUT116), .A3(G106gat), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT116), .B1(new_n811), .B2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(new_n809), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n816), .B1(new_n778), .B2(new_n779), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n814), .A2(new_n815), .A3(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n813), .B1(new_n818), .B2(new_n819), .ZN(G1339gat));
  NOR2_X1   g619(.A1(new_n720), .A2(G113gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n666), .A2(new_n689), .A3(new_n663), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n675), .A2(new_n676), .A3(new_n674), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n670), .B1(new_n668), .B2(new_n669), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n684), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n688), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n826), .B1(new_n626), .B2(new_n630), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT54), .ZN(new_n828));
  AND2_X1   g627(.A1(new_n657), .A2(new_n654), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n656), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n661), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n637), .B1(new_n658), .B2(new_n828), .ZN(new_n832));
  AOI21_X1  g631(.A(KEYINPUT55), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT117), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(new_n832), .A3(KEYINPUT55), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n662), .ZN(new_n837));
  INV_X1    g636(.A(new_n830), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT55), .B1(new_n838), .B2(new_n660), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n658), .A2(new_n828), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n638), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n835), .B(new_n662), .C1(new_n839), .C2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n827), .B(new_n834), .C1(new_n837), .C2(new_n843), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n664), .A2(new_n826), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n662), .B1(new_n839), .B2(new_n841), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n846), .A2(KEYINPUT117), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n833), .B1(new_n847), .B2(new_n842), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n845), .B1(new_n848), .B2(new_n689), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n844), .B1(new_n849), .B2(new_n631), .ZN(new_n850));
  INV_X1    g649(.A(new_n578), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n822), .B1(new_n850), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n852), .A2(new_n475), .ZN(new_n853));
  INV_X1    g652(.A(new_n465), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(new_n696), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT118), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n855), .A2(KEYINPUT118), .A3(new_n696), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n821), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n852), .A2(new_n508), .A3(new_n711), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n696), .A2(new_n475), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(G113gat), .B1(new_n863), .B2(new_n720), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1340gat));
  NOR2_X1   g664(.A1(new_n664), .A2(G120gat), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n858), .B2(new_n859), .ZN(new_n867));
  OAI21_X1  g666(.A(G120gat), .B1(new_n863), .B2(new_n664), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  INV_X1    g668(.A(G127gat), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n856), .A2(new_n870), .A3(new_n578), .ZN(new_n871));
  OAI21_X1  g670(.A(G127gat), .B1(new_n863), .B2(new_n851), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(G1342gat));
  INV_X1    g672(.A(G134gat), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n632), .A2(new_n696), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n853), .A2(new_n874), .A3(new_n854), .A4(new_n875), .ZN(new_n876));
  XNOR2_X1  g675(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n877), .ZN(new_n879));
  OAI21_X1  g678(.A(G134gat), .B1(new_n863), .B2(new_n632), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G1343gat));
  NOR2_X1   g680(.A1(new_n742), .A2(new_n393), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n852), .A2(new_n883), .A3(new_n475), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n884), .A2(new_n471), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n885), .A2(new_n340), .A3(new_n689), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n482), .A2(new_n862), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n720), .A2(new_n833), .A3(new_n846), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n632), .B1(new_n888), .B2(new_n845), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n578), .B1(new_n889), .B2(new_n844), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n508), .B1(new_n890), .B2(new_n822), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n887), .B1(new_n891), .B2(KEYINPUT57), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n689), .B(new_n834), .C1(new_n843), .C2(new_n837), .ZN(new_n893));
  INV_X1    g692(.A(new_n845), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n631), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n844), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n851), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n822), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n393), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n892), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(G141gat), .B1(new_n902), .B2(new_n720), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n886), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n886), .A2(new_n903), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1344gat));
  NOR2_X1   g707(.A1(new_n354), .A2(KEYINPUT59), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n909), .B1(new_n902), .B2(new_n664), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT120), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT120), .B(new_n909), .C1(new_n902), .C2(new_n664), .ZN(new_n913));
  XNOR2_X1  g712(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n665), .A2(new_n667), .A3(new_n720), .ZN(new_n915));
  OAI211_X1 g714(.A(new_n900), .B(new_n508), .C1(new_n890), .C2(new_n915), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n887), .A2(new_n664), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n916), .B(new_n917), .C1(new_n899), .C2(new_n900), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n914), .B1(new_n919), .B2(new_n342), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n912), .A2(new_n913), .A3(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n885), .A2(new_n354), .A3(new_n663), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n921), .A2(new_n922), .ZN(G1345gat));
  AOI21_X1  g722(.A(G155gat), .B1(new_n885), .B2(new_n578), .ZN(new_n924));
  INV_X1    g723(.A(new_n902), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n578), .A2(G155gat), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT122), .Z(new_n927));
  AOI21_X1  g726(.A(new_n924), .B1(new_n925), .B2(new_n927), .ZN(G1346gat));
  OAI21_X1  g727(.A(G162gat), .B1(new_n902), .B2(new_n632), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n884), .A2(new_n348), .A3(new_n875), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(G1347gat));
  NOR2_X1   g730(.A1(new_n693), .A2(new_n471), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n861), .A2(new_n932), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n933), .A2(new_n213), .A3(new_n720), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT123), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n935), .B1(new_n852), .B2(new_n693), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n897), .A2(new_n898), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n937), .A2(KEYINPUT123), .A3(new_n475), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n465), .A2(new_n471), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(new_n689), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n934), .B1(new_n942), .B2(new_n213), .ZN(G1348gat));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n214), .A3(new_n663), .ZN(new_n944));
  OAI21_X1  g743(.A(G176gat), .B1(new_n933), .B2(new_n664), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(G1349gat));
  OAI21_X1  g745(.A(G183gat), .B1(new_n933), .B2(new_n851), .ZN(new_n947));
  NAND4_X1  g746(.A1(new_n939), .A2(new_n272), .A3(new_n578), .A4(new_n940), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(KEYINPUT60), .ZN(new_n950));
  INV_X1    g749(.A(KEYINPUT60), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n947), .A2(new_n948), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n950), .A2(new_n952), .ZN(G1350gat));
  NAND3_X1  g752(.A1(new_n941), .A2(new_n273), .A3(new_n631), .ZN(new_n954));
  INV_X1    g753(.A(KEYINPUT124), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n861), .A2(new_n631), .A3(new_n932), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT61), .ZN(new_n957));
  AND4_X1   g756(.A1(new_n955), .A2(new_n956), .A3(new_n957), .A4(G190gat), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n273), .B1(KEYINPUT124), .B2(KEYINPUT61), .ZN(new_n959));
  AOI22_X1  g758(.A1(new_n956), .A2(new_n959), .B1(new_n955), .B2(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n954), .B1(new_n958), .B2(new_n960), .ZN(G1351gat));
  AND2_X1   g760(.A1(new_n482), .A2(new_n932), .ZN(new_n962));
  OAI211_X1 g761(.A(new_n916), .B(new_n962), .C1(new_n899), .C2(new_n900), .ZN(new_n963));
  OAI21_X1  g762(.A(G197gat), .B1(new_n963), .B2(new_n720), .ZN(new_n964));
  INV_X1    g763(.A(KEYINPUT125), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n883), .A2(new_n471), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n939), .A2(new_n966), .ZN(new_n967));
  INV_X1    g766(.A(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n720), .A2(G197gat), .ZN(new_n969));
  AOI21_X1  g768(.A(new_n965), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NOR4_X1   g769(.A1(new_n967), .A2(KEYINPUT125), .A3(G197gat), .A4(new_n720), .ZN(new_n971));
  OAI21_X1  g770(.A(new_n964), .B1(new_n970), .B2(new_n971), .ZN(G1352gat));
  NOR2_X1   g771(.A1(new_n664), .A2(G204gat), .ZN(new_n973));
  AOI21_X1  g772(.A(KEYINPUT123), .B1(new_n937), .B2(new_n475), .ZN(new_n974));
  AOI211_X1 g773(.A(new_n935), .B(new_n693), .C1(new_n897), .C2(new_n898), .ZN(new_n975));
  OAI211_X1 g774(.A(new_n966), .B(new_n973), .C1(new_n974), .C2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT62), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n939), .A2(new_n978), .A3(new_n966), .A4(new_n973), .ZN(new_n979));
  OAI21_X1  g778(.A(G204gat), .B1(new_n963), .B2(new_n664), .ZN(new_n980));
  NAND3_X1  g779(.A1(new_n977), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n981), .A2(KEYINPUT126), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT126), .ZN(new_n983));
  NAND4_X1  g782(.A1(new_n977), .A2(new_n979), .A3(new_n983), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n982), .A2(new_n984), .ZN(G1353gat));
  NAND3_X1  g784(.A1(new_n968), .A2(new_n327), .A3(new_n578), .ZN(new_n986));
  AND2_X1   g785(.A1(KEYINPUT127), .A2(KEYINPUT63), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n963), .A2(new_n851), .ZN(new_n988));
  OAI21_X1  g787(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n989));
  INV_X1    g788(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g789(.A(new_n987), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g790(.A(new_n987), .B(new_n990), .C1(new_n963), .C2(new_n851), .ZN(new_n992));
  INV_X1    g791(.A(new_n992), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n986), .B1(new_n991), .B2(new_n993), .ZN(G1354gat));
  OAI21_X1  g793(.A(G218gat), .B1(new_n963), .B2(new_n632), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n631), .A2(new_n328), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n995), .B1(new_n967), .B2(new_n996), .ZN(G1355gat));
endmodule


