//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 0 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:45 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n783, new_n784, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XOR2_X1   g002(.A(new_n188), .B(KEYINPUT79), .Z(new_n189));
  INV_X1    g003(.A(G469), .ZN(new_n190));
  INV_X1    g004(.A(G902), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G110), .B(G140), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT80), .ZN(new_n194));
  INV_X1    g008(.A(G227), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G953), .ZN(new_n196));
  XNOR2_X1  g010(.A(new_n194), .B(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT3), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT3), .ZN(new_n201));
  INV_X1    g015(.A(G107), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n202), .A3(G104), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n199), .A2(G107), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n200), .A2(new_n203), .A3(new_n204), .A4(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n199), .A2(G107), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n202), .A2(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(G101), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(KEYINPUT1), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  INV_X1    g026(.A(G143), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  AND4_X1   g028(.A1(new_n210), .A2(new_n212), .A3(new_n214), .A4(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(KEYINPUT1), .B1(new_n213), .B2(G146), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n216), .A2(G128), .B1(new_n212), .B2(new_n214), .ZN(new_n217));
  OAI211_X1 g031(.A(new_n206), .B(new_n209), .C1(new_n215), .C2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT10), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(KEYINPUT81), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT81), .B1(new_n218), .B2(new_n219), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT11), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n224), .B1(new_n225), .B2(G137), .ZN(new_n226));
  INV_X1    g040(.A(G137), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n227), .A2(KEYINPUT11), .A3(G134), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(G137), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n226), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G131), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n226), .A2(new_n228), .A3(new_n232), .A4(new_n229), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT65), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n230), .A2(new_n235), .A3(G131), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n200), .A2(new_n203), .A3(new_n205), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G101), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(KEYINPUT4), .A3(new_n206), .ZN(new_n241));
  AND3_X1   g055(.A1(new_n213), .A2(KEYINPUT64), .A3(G146), .ZN(new_n242));
  AOI21_X1  g056(.A(KEYINPUT64), .B1(new_n213), .B2(G146), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n212), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  AND2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NOR2_X1   g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n212), .A2(new_n214), .ZN(new_n248));
  AOI22_X1  g062(.A1(new_n244), .A2(new_n247), .B1(new_n248), .B2(new_n245), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n239), .A2(new_n250), .A3(G101), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n241), .A2(new_n249), .A3(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G128), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(new_n212), .B2(KEYINPUT1), .ZN(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n244), .A2(new_n255), .A3(KEYINPUT66), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT66), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n213), .A2(G146), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n259));
  OAI21_X1  g073(.A(new_n259), .B1(new_n211), .B2(G143), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n213), .A2(KEYINPUT64), .A3(G146), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n258), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n257), .B1(new_n262), .B2(new_n254), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n215), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n206), .A2(new_n209), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n265), .A2(new_n219), .ZN(new_n266));
  INV_X1    g080(.A(new_n266), .ZN(new_n267));
  OAI21_X1  g081(.A(new_n252), .B1(new_n264), .B2(new_n267), .ZN(new_n268));
  NOR3_X1   g082(.A1(new_n223), .A2(new_n238), .A3(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n241), .A2(new_n251), .ZN(new_n270));
  INV_X1    g084(.A(new_n215), .ZN(new_n271));
  AOI21_X1  g085(.A(KEYINPUT66), .B1(new_n244), .B2(new_n255), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n262), .A2(new_n257), .A3(new_n254), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n270), .A2(new_n249), .B1(new_n274), .B2(new_n266), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n218), .A2(new_n219), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT81), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n220), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n237), .B1(new_n275), .B2(new_n279), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n198), .B1(new_n269), .B2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n275), .A2(new_n237), .A3(new_n279), .ZN(new_n282));
  AND2_X1   g096(.A1(new_n206), .A2(new_n209), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n218), .B1(new_n274), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT12), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n285), .A3(new_n238), .ZN(new_n286));
  INV_X1    g100(.A(new_n218), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n264), .B2(new_n265), .ZN(new_n288));
  OAI21_X1  g102(.A(KEYINPUT12), .B1(new_n288), .B2(new_n237), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n282), .A2(new_n197), .A3(new_n286), .A4(new_n289), .ZN(new_n290));
  AOI21_X1  g104(.A(G902), .B1(new_n281), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n192), .B1(new_n291), .B2(new_n190), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n282), .A2(new_n286), .A3(new_n289), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n198), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n238), .B1(new_n223), .B2(new_n268), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n295), .A2(new_n282), .A3(new_n197), .ZN(new_n296));
  AND2_X1   g110(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(G469), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n189), .B1(new_n292), .B2(new_n298), .ZN(new_n299));
  NOR2_X1   g113(.A1(G475), .A2(G902), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(G113), .B(G122), .ZN(new_n302));
  XNOR2_X1  g116(.A(new_n302), .B(new_n199), .ZN(new_n303));
  INV_X1    g117(.A(G237), .ZN(new_n304));
  INV_X1    g118(.A(G953), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(G214), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(G143), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(KEYINPUT18), .A3(G131), .ZN(new_n309));
  XNOR2_X1  g123(.A(G125), .B(G140), .ZN(new_n310));
  XNOR2_X1  g124(.A(new_n310), .B(new_n211), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT18), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n307), .B1(new_n312), .B2(new_n232), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G125), .ZN(new_n315));
  NOR3_X1   g129(.A1(new_n315), .A2(KEYINPUT16), .A3(G140), .ZN(new_n316));
  INV_X1    g130(.A(G140), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G125), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n315), .A2(G140), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n318), .A2(new_n319), .A3(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT74), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n318), .A2(KEYINPUT74), .A3(KEYINPUT16), .ZN(new_n323));
  OAI211_X1 g137(.A(KEYINPUT76), .B(new_n211), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT76), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n322), .A2(new_n323), .ZN(new_n326));
  OAI21_X1  g140(.A(new_n325), .B1(new_n326), .B2(G146), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT75), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n328), .B1(new_n326), .B2(G146), .ZN(new_n329));
  NOR4_X1   g143(.A1(new_n322), .A2(KEYINPUT75), .A3(new_n211), .A4(new_n323), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n324), .B(new_n327), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n308), .A2(KEYINPUT17), .A3(G131), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n307), .B(new_n232), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n332), .B1(new_n333), .B2(KEYINPUT17), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n303), .B(new_n314), .C1(new_n331), .C2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n323), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT74), .B1(new_n310), .B2(KEYINPUT16), .ZN(new_n337));
  OAI211_X1 g151(.A(G146), .B(new_n336), .C1(new_n337), .C2(new_n316), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT86), .ZN(new_n339));
  AND3_X1   g153(.A1(new_n310), .A2(new_n339), .A3(KEYINPUT19), .ZN(new_n340));
  AOI21_X1  g154(.A(KEYINPUT19), .B1(new_n310), .B2(new_n339), .ZN(new_n341));
  OAI21_X1  g155(.A(new_n211), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n333), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n314), .ZN(new_n344));
  INV_X1    g158(.A(new_n303), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g160(.A(new_n301), .B1(new_n335), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI211_X1 g163(.A(KEYINPUT20), .B(new_n301), .C1(new_n335), .C2(new_n346), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n314), .B1(new_n331), .B2(new_n334), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n351), .A2(new_n345), .ZN(new_n352));
  AOI21_X1  g166(.A(G902), .B1(new_n352), .B2(new_n335), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT87), .B(G475), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n349), .A2(new_n350), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G217), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n187), .A2(new_n357), .A3(G953), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  INV_X1    g173(.A(G116), .ZN(new_n360));
  OR2_X1    g174(.A1(new_n360), .A2(G122), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(G122), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G107), .ZN(new_n364));
  NAND3_X1  g178(.A1(new_n361), .A2(new_n362), .A3(new_n202), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G128), .B(G143), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(new_n225), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n367), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT88), .B(KEYINPUT13), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n372), .A2(G128), .A3(new_n213), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(G134), .A3(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT89), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n374), .A2(new_n375), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n369), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OR2_X1    g193(.A1(new_n367), .A2(new_n225), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n368), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT90), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n365), .B(KEYINPUT91), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n380), .A2(KEYINPUT90), .A3(new_n368), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n361), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n388));
  OAI21_X1  g202(.A(G107), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n383), .A2(new_n384), .A3(new_n385), .A4(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n359), .B1(new_n379), .B2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(new_n378), .ZN(new_n393));
  OAI211_X1 g207(.A(new_n368), .B(new_n366), .C1(new_n393), .C2(new_n376), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n390), .A3(new_n358), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n392), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n191), .ZN(new_n397));
  INV_X1    g211(.A(G478), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n398), .A2(KEYINPUT15), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(new_n399), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n191), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n305), .A2(G952), .ZN(new_n404));
  INV_X1    g218(.A(G234), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n304), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  AOI211_X1 g221(.A(new_n191), .B(new_n305), .C1(G234), .C2(G237), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT21), .B(G898), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n407), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n356), .A2(new_n403), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(G214), .B1(G237), .B2(G902), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(G110), .B(G122), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n414), .B(KEYINPUT82), .ZN(new_n415));
  XNOR2_X1  g229(.A(KEYINPUT2), .B(G113), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G116), .B(G119), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(G119), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(G116), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n360), .A2(G119), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n419), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n241), .A2(new_n425), .A3(new_n251), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n418), .A2(KEYINPUT5), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n427), .B(G113), .C1(KEYINPUT5), .C2(new_n421), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n283), .A3(new_n419), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n415), .B1(new_n426), .B2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(KEYINPUT6), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n426), .A2(new_n429), .A3(new_n414), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT83), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g249(.A1(new_n426), .A2(new_n429), .A3(KEYINPUT83), .A4(new_n414), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n432), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n431), .B1(new_n437), .B2(new_n430), .ZN(new_n438));
  AOI211_X1 g252(.A(G125), .B(new_n215), .C1(new_n256), .C2(new_n263), .ZN(new_n439));
  NOR2_X1   g253(.A1(new_n249), .A2(new_n315), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n305), .A2(G224), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n443), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n414), .B(KEYINPUT8), .ZN(new_n445));
  INV_X1    g259(.A(new_n427), .ZN(new_n446));
  OAI21_X1  g260(.A(G113), .B1(new_n421), .B2(KEYINPUT5), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n419), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n265), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n447), .A2(KEYINPUT84), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT84), .ZN(new_n451));
  OAI211_X1 g265(.A(new_n451), .B(G113), .C1(new_n421), .C2(KEYINPUT5), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n427), .A3(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n453), .A2(new_n283), .A3(new_n419), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT85), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n449), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n265), .B1(new_n418), .B2(new_n417), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT85), .B1(new_n457), .B2(new_n453), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n445), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n460), .B1(new_n439), .B2(new_n440), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n264), .A2(new_n315), .ZN(new_n462));
  INV_X1    g276(.A(new_n440), .ZN(new_n463));
  NAND4_X1  g277(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT7), .A4(new_n442), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n459), .A2(new_n461), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n435), .A2(new_n436), .ZN(new_n466));
  AOI21_X1  g280(.A(G902), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n444), .A2(new_n467), .ZN(new_n468));
  OAI21_X1  g282(.A(G210), .B1(G237), .B2(G902), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n444), .A2(new_n467), .A3(new_n469), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n413), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NAND3_X1  g287(.A1(new_n299), .A2(new_n411), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT92), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT68), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n234), .A2(new_n249), .A3(new_n236), .ZN(new_n477));
  INV_X1    g291(.A(new_n229), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n225), .A2(G137), .ZN(new_n479));
  OAI21_X1  g293(.A(G131), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n233), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n477), .B(KEYINPUT30), .C1(new_n264), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n425), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n484));
  INV_X1    g298(.A(new_n481), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n274), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(KEYINPUT67), .B1(new_n264), .B2(new_n481), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n486), .A2(new_n487), .A3(new_n477), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT30), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n483), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n425), .ZN(new_n491));
  OAI211_X1 g305(.A(new_n477), .B(new_n491), .C1(new_n264), .C2(new_n481), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n304), .A2(new_n305), .A3(G210), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(KEYINPUT27), .ZN(new_n494));
  XNOR2_X1  g308(.A(KEYINPUT26), .B(G101), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n494), .B(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n492), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n476), .B1(new_n490), .B2(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n497), .ZN(new_n499));
  INV_X1    g313(.A(new_n477), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n274), .A2(new_n485), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(KEYINPUT67), .ZN(new_n502));
  AOI21_X1  g316(.A(KEYINPUT30), .B1(new_n502), .B2(new_n486), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT68), .B(new_n499), .C1(new_n503), .C2(new_n483), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n504), .A3(KEYINPUT31), .ZN(new_n505));
  INV_X1    g319(.A(new_n492), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n506), .B1(new_n488), .B2(new_n425), .ZN(new_n507));
  XOR2_X1   g321(.A(KEYINPUT70), .B(KEYINPUT28), .Z(new_n508));
  OAI22_X1  g322(.A1(new_n507), .A2(new_n508), .B1(KEYINPUT28), .B2(new_n506), .ZN(new_n509));
  INV_X1    g323(.A(new_n496), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NOR4_X1   g325(.A1(new_n490), .A2(KEYINPUT69), .A3(KEYINPUT31), .A4(new_n497), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n488), .A2(new_n489), .ZN(new_n514));
  INV_X1    g328(.A(new_n483), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n497), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT31), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n505), .B(new_n511), .C1(new_n512), .C2(new_n518), .ZN(new_n519));
  NOR2_X1   g333(.A1(G472), .A2(G902), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT32), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n519), .A2(KEYINPUT32), .A3(new_n520), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n510), .B1(new_n490), .B2(new_n506), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT29), .ZN(new_n526));
  OAI211_X1 g340(.A(new_n525), .B(new_n526), .C1(new_n509), .C2(new_n510), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n506), .A2(KEYINPUT28), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n501), .A2(new_n477), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n425), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(new_n492), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n528), .B1(new_n531), .B2(KEYINPUT28), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n510), .A2(new_n526), .ZN(new_n533));
  AOI21_X1  g347(.A(G902), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n527), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(G472), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n523), .A2(new_n524), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n253), .A2(G119), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n420), .A2(G128), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT72), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n540), .B1(new_n538), .B2(new_n539), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT24), .B(G110), .ZN(new_n544));
  OR2_X1    g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT23), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n546), .B1(new_n420), .B2(G128), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT73), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n420), .B2(G128), .ZN(new_n549));
  NOR2_X1   g363(.A1(KEYINPUT73), .A2(KEYINPUT23), .ZN(new_n550));
  OAI22_X1  g364(.A1(new_n547), .A2(new_n549), .B1(new_n538), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(G110), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n336), .B1(new_n337), .B2(new_n316), .ZN(new_n554));
  AOI21_X1  g368(.A(KEYINPUT76), .B1(new_n554), .B2(new_n211), .ZN(new_n555));
  INV_X1    g369(.A(new_n324), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n326), .A2(new_n328), .A3(G146), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n338), .A2(KEYINPUT75), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n553), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n310), .A2(new_n211), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n338), .A2(new_n562), .ZN(new_n563));
  OR2_X1    g377(.A1(new_n551), .A2(G110), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n544), .B1(new_n541), .B2(new_n542), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT77), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(KEYINPUT77), .A3(new_n565), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n563), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g384(.A(KEYINPUT78), .B1(new_n561), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n553), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n331), .A2(new_n572), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT78), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n568), .A2(new_n569), .ZN(new_n575));
  INV_X1    g389(.A(new_n563), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n573), .A2(new_n574), .A3(new_n577), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT22), .B(G137), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n305), .A2(G221), .A3(G234), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n579), .B(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n571), .A2(new_n578), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n573), .A2(new_n577), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(KEYINPUT78), .A3(new_n581), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n357), .B1(G234), .B2(new_n191), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(G902), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n586), .A2(new_n191), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT25), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n586), .A2(KEYINPUT25), .A3(new_n191), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n588), .B(KEYINPUT71), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n591), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT92), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n299), .A2(new_n411), .A3(new_n473), .A4(new_n599), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n475), .A2(new_n537), .A3(new_n598), .A4(new_n600), .ZN(new_n601));
  XOR2_X1   g415(.A(KEYINPUT93), .B(G101), .Z(new_n602));
  XNOR2_X1  g416(.A(new_n601), .B(new_n602), .ZN(G3));
  AOI21_X1  g417(.A(KEYINPUT25), .B1(new_n586), .B2(new_n191), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n593), .B(G902), .C1(new_n583), .C2(new_n585), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n597), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n587), .B2(new_n590), .ZN(new_n607));
  INV_X1    g421(.A(new_n299), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(KEYINPUT94), .A2(G472), .ZN(new_n610));
  AND3_X1   g424(.A1(new_n519), .A2(new_n191), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n610), .B1(new_n519), .B2(new_n191), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n609), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n410), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n394), .A2(new_n390), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT95), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(KEYINPUT33), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n618), .A2(new_n396), .ZN(new_n619));
  NAND4_X1  g433(.A1(new_n617), .A2(KEYINPUT33), .A3(new_n395), .A4(new_n392), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n398), .A2(G902), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT96), .B(G478), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n397), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n622), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n356), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n614), .A2(new_n473), .A3(new_n615), .A4(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(G6));
  INV_X1    g444(.A(KEYINPUT97), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n401), .B1(new_n396), .B2(new_n191), .ZN(new_n632));
  AOI211_X1 g446(.A(G902), .B(new_n399), .C1(new_n392), .C2(new_n395), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n356), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AND3_X1   g450(.A1(new_n444), .A2(new_n467), .A3(new_n469), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n469), .B1(new_n444), .B2(new_n467), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n412), .B(new_n615), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n631), .B1(new_n636), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n473), .A2(KEYINPUT97), .A3(new_n615), .A4(new_n635), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n614), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT98), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT35), .B(G107), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G9));
  INV_X1    g459(.A(KEYINPUT36), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n581), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT100), .ZN(new_n648));
  XOR2_X1   g462(.A(new_n648), .B(KEYINPUT99), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n584), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n589), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n606), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n475), .A2(new_n613), .A3(new_n600), .A4(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  AND3_X1   g469(.A1(new_n652), .A2(new_n473), .A3(new_n299), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n537), .ZN(new_n657));
  INV_X1    g471(.A(G900), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n407), .B1(new_n408), .B2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n635), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n253), .ZN(G30));
  XOR2_X1   g477(.A(new_n659), .B(KEYINPUT39), .Z(new_n664));
  NAND2_X1  g478(.A1(new_n299), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g479(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n665), .A2(KEYINPUT40), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n471), .A2(new_n472), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT38), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n413), .B1(new_n400), .B2(new_n402), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n356), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n652), .A2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n666), .A2(new_n667), .A3(new_n669), .A4(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n524), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT32), .B1(new_n519), .B2(new_n520), .ZN(new_n675));
  INV_X1    g489(.A(G472), .ZN(new_n676));
  AND2_X1   g490(.A1(new_n498), .A2(new_n504), .ZN(new_n677));
  INV_X1    g491(.A(new_n531), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n677), .B1(new_n496), .B2(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n676), .B1(new_n679), .B2(new_n191), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n673), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT101), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT102), .B(G143), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G45));
  NOR2_X1   g499(.A1(new_n626), .A2(new_n659), .ZN(new_n686));
  INV_X1    g500(.A(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n657), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(new_n211), .ZN(G48));
  AND4_X1   g503(.A1(new_n282), .A2(new_n197), .A3(new_n286), .A4(new_n289), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n197), .B1(new_n295), .B2(new_n282), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n191), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(G469), .ZN(new_n693));
  OAI211_X1 g507(.A(new_n190), .B(new_n191), .C1(new_n690), .C2(new_n691), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n693), .A2(new_n694), .A3(new_n188), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n639), .A2(new_n626), .A3(new_n695), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n524), .A2(new_n536), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n696), .B(new_n598), .C1(new_n675), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(KEYINPUT41), .B(G113), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G15));
  INV_X1    g514(.A(new_n695), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n598), .B(new_n701), .C1(new_n697), .C2(new_n675), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n640), .A2(new_n641), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  XOR2_X1   g518(.A(KEYINPUT103), .B(G116), .Z(new_n705));
  XNOR2_X1  g519(.A(new_n704), .B(new_n705), .ZN(G18));
  XNOR2_X1  g520(.A(new_n347), .B(new_n348), .ZN(new_n707));
  OR2_X1    g521(.A1(new_n353), .A2(new_n355), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n707), .A2(new_n708), .A3(new_n615), .A4(new_n634), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n709), .B1(new_n606), .B2(new_n651), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n637), .A2(new_n638), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n711), .A2(new_n695), .A3(new_n413), .ZN(new_n712));
  OAI211_X1 g526(.A(new_n710), .B(new_n712), .C1(new_n697), .C2(new_n675), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G119), .ZN(G21));
  OAI21_X1  g528(.A(KEYINPUT105), .B1(new_n711), .B2(new_n671), .ZN(new_n715));
  INV_X1    g529(.A(KEYINPUT105), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n668), .A2(new_n716), .A3(new_n356), .A4(new_n670), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n519), .A2(new_n191), .ZN(new_n719));
  OAI221_X1 g533(.A(new_n505), .B1(new_n496), .B2(new_n532), .C1(new_n512), .C2(new_n518), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n520), .B(KEYINPUT104), .ZN(new_n721));
  AOI22_X1  g535(.A1(new_n719), .A2(G472), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n695), .A2(new_n410), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n718), .A2(new_n598), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  NAND2_X1  g539(.A1(new_n712), .A2(new_n686), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n719), .A2(G472), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT106), .ZN(new_n729));
  OAI22_X1  g543(.A1(new_n518), .A2(new_n512), .B1(new_n496), .B2(new_n532), .ZN(new_n730));
  INV_X1    g544(.A(new_n505), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n721), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n728), .A2(new_n652), .A3(new_n729), .A4(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n729), .B1(new_n722), .B2(new_n652), .ZN(new_n735));
  OAI21_X1  g549(.A(new_n727), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n736), .A2(KEYINPUT107), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n517), .B(new_n499), .C1(new_n503), .C2(new_n483), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(KEYINPUT69), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n516), .A2(new_n513), .A3(new_n517), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n739), .A2(new_n740), .B1(new_n510), .B2(new_n509), .ZN(new_n741));
  AOI21_X1  g555(.A(G902), .B1(new_n741), .B2(new_n505), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n732), .B1(new_n742), .B2(new_n676), .ZN(new_n743));
  INV_X1    g557(.A(new_n651), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n744), .B1(new_n596), .B2(new_n597), .ZN(new_n745));
  OAI21_X1  g559(.A(KEYINPUT106), .B1(new_n743), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n746), .A2(new_n733), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT107), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n747), .A2(new_n748), .A3(new_n727), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n737), .A2(new_n749), .ZN(new_n750));
  XNOR2_X1  g564(.A(new_n750), .B(G125), .ZN(G27));
  NAND2_X1  g565(.A1(new_n523), .A2(KEYINPUT109), .ZN(new_n752));
  AND2_X1   g566(.A1(new_n524), .A2(new_n536), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT109), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n675), .A2(new_n754), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n752), .A2(new_n753), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(new_n188), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT108), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n293), .B2(new_n198), .ZN(new_n759));
  INV_X1    g573(.A(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n293), .A2(new_n758), .A3(new_n198), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n760), .A2(G469), .A3(new_n296), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n757), .B1(new_n762), .B2(new_n292), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n471), .A2(new_n412), .A3(new_n472), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  AND4_X1   g579(.A1(KEYINPUT42), .A2(new_n686), .A3(new_n763), .A4(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n756), .A2(new_n598), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(KEYINPUT110), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT110), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n756), .A2(new_n769), .A3(new_n598), .A4(new_n766), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT42), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n761), .A2(new_n296), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n772), .A2(new_n190), .A3(new_n759), .ZN(new_n773));
  INV_X1    g587(.A(new_n192), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n694), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n188), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n764), .ZN(new_n777));
  OAI211_X1 g591(.A(new_n777), .B(new_n598), .C1(new_n697), .C2(new_n675), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n686), .ZN(new_n780));
  AOI22_X1  g594(.A1(new_n768), .A2(new_n770), .B1(new_n771), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g595(.A(new_n781), .B(new_n232), .ZN(G33));
  INV_X1    g596(.A(new_n661), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n779), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G134), .ZN(G36));
  NAND4_X1  g599(.A1(new_n760), .A2(KEYINPUT45), .A3(new_n296), .A4(new_n761), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n786), .B(G469), .C1(KEYINPUT45), .C2(new_n297), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n787), .A2(new_n774), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(KEYINPUT46), .ZN(new_n789));
  OAI21_X1  g603(.A(new_n694), .B1(new_n788), .B2(KEYINPUT46), .ZN(new_n790));
  OAI211_X1 g604(.A(new_n188), .B(new_n664), .C1(new_n789), .C2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n764), .B(KEYINPUT112), .ZN(new_n793));
  AND2_X1   g607(.A1(new_n622), .A2(new_n624), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n356), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT43), .ZN(new_n798));
  OAI22_X1  g612(.A1(new_n794), .A2(new_n356), .B1(KEYINPUT111), .B2(new_n798), .ZN(new_n799));
  AOI21_X1  g613(.A(new_n745), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(new_n613), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n802), .A2(KEYINPUT44), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(KEYINPUT44), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n792), .B(new_n793), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G137), .ZN(G39));
  OAI21_X1  g620(.A(new_n188), .B1(new_n789), .B2(new_n790), .ZN(new_n807));
  XOR2_X1   g621(.A(KEYINPUT113), .B(KEYINPUT47), .Z(new_n808));
  OR2_X1    g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n807), .B1(KEYINPUT113), .B2(KEYINPUT47), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n537), .A2(new_n598), .A3(new_n687), .A4(new_n764), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G140), .ZN(G42));
  NAND2_X1  g627(.A1(new_n693), .A2(new_n694), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(KEYINPUT49), .ZN(new_n815));
  INV_X1    g629(.A(new_n189), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n795), .A2(new_n412), .A3(new_n816), .ZN(new_n817));
  NOR3_X1   g631(.A1(new_n815), .A2(new_n817), .A3(new_n607), .ZN(new_n818));
  INV_X1    g632(.A(new_n669), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n681), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n777), .A2(new_n686), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(new_n746), .B2(new_n733), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n356), .A2(new_n403), .A3(new_n659), .ZN(new_n823));
  AND2_X1   g637(.A1(new_n299), .A2(new_n823), .ZN(new_n824));
  AOI21_X1  g638(.A(new_n764), .B1(new_n606), .B2(new_n651), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n824), .B(new_n825), .C1(new_n697), .C2(new_n675), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n778), .B2(new_n661), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n822), .A2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n724), .A2(new_n698), .A3(new_n713), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n829), .A2(new_n704), .ZN(new_n830));
  AOI21_X1  g644(.A(new_n639), .B1(new_n636), .B2(new_n626), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n609), .A2(new_n613), .A3(new_n831), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n601), .A2(new_n653), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n828), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n834), .A2(new_n781), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n656), .B(new_n537), .C1(new_n783), .C2(new_n686), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n718), .A2(new_n745), .A3(new_n660), .A4(new_n763), .ZN(new_n837));
  OR2_X1    g651(.A1(new_n837), .A2(new_n681), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n748), .B1(new_n747), .B2(new_n727), .ZN(new_n839));
  AOI211_X1 g653(.A(KEYINPUT107), .B(new_n726), .C1(new_n746), .C2(new_n733), .ZN(new_n840));
  OAI211_X1 g654(.A(new_n836), .B(new_n838), .C1(new_n839), .C2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n841), .A2(KEYINPUT52), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT52), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n750), .A2(new_n843), .A3(new_n836), .A4(new_n838), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n835), .A2(new_n842), .A3(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT54), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  OR3_X1    g663(.A1(new_n829), .A2(KEYINPUT114), .A3(new_n704), .ZN(new_n850));
  AND4_X1   g664(.A1(KEYINPUT53), .A2(new_n601), .A3(new_n653), .A4(new_n832), .ZN(new_n851));
  OAI21_X1  g665(.A(KEYINPUT114), .B1(new_n829), .B2(new_n704), .ZN(new_n852));
  AND4_X1   g666(.A1(new_n828), .A2(new_n850), .A3(new_n851), .A4(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n781), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n853), .A2(new_n854), .A3(new_n842), .A4(new_n844), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n848), .B1(KEYINPUT54), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n764), .A2(new_n695), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n681), .A2(new_n598), .A3(new_n407), .A4(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n797), .A2(new_n799), .ZN(new_n860));
  AOI21_X1  g674(.A(KEYINPUT115), .B1(new_n860), .B2(new_n407), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n860), .A2(KEYINPUT115), .A3(new_n407), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n743), .A2(new_n607), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n712), .ZN(new_n867));
  OAI221_X1 g681(.A(new_n404), .B1(new_n626), .B2(new_n859), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n864), .A2(new_n858), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(new_n598), .A3(new_n756), .ZN(new_n871));
  INV_X1    g685(.A(new_n871), .ZN(new_n872));
  OR2_X1    g686(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n872), .A2(KEYINPUT48), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n868), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g689(.A(new_n866), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n669), .A2(new_n412), .A3(new_n695), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n876), .A2(KEYINPUT50), .A3(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT50), .ZN(new_n879));
  INV_X1    g693(.A(new_n877), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n866), .B2(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n878), .A2(new_n881), .B1(new_n747), .B2(new_n870), .ZN(new_n882));
  AND2_X1   g696(.A1(new_n809), .A2(new_n810), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n814), .A2(new_n816), .ZN(new_n884));
  OAI211_X1 g698(.A(new_n876), .B(new_n793), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n859), .A2(new_n356), .A3(new_n625), .ZN(new_n886));
  XOR2_X1   g700(.A(new_n886), .B(KEYINPUT116), .Z(new_n887));
  NAND3_X1  g701(.A1(new_n882), .A2(new_n885), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT51), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n875), .A2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n888), .A2(new_n889), .ZN(new_n892));
  NOR3_X1   g706(.A1(new_n857), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(G952), .A2(G953), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n820), .B1(new_n893), .B2(new_n894), .ZN(G75));
  NAND3_X1  g709(.A1(new_n856), .A2(G210), .A3(G902), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n438), .B(new_n443), .ZN(new_n898));
  XNOR2_X1  g712(.A(KEYINPUT117), .B(KEYINPUT55), .ZN(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n896), .A2(new_n897), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n191), .B1(new_n849), .B2(new_n855), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT56), .B1(new_n905), .B2(G210), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(KEYINPUT119), .A3(new_n901), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n909), .B1(new_n906), .B2(new_n901), .ZN(new_n910));
  INV_X1    g724(.A(G210), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n911), .B(new_n191), .C1(new_n849), .C2(new_n855), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT118), .B(new_n900), .C1(new_n912), .C2(KEYINPUT56), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n910), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n305), .A2(G952), .ZN(new_n915));
  INV_X1    g729(.A(new_n915), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n908), .A2(new_n914), .A3(new_n916), .ZN(G51));
  XNOR2_X1  g731(.A(new_n856), .B(KEYINPUT54), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n192), .B(KEYINPUT57), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n920), .B1(new_n691), .B2(new_n690), .ZN(new_n921));
  INV_X1    g735(.A(new_n905), .ZN(new_n922));
  OR2_X1    g736(.A1(new_n922), .A2(new_n787), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n915), .B1(new_n921), .B2(new_n923), .ZN(G54));
  AND3_X1   g738(.A1(new_n905), .A2(KEYINPUT58), .A3(G475), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n335), .A2(new_n346), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n916), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n926), .B2(new_n925), .ZN(G60));
  AND2_X1   g742(.A1(new_n619), .A2(new_n620), .ZN(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT59), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n918), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n916), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n929), .B1(new_n857), .B2(new_n931), .ZN(new_n934));
  NOR2_X1   g748(.A1(new_n933), .A2(new_n934), .ZN(G63));
  XNOR2_X1  g749(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n357), .A2(new_n191), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n936), .B(new_n937), .Z(new_n938));
  AOI21_X1  g752(.A(new_n938), .B1(new_n849), .B2(new_n855), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(new_n586), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(new_n650), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n916), .A3(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(KEYINPUT61), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n942), .B(new_n943), .ZN(G66));
  INV_X1    g758(.A(G224), .ZN(new_n945));
  OAI21_X1  g759(.A(G953), .B1(new_n409), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n830), .A2(new_n833), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n946), .B1(new_n948), .B2(G953), .ZN(new_n949));
  INV_X1    g763(.A(new_n438), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(G898), .B2(new_n305), .ZN(new_n951));
  XOR2_X1   g765(.A(new_n951), .B(KEYINPUT121), .Z(new_n952));
  XNOR2_X1  g766(.A(new_n949), .B(new_n952), .ZN(G69));
  INV_X1    g767(.A(KEYINPUT123), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n764), .B1(new_n636), .B2(new_n626), .ZN(new_n955));
  INV_X1    g769(.A(new_n665), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n537), .A2(new_n955), .A3(new_n598), .A4(new_n956), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n812), .A2(new_n805), .A3(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n836), .B1(new_n839), .B2(new_n840), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(KEYINPUT122), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT122), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n750), .A2(new_n961), .A3(new_n836), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n683), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT62), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n958), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  AOI211_X1 g779(.A(KEYINPUT62), .B(new_n683), .C1(new_n960), .C2(new_n962), .ZN(new_n966));
  OAI21_X1  g780(.A(new_n954), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n960), .A2(new_n962), .ZN(new_n968));
  OAI21_X1  g782(.A(KEYINPUT62), .B1(new_n968), .B2(new_n683), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n964), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n969), .A2(KEYINPUT123), .A3(new_n970), .A4(new_n958), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n967), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n514), .A2(new_n482), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n340), .A2(new_n341), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n973), .B(new_n974), .Z(new_n975));
  NAND3_X1  g789(.A1(new_n972), .A2(new_n305), .A3(new_n975), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n792), .A2(new_n598), .A3(new_n718), .A4(new_n756), .ZN(new_n977));
  NAND4_X1  g791(.A1(new_n812), .A2(new_n784), .A3(new_n805), .A4(new_n977), .ZN(new_n978));
  OR3_X1    g792(.A1(new_n968), .A2(new_n978), .A3(new_n781), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(new_n305), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n975), .B1(new_n195), .B2(G953), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n658), .B1(new_n975), .B2(new_n195), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n976), .B(new_n982), .C1(new_n305), .C2(new_n983), .ZN(G72));
  NAND2_X1  g798(.A1(G472), .A2(G902), .ZN(new_n985));
  XOR2_X1   g799(.A(new_n985), .B(KEYINPUT63), .Z(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n979), .B2(new_n947), .ZN(new_n987));
  NOR2_X1   g801(.A1(new_n490), .A2(new_n506), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n988), .B(KEYINPUT125), .Z(new_n989));
  NOR2_X1   g803(.A1(new_n989), .A2(new_n496), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT126), .Z(new_n991));
  NAND2_X1  g805(.A1(new_n987), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n677), .A2(new_n525), .ZN(new_n993));
  NAND3_X1  g807(.A1(new_n847), .A2(new_n986), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n992), .A2(new_n916), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n989), .A2(new_n496), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n967), .A2(new_n971), .A3(new_n948), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n986), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT124), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n997), .A2(KEYINPUT124), .A3(new_n986), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n995), .B1(new_n1000), .B2(new_n1001), .ZN(G57));
endmodule


