//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 0 1 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 0 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:03 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n445, new_n450, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n459, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT64), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g021(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g022(.A(KEYINPUT66), .B(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g026(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g028(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n454), .B(KEYINPUT2), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NAND4_X1  g031(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n457));
  XOR2_X1   g032(.A(new_n457), .B(KEYINPUT67), .Z(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g034(.A1(new_n456), .A2(new_n459), .ZN(G325));
  INV_X1    g035(.A(G325), .ZN(G261));
  AOI22_X1  g036(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n459), .ZN(G319));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(G113), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(KEYINPUT68), .ZN(new_n469));
  XNOR2_X1  g044(.A(new_n468), .B(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n467), .B2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n472), .B1(new_n463), .B2(new_n464), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n472), .A2(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n474), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n465), .A2(KEYINPUT69), .ZN(new_n479));
  OR2_X1    g054(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n480));
  NAND2_X1  g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n480), .A2(KEYINPUT69), .A3(new_n481), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n472), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n479), .B2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OR2_X1    g063(.A1(G100), .A2(G2105), .ZN(new_n489));
  OAI211_X1 g064(.A(new_n489), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  NOR2_X1   g067(.A1(KEYINPUT70), .A2(KEYINPUT4), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  OAI21_X1  g070(.A(G138), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n493), .B1(new_n473), .B2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(G126), .A2(G2105), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n498), .B1(new_n480), .B2(new_n481), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n472), .A2(G114), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  NOR2_X1   g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n480), .A2(new_n481), .ZN(new_n504));
  INV_X1    g079(.A(G138), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n505), .B1(KEYINPUT70), .B2(KEYINPUT4), .ZN(new_n506));
  INV_X1    g081(.A(new_n493), .ZN(new_n507));
  NAND4_X1  g082(.A1(new_n504), .A2(new_n506), .A3(new_n472), .A4(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n497), .A2(new_n503), .A3(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(G164));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n511), .B1(new_n512), .B2(KEYINPUT72), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n514));
  NAND4_X1  g089(.A1(new_n514), .A2(KEYINPUT71), .A3(KEYINPUT5), .A4(G543), .ZN(new_n515));
  OR2_X1    g090(.A1(KEYINPUT71), .A2(G543), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n513), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  INV_X1    g095(.A(G50), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n518), .A2(G543), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g098(.A(G651), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n517), .A2(G62), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n526), .B(KEYINPUT73), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G166));
  AND2_X1   g104(.A1(new_n518), .A2(G543), .ZN(new_n530));
  NAND3_X1  g105(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n532));
  OR2_X1    g107(.A1(new_n531), .A2(KEYINPUT7), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n530), .A2(G51), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n535));
  AND2_X1   g110(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n519), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G89), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  AOI22_X1  g115(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n524), .ZN(new_n542));
  INV_X1    g117(.A(G90), .ZN(new_n543));
  INV_X1    g118(.A(G52), .ZN(new_n544));
  OAI22_X1  g119(.A1(new_n519), .A2(new_n543), .B1(new_n544), .B2(new_n522), .ZN(new_n545));
  OR3_X1    g120(.A1(new_n542), .A2(new_n545), .A3(KEYINPUT74), .ZN(new_n546));
  OAI21_X1  g121(.A(KEYINPUT74), .B1(new_n542), .B2(new_n545), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(G171));
  INV_X1    g123(.A(G81), .ZN(new_n549));
  INV_X1    g124(.A(G43), .ZN(new_n550));
  OAI22_X1  g125(.A1(new_n519), .A2(new_n549), .B1(new_n550), .B2(new_n522), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT75), .ZN(new_n552));
  AOI22_X1  g127(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n553), .A2(new_n524), .ZN(new_n554));
  AND2_X1   g129(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT76), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n557), .A2(new_n561), .ZN(G188));
  INV_X1    g137(.A(G53), .ZN(new_n563));
  OR3_X1    g138(.A1(new_n522), .A2(KEYINPUT9), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g139(.A(KEYINPUT9), .B1(new_n522), .B2(new_n563), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(KEYINPUT77), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT77), .ZN(new_n568));
  NAND3_X1  g143(.A1(new_n564), .A2(new_n568), .A3(new_n565), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n517), .A2(G65), .ZN(new_n571));
  INV_X1    g146(.A(G78), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n572), .B2(new_n512), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(G91), .B2(new_n537), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G166), .ZN(G303));
  INV_X1    g152(.A(G87), .ZN(new_n578));
  INV_X1    g153(.A(G49), .ZN(new_n579));
  OAI22_X1  g154(.A1(new_n519), .A2(new_n578), .B1(new_n579), .B2(new_n522), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n582));
  INV_X1    g157(.A(KEYINPUT78), .ZN(new_n583));
  AND2_X1   g158(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g159(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(G288));
  NAND3_X1  g161(.A1(new_n517), .A2(G86), .A3(new_n518), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n518), .A2(G48), .A3(G543), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n590), .B1(new_n517), .B2(G61), .ZN(new_n591));
  OAI211_X1 g166(.A(new_n587), .B(new_n588), .C1(new_n591), .C2(new_n524), .ZN(G305));
  XNOR2_X1  g167(.A(KEYINPUT79), .B(G85), .ZN(new_n593));
  AOI22_X1  g168(.A1(new_n537), .A2(new_n593), .B1(G47), .B2(new_n530), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n524), .B2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(new_n537), .A2(G92), .ZN(new_n597));
  XOR2_X1   g172(.A(new_n597), .B(KEYINPUT10), .Z(new_n598));
  AOI22_X1  g173(.A1(new_n517), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n599));
  NOR2_X1   g174(.A1(new_n599), .A2(new_n524), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n600), .B1(G54), .B2(new_n530), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  MUX2_X1   g178(.A(G301), .B(new_n602), .S(new_n603), .Z(G284));
  MUX2_X1   g179(.A(G301), .B(new_n602), .S(new_n603), .Z(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  INV_X1    g181(.A(G299), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G280));
  XOR2_X1   g183(.A(G280), .B(KEYINPUT80), .Z(G297));
  NOR2_X1   g184(.A1(new_n602), .A2(G559), .ZN(new_n610));
  AND2_X1   g185(.A1(new_n598), .A2(new_n601), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(G860), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT81), .ZN(G148));
  NAND2_X1  g188(.A1(new_n552), .A2(new_n554), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(new_n603), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(new_n610), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n504), .A2(new_n475), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT83), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT82), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT13), .Z(new_n622));
  INV_X1    g197(.A(G2100), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n484), .A2(G135), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n487), .A2(G123), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n472), .A2(G111), .ZN(new_n628));
  OAI21_X1  g203(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n629));
  OAI211_X1 g204(.A(new_n626), .B(new_n627), .C1(new_n628), .C2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  NAND3_X1  g206(.A1(new_n624), .A2(new_n625), .A3(new_n631), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2067), .B(G2678), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT84), .ZN(new_n649));
  XOR2_X1   g224(.A(G2072), .B(G2078), .Z(new_n650));
  XNOR2_X1  g225(.A(G2084), .B(G2090), .ZN(new_n651));
  NOR3_X1   g226(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT18), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n650), .A2(KEYINPUT85), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(KEYINPUT85), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT86), .B(KEYINPUT17), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n650), .B(new_n657), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n656), .B(new_n651), .C1(new_n658), .C2(new_n649), .ZN(new_n659));
  INV_X1    g234(.A(new_n651), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n658), .A2(new_n649), .A3(new_n660), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n653), .A2(new_n659), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(KEYINPUT87), .B(KEYINPUT19), .Z(new_n665));
  XNOR2_X1  g240(.A(G1971), .B(G1976), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1956), .B(G2474), .ZN(new_n668));
  XNOR2_X1  g243(.A(G1961), .B(G1966), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT20), .ZN(new_n672));
  NAND3_X1  g247(.A1(new_n667), .A2(new_n668), .A3(new_n669), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(new_n669), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n672), .B(new_n673), .C1(new_n667), .C2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G1991), .B(G1996), .Z(new_n678));
  INV_X1    g253(.A(new_n678), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n679), .ZN(new_n682));
  AND3_X1   g257(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g258(.A(new_n681), .B1(new_n680), .B2(new_n682), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(G229));
  INV_X1    g260(.A(G16), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n686), .A2(G23), .ZN(new_n687));
  INV_X1    g262(.A(G288), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(new_n686), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT33), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n686), .A2(G22), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G166), .B2(new_n686), .ZN(new_n693));
  INV_X1    g268(.A(G1971), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  NOR2_X1   g270(.A1(G6), .A2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G305), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  AND3_X1   g275(.A1(new_n691), .A2(new_n695), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT34), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n701), .A2(new_n702), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n484), .A2(G131), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT88), .Z(new_n706));
  OAI21_X1  g281(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n707));
  INV_X1    g282(.A(G107), .ZN(new_n708));
  AOI21_X1  g283(.A(new_n707), .B1(new_n708), .B2(G2105), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(new_n487), .B2(G119), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  MUX2_X1   g286(.A(G25), .B(new_n711), .S(G29), .Z(new_n712));
  XOR2_X1   g287(.A(KEYINPUT35), .B(G1991), .Z(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  MUX2_X1   g289(.A(G24), .B(G290), .S(G16), .Z(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(G1986), .Z(new_n716));
  NAND4_X1  g291(.A1(new_n703), .A2(new_n704), .A3(new_n714), .A4(new_n716), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT36), .ZN(new_n718));
  OR2_X1    g293(.A1(KEYINPUT30), .A2(G28), .ZN(new_n719));
  NAND2_X1  g294(.A1(KEYINPUT30), .A2(G28), .ZN(new_n720));
  AOI21_X1  g295(.A(G29), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  XOR2_X1   g296(.A(KEYINPUT31), .B(G11), .Z(new_n722));
  INV_X1    g297(.A(G34), .ZN(new_n723));
  AOI21_X1  g298(.A(G29), .B1(new_n723), .B2(KEYINPUT24), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(KEYINPUT24), .B2(new_n723), .ZN(new_n725));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n477), .B2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G2084), .ZN(new_n728));
  AOI211_X1 g303(.A(new_n721), .B(new_n722), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  OAI221_X1 g304(.A(new_n729), .B1(new_n726), .B2(new_n630), .C1(new_n728), .C2(new_n727), .ZN(new_n730));
  NAND3_X1  g305(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n731));
  INV_X1    g306(.A(KEYINPUT26), .ZN(new_n732));
  OR2_X1    g307(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n731), .A2(new_n732), .ZN(new_n734));
  AOI22_X1  g309(.A1(new_n733), .A2(new_n734), .B1(G105), .B2(new_n475), .ZN(new_n735));
  INV_X1    g310(.A(G141), .ZN(new_n736));
  INV_X1    g311(.A(G129), .ZN(new_n737));
  OAI221_X1 g312(.A(new_n735), .B1(new_n483), .B2(new_n736), .C1(new_n737), .C2(new_n486), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(G29), .ZN(new_n739));
  INV_X1    g314(.A(G32), .ZN(new_n740));
  OAI21_X1  g315(.A(new_n739), .B1(G29), .B2(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(new_n741), .ZN(new_n742));
  XNOR2_X1  g317(.A(KEYINPUT27), .B(G1996), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n730), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  AND2_X1   g319(.A1(new_n686), .A2(G21), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G286), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1966), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT96), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n726), .A2(G27), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G164), .B2(new_n726), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n751), .A2(G2078), .ZN(new_n752));
  AND2_X1   g327(.A1(new_n751), .A2(G2078), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n752), .B(new_n753), .C1(new_n746), .C2(new_n747), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n744), .A2(new_n749), .A3(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(new_n743), .ZN(new_n756));
  AND2_X1   g331(.A1(new_n726), .A2(G33), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n484), .A2(G139), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n472), .A2(G103), .A3(G2104), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n759), .A2(KEYINPUT95), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT25), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n504), .A2(G127), .ZN(new_n764));
  AND2_X1   g339(.A1(G115), .A2(G2104), .ZN(new_n765));
  OAI21_X1  g340(.A(G2105), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n758), .A2(new_n763), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g342(.A(new_n757), .B1(new_n767), .B2(G29), .ZN(new_n768));
  AOI22_X1  g343(.A1(new_n741), .A2(new_n756), .B1(new_n768), .B2(new_n442), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n686), .A2(G5), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(G171), .B2(new_n686), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n769), .B1(new_n442), .B2(new_n768), .C1(new_n771), .C2(G1961), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n755), .A2(new_n772), .ZN(new_n773));
  INV_X1    g348(.A(KEYINPUT98), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(G1961), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT97), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n773), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n774), .B1(new_n773), .B2(new_n776), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n686), .A2(G20), .ZN(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT23), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n607), .B2(new_n686), .ZN(new_n782));
  XOR2_X1   g357(.A(KEYINPUT100), .B(G1956), .Z(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n726), .A2(G35), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT99), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n491), .B2(G29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(KEYINPUT29), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n788), .B(G2090), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT93), .B(KEYINPUT28), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n726), .A2(G26), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(G128), .A2(new_n487), .B1(new_n484), .B2(G140), .ZN(new_n793));
  OAI21_X1  g368(.A(KEYINPUT90), .B1(G104), .B2(G2105), .ZN(new_n794));
  INV_X1    g369(.A(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(KEYINPUT90), .A2(G104), .A3(G2105), .ZN(new_n796));
  OAI221_X1 g371(.A(G2104), .B1(G116), .B2(new_n472), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n793), .A2(new_n798), .ZN(new_n799));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g376(.A1(new_n793), .A2(KEYINPUT92), .A3(new_n798), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g378(.A(new_n792), .B1(new_n803), .B2(G29), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2067), .ZN(new_n805));
  NOR2_X1   g380(.A1(G4), .A2(G16), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n611), .B2(G16), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT89), .B(G1348), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n686), .A2(G19), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n555), .B2(new_n686), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n811), .A2(G1341), .ZN(new_n812));
  OR2_X1    g387(.A1(new_n811), .A2(G1341), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n805), .A2(new_n809), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(KEYINPUT94), .ZN(new_n815));
  OAI211_X1 g390(.A(new_n784), .B(new_n789), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n815), .B2(new_n814), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n718), .A2(new_n779), .A3(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n611), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n822), .A2(new_n524), .ZN(new_n823));
  INV_X1    g398(.A(G93), .ZN(new_n824));
  INV_X1    g399(.A(G55), .ZN(new_n825));
  OAI22_X1  g400(.A1(new_n519), .A2(new_n824), .B1(new_n825), .B2(new_n522), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n555), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n827), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n614), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n821), .B(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT39), .ZN(new_n833));
  AOI21_X1  g408(.A(G860), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g409(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(G860), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT37), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n835), .A2(new_n837), .ZN(G145));
  NAND2_X1  g413(.A1(new_n767), .A2(KEYINPUT102), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n738), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n840), .A2(new_n803), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT101), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n842), .B1(new_n499), .B2(new_n502), .ZN(new_n843));
  OR2_X1    g418(.A1(G102), .A2(G2105), .ZN(new_n844));
  INV_X1    g419(.A(G114), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n845), .A2(G2105), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n844), .A2(new_n846), .A3(G2104), .ZN(new_n847));
  AND2_X1   g422(.A1(G126), .A2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n848), .B1(new_n463), .B2(new_n464), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n849), .A3(KEYINPUT101), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n843), .A2(new_n497), .A3(new_n508), .A4(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n840), .A2(new_n803), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n841), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n852), .B1(new_n841), .B2(new_n853), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  INV_X1    g432(.A(G118), .ZN(new_n858));
  AOI22_X1  g433(.A1(new_n857), .A2(KEYINPUT103), .B1(new_n858), .B2(G2105), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n859), .B1(KEYINPUT103), .B2(new_n857), .ZN(new_n860));
  INV_X1    g435(.A(G130), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n860), .B1(new_n486), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n862), .B1(G142), .B2(new_n484), .ZN(new_n863));
  XOR2_X1   g438(.A(new_n621), .B(new_n863), .Z(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n711), .ZN(new_n865));
  OAI22_X1  g440(.A1(new_n855), .A2(new_n856), .B1(KEYINPUT104), .B2(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n856), .ZN(new_n867));
  NOR2_X1   g442(.A1(new_n865), .A2(KEYINPUT104), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n867), .A2(new_n854), .A3(new_n868), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n630), .B(G160), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(G162), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n866), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n865), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n874), .B1(new_n855), .B2(new_n856), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n867), .A2(new_n854), .A3(new_n865), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n871), .ZN(new_n877));
  INV_X1    g452(.A(G37), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n873), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XOR2_X1   g454(.A(KEYINPUT105), .B(KEYINPUT40), .Z(new_n880));
  XNOR2_X1  g455(.A(new_n879), .B(new_n880), .ZN(G395));
  INV_X1    g456(.A(KEYINPUT109), .ZN(new_n882));
  OAI21_X1  g457(.A(new_n882), .B1(new_n827), .B2(G868), .ZN(new_n883));
  XNOR2_X1  g458(.A(G290), .B(G288), .ZN(new_n884));
  OR2_X1    g459(.A1(new_n884), .A2(KEYINPUT107), .ZN(new_n885));
  XNOR2_X1  g460(.A(G166), .B(KEYINPUT106), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n886), .B(G305), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n884), .A2(KEYINPUT107), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n885), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n886), .B(new_n697), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(KEYINPUT107), .A3(new_n884), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n892), .A2(KEYINPUT42), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n611), .A2(new_n607), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n598), .A2(new_n601), .B1(new_n570), .B2(new_n574), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n894), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n602), .A2(G299), .ZN(new_n899));
  OAI21_X1  g474(.A(KEYINPUT41), .B1(new_n899), .B2(new_n895), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n831), .A2(new_n610), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n831), .A2(new_n610), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n904), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n899), .A2(new_n895), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n906), .A2(new_n902), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n905), .A2(new_n908), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT108), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n892), .A2(KEYINPUT42), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n893), .A2(new_n909), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  AND2_X1   g487(.A1(new_n912), .A2(G868), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n893), .A2(new_n911), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n909), .A2(new_n910), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n905), .A2(new_n908), .A3(KEYINPUT108), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n883), .B1(new_n913), .B2(new_n917), .ZN(new_n918));
  AND4_X1   g493(.A1(KEYINPUT109), .A2(new_n917), .A3(G868), .A4(new_n912), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n918), .A2(new_n919), .ZN(G295));
  NOR2_X1   g495(.A1(new_n918), .A2(new_n919), .ZN(G331));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n922));
  INV_X1    g497(.A(new_n892), .ZN(new_n923));
  NAND2_X1  g498(.A1(G171), .A2(G168), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(G171), .A2(G168), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n831), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n926), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n928), .A2(new_n830), .A3(new_n828), .A4(new_n924), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n927), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n930), .A2(new_n901), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n927), .A2(new_n929), .A3(new_n907), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n923), .A2(new_n931), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(new_n878), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n907), .A2(KEYINPUT111), .A3(new_n897), .ZN(new_n935));
  OAI211_X1 g510(.A(new_n930), .B(new_n935), .C1(new_n901), .C2(KEYINPUT111), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n923), .B1(new_n936), .B2(new_n932), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT43), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n932), .ZN(new_n939));
  AOI22_X1  g514(.A1(new_n927), .A2(new_n929), .B1(new_n898), .B2(new_n900), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n892), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT110), .B(KEYINPUT43), .Z(new_n942));
  NAND4_X1  g517(.A1(new_n941), .A2(new_n933), .A3(new_n878), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n922), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n936), .A2(new_n932), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(new_n892), .ZN(new_n946));
  NAND4_X1  g521(.A1(new_n946), .A2(new_n878), .A3(new_n933), .A4(new_n942), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n941), .A2(new_n933), .A3(new_n878), .ZN(new_n948));
  INV_X1    g523(.A(new_n942), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n944), .B1(new_n951), .B2(new_n922), .ZN(G397));
  INV_X1    g527(.A(G2067), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n801), .A2(new_n953), .A3(new_n802), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n803), .A2(G2067), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  XNOR2_X1  g531(.A(new_n738), .B(new_n956), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n955), .A2(new_n954), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n706), .A2(new_n713), .A3(new_n710), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n954), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G1384), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n851), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT45), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n471), .A2(new_n476), .A3(G40), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n960), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(new_n711), .B(new_n713), .Z(new_n968));
  NOR2_X1   g543(.A1(new_n968), .A2(new_n958), .ZN(new_n969));
  INV_X1    g544(.A(new_n966), .ZN(new_n970));
  NOR2_X1   g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g546(.A1(G290), .A2(G1986), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT112), .Z(new_n973));
  NAND2_X1  g548(.A1(new_n973), .A2(new_n966), .ZN(new_n974));
  XOR2_X1   g549(.A(new_n974), .B(KEYINPUT48), .Z(new_n975));
  OAI21_X1  g550(.A(new_n967), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n955), .A2(new_n954), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n966), .B1(new_n977), .B2(new_n738), .ZN(new_n978));
  NAND2_X1  g553(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n966), .A2(new_n956), .ZN(new_n980));
  NOR2_X1   g555(.A1(KEYINPUT124), .A2(KEYINPUT46), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  OAI211_X1 g557(.A(new_n978), .B(new_n982), .C1(new_n979), .C2(new_n980), .ZN(new_n983));
  XNOR2_X1  g558(.A(KEYINPUT125), .B(KEYINPUT47), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  OR2_X1    g560(.A1(new_n983), .A2(new_n984), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n976), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n517), .A2(G61), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n524), .B1(new_n988), .B2(new_n589), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n587), .A2(new_n588), .ZN(new_n990));
  OAI21_X1  g565(.A(G1981), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT115), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  NAND3_X1  g568(.A1(G305), .A2(KEYINPUT115), .A3(G1981), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT114), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n996), .B1(G305), .B2(G1981), .ZN(new_n997));
  INV_X1    g572(.A(new_n989), .ZN(new_n998));
  INV_X1    g573(.A(new_n990), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  NAND4_X1  g575(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT114), .A4(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n997), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g577(.A(KEYINPUT49), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n962), .A2(KEYINPUT113), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n851), .A2(new_n1005), .A3(new_n961), .ZN(new_n1006));
  INV_X1    g581(.A(new_n965), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1003), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n995), .A2(new_n1002), .A3(KEYINPUT49), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(G288), .A2(G1976), .ZN(new_n1013));
  AOI22_X1  g588(.A1(new_n1012), .A2(new_n1013), .B1(new_n997), .B2(new_n1001), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n581), .B(G1976), .C1(new_n584), .C2(new_n585), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1008), .A2(G8), .A3(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT52), .ZN(new_n1017));
  INV_X1    g592(.A(G1976), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT52), .B1(G288), .B2(new_n1018), .ZN(new_n1019));
  NAND4_X1  g594(.A1(new_n1019), .A2(new_n1008), .A3(G8), .A4(new_n1015), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1012), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1004), .A2(new_n1022), .A3(new_n1006), .ZN(new_n1023));
  INV_X1    g598(.A(G2090), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n509), .A2(new_n961), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n965), .B1(KEYINPUT50), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1023), .A2(new_n1024), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n963), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n1007), .C1(new_n963), .C2(new_n962), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(new_n694), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1027), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1032));
  NAND3_X1  g607(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1033));
  INV_X1    g608(.A(new_n1033), .ZN(new_n1034));
  OAI211_X1 g609(.A(new_n1031), .B(G8), .C1(new_n1032), .C2(new_n1034), .ZN(new_n1035));
  OAI22_X1  g610(.A1(new_n1014), .A2(new_n1009), .B1(new_n1021), .B2(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n995), .A2(new_n1002), .A3(KEYINPUT49), .ZN(new_n1037));
  NOR3_X1   g612(.A1(new_n1037), .A2(new_n1003), .A3(new_n1009), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1034), .A2(new_n1032), .ZN(new_n1041));
  AND3_X1   g616(.A1(new_n851), .A2(new_n1005), .A3(new_n961), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n1005), .B1(new_n851), .B2(new_n961), .ZN(new_n1043));
  OAI21_X1  g618(.A(KEYINPUT50), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1025), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n965), .B1(new_n1045), .B2(new_n1022), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1044), .A2(new_n1024), .A3(new_n1046), .ZN(new_n1047));
  AND2_X1   g622(.A1(new_n1047), .A2(new_n1030), .ZN(new_n1048));
  INV_X1    g623(.A(G8), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1041), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(KEYINPUT45), .B1(new_n1004), .B2(new_n1006), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1007), .B1(new_n963), .B2(new_n1025), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n747), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1023), .A2(new_n728), .A3(new_n1026), .ZN(new_n1054));
  AOI211_X1 g629(.A(new_n1049), .B(G286), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1040), .A2(new_n1050), .A3(new_n1035), .A4(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT116), .B(KEYINPUT63), .Z(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AND3_X1   g633(.A1(new_n1023), .A2(new_n728), .A3(new_n1026), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n963), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n965), .B1(new_n1045), .B2(KEYINPUT45), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1966), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(G8), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT63), .ZN(new_n1064));
  NOR3_X1   g639(.A1(new_n1063), .A2(new_n1064), .A3(G286), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1031), .A2(G8), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1041), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1065), .A2(new_n1040), .A3(new_n1035), .A4(new_n1067), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1036), .B1(new_n1058), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1040), .A2(new_n1050), .A3(new_n1035), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1042), .A2(new_n1043), .A3(KEYINPUT50), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1026), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT119), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(G1961), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT119), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1023), .A2(new_n1075), .A3(new_n1026), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1074), .A3(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT53), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1029), .B2(G2078), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n1060), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n1061), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1077), .A2(new_n1079), .A3(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(G171), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1070), .A2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G286), .A2(G8), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT121), .B1(new_n1059), .B2(new_n1062), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT121), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1053), .A2(new_n1086), .A3(new_n1054), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1084), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1085), .A2(G168), .A3(new_n1087), .ZN(new_n1089));
  AND2_X1   g664(.A1(KEYINPUT51), .A2(G8), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT51), .B1(G286), .B2(G8), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1063), .A2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g668(.A(new_n1088), .B1(new_n1091), .B2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT62), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1083), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  AOI22_X1  g671(.A1(new_n1089), .A2(new_n1090), .B1(new_n1063), .B2(new_n1092), .ZN(new_n1097));
  NOR3_X1   g672(.A1(new_n1097), .A2(KEYINPUT62), .A3(new_n1088), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1069), .B1(new_n1096), .B2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1008), .A2(KEYINPUT118), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1008), .A2(KEYINPUT118), .ZN(new_n1102));
  XOR2_X1   g677(.A(KEYINPUT58), .B(G1341), .Z(new_n1103));
  NAND3_X1  g678(.A1(new_n1101), .A2(new_n1102), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1104), .B1(G1996), .B2(new_n1029), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n555), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT59), .ZN(new_n1107));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1108), .A3(new_n555), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1107), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g685(.A(new_n1102), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n953), .B1(new_n1111), .B2(new_n1100), .ZN(new_n1112));
  INV_X1    g687(.A(G1348), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1073), .A2(new_n1113), .A3(new_n1076), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1112), .A2(new_n602), .A3(new_n1114), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n602), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1116));
  OAI21_X1  g691(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  XNOR2_X1  g692(.A(KEYINPUT56), .B(G2072), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1118), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1029), .A2(new_n1119), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1121), .B2(G1956), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n574), .A2(new_n566), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT117), .B(KEYINPUT57), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1125), .B1(G299), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1122), .A2(new_n1128), .ZN(new_n1129));
  OAI211_X1 g704(.A(new_n1127), .B(new_n1120), .C1(new_n1121), .C2(G1956), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1129), .A2(KEYINPUT120), .A3(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT61), .ZN(new_n1132));
  INV_X1    g707(.A(KEYINPUT120), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1122), .A2(new_n1133), .A3(new_n1128), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1131), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(KEYINPUT61), .A3(new_n1130), .ZN(new_n1136));
  NOR2_X1   g711(.A1(new_n602), .A2(KEYINPUT60), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1112), .A2(new_n1114), .A3(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND4_X1  g714(.A1(new_n1110), .A2(new_n1117), .A3(new_n1135), .A4(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1129), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1130), .B1(new_n1141), .B2(new_n1116), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1070), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1077), .A2(G301), .A3(new_n1079), .A4(new_n1080), .ZN(new_n1145));
  INV_X1    g720(.A(new_n962), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n965), .B1(new_n1146), .B2(KEYINPUT45), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1147), .A2(KEYINPUT53), .A3(new_n443), .A4(new_n964), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1077), .A2(new_n1079), .A3(new_n1148), .ZN(new_n1149));
  OAI211_X1 g724(.A(KEYINPUT54), .B(new_n1145), .C1(new_n1149), .C2(G301), .ZN(new_n1150));
  OAI211_X1 g725(.A(new_n1144), .B(new_n1150), .C1(new_n1088), .C2(new_n1097), .ZN(new_n1151));
  XOR2_X1   g726(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1152));
  NAND4_X1  g727(.A1(new_n1077), .A2(G301), .A3(new_n1079), .A4(new_n1148), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1152), .B1(new_n1082), .B2(new_n1153), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1154), .A2(KEYINPUT123), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT123), .ZN(new_n1156));
  AOI211_X1 g731(.A(new_n1156), .B(new_n1152), .C1(new_n1082), .C2(new_n1153), .ZN(new_n1157));
  NOR3_X1   g732(.A1(new_n1151), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1099), .B1(new_n1143), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g734(.A(new_n973), .B1(G1986), .B2(G290), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n970), .B1(new_n969), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n987), .B1(new_n1159), .B2(new_n1161), .ZN(G329));
  assign    G231 = 1'b0;
  NAND2_X1  g737(.A1(new_n947), .A2(new_n950), .ZN(new_n1164));
  INV_X1    g738(.A(G319), .ZN(new_n1165));
  NOR3_X1   g739(.A1(G401), .A2(new_n1165), .A3(G227), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1166), .B1(new_n683), .B2(new_n684), .ZN(new_n1167));
  NAND2_X1  g741(.A1(new_n1167), .A2(KEYINPUT126), .ZN(new_n1168));
  INV_X1    g742(.A(KEYINPUT126), .ZN(new_n1169));
  OAI211_X1 g743(.A(new_n1169), .B(new_n1166), .C1(new_n683), .C2(new_n684), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND3_X1  g745(.A1(new_n1164), .A2(new_n1171), .A3(new_n879), .ZN(G225));
  INV_X1    g746(.A(G225), .ZN(G308));
endmodule


