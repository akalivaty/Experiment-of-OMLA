

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584;

  XOR2_X1 U323 ( .A(n345), .B(n344), .Z(n579) );
  XNOR2_X1 U324 ( .A(n407), .B(KEYINPUT113), .ZN(n408) );
  XNOR2_X1 U325 ( .A(KEYINPUT48), .B(KEYINPUT115), .ZN(n419) );
  XOR2_X1 U326 ( .A(n335), .B(n334), .Z(n291) );
  XOR2_X1 U327 ( .A(n340), .B(n374), .Z(n292) );
  XNOR2_X1 U328 ( .A(n409), .B(n408), .ZN(n418) );
  XNOR2_X1 U329 ( .A(n435), .B(KEYINPUT121), .ZN(n436) );
  XNOR2_X1 U330 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U331 ( .A(n370), .B(n369), .ZN(n373) );
  XNOR2_X1 U332 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U333 ( .A(n381), .B(n380), .ZN(n413) );
  NOR2_X1 U334 ( .A1(n569), .A2(n568), .ZN(n581) );
  XNOR2_X1 U335 ( .A(n364), .B(n363), .ZN(n570) );
  XNOR2_X1 U336 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U337 ( .A(n464), .B(n463), .ZN(G1349GAT) );
  XOR2_X1 U338 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n294) );
  XNOR2_X1 U339 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n293) );
  XNOR2_X1 U340 ( .A(n294), .B(n293), .ZN(n429) );
  XOR2_X1 U341 ( .A(G120GAT), .B(G71GAT), .Z(n375) );
  XOR2_X1 U342 ( .A(n429), .B(n375), .Z(n296) );
  XNOR2_X1 U343 ( .A(G43GAT), .B(G190GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U345 ( .A(G183GAT), .B(G176GAT), .Z(n298) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U347 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U348 ( .A(n300), .B(n299), .Z(n305) );
  XOR2_X1 U349 ( .A(KEYINPUT90), .B(KEYINPUT20), .Z(n302) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(KEYINPUT89), .ZN(n301) );
  XNOR2_X1 U351 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U352 ( .A(G15GAT), .B(n303), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U354 ( .A(KEYINPUT88), .B(G134GAT), .Z(n307) );
  XNOR2_X1 U355 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n306) );
  XNOR2_X1 U356 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U357 ( .A(G113GAT), .B(n308), .ZN(n450) );
  XOR2_X1 U358 ( .A(n309), .B(n450), .Z(n524) );
  INV_X1 U359 ( .A(n524), .ZN(n532) );
  XOR2_X1 U360 ( .A(KEYINPUT3), .B(KEYINPUT94), .Z(n311) );
  XNOR2_X1 U361 ( .A(KEYINPUT93), .B(G155GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U363 ( .A(KEYINPUT2), .B(n312), .Z(n443) );
  XOR2_X1 U364 ( .A(KEYINPUT92), .B(G218GAT), .Z(n314) );
  XNOR2_X1 U365 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U367 ( .A(G197GAT), .B(n315), .Z(n432) );
  XNOR2_X1 U368 ( .A(n443), .B(n432), .ZN(n327) );
  XOR2_X1 U369 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n317) );
  XNOR2_X1 U370 ( .A(G204GAT), .B(KEYINPUT91), .ZN(n316) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U372 ( .A(G50GAT), .B(G162GAT), .Z(n399) );
  XOR2_X1 U373 ( .A(n318), .B(n399), .Z(n325) );
  XOR2_X1 U374 ( .A(G141GAT), .B(G22GAT), .Z(n349) );
  XOR2_X1 U375 ( .A(G78GAT), .B(G148GAT), .Z(n320) );
  XNOR2_X1 U376 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n319) );
  XNOR2_X1 U377 ( .A(n320), .B(n319), .ZN(n371) );
  XOR2_X1 U378 ( .A(KEYINPUT22), .B(n371), .Z(n322) );
  NAND2_X1 U379 ( .A1(G228GAT), .A2(G233GAT), .ZN(n321) );
  XNOR2_X1 U380 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n349), .B(n323), .ZN(n324) );
  XNOR2_X1 U382 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U383 ( .A(n327), .B(n326), .ZN(n468) );
  XOR2_X1 U384 ( .A(KEYINPUT14), .B(KEYINPUT85), .Z(n329) );
  XNOR2_X1 U385 ( .A(KEYINPUT83), .B(KEYINPUT84), .ZN(n328) );
  XNOR2_X1 U386 ( .A(n329), .B(n328), .ZN(n345) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G211GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G22GAT), .B(G155GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U390 ( .A(KEYINPUT12), .B(KEYINPUT82), .Z(n333) );
  XNOR2_X1 U391 ( .A(G127GAT), .B(G71GAT), .ZN(n332) );
  XNOR2_X1 U392 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U393 ( .A(KEYINPUT86), .B(G64GAT), .Z(n337) );
  NAND2_X1 U394 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U395 ( .A(n337), .B(n336), .ZN(n338) );
  XNOR2_X1 U396 ( .A(KEYINPUT15), .B(n338), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n291), .B(n339), .ZN(n340) );
  XOR2_X1 U398 ( .A(KEYINPUT13), .B(G57GAT), .Z(n374) );
  XOR2_X1 U399 ( .A(G1GAT), .B(KEYINPUT70), .Z(n342) );
  XNOR2_X1 U400 ( .A(G15GAT), .B(KEYINPUT71), .ZN(n341) );
  XNOR2_X1 U401 ( .A(n342), .B(n341), .ZN(n360) );
  XOR2_X1 U402 ( .A(G8GAT), .B(G183GAT), .Z(n424) );
  XNOR2_X1 U403 ( .A(n360), .B(n424), .ZN(n343) );
  XNOR2_X1 U404 ( .A(n292), .B(n343), .ZN(n344) );
  XOR2_X1 U405 ( .A(G113GAT), .B(G197GAT), .Z(n347) );
  XNOR2_X1 U406 ( .A(G36GAT), .B(G50GAT), .ZN(n346) );
  XNOR2_X1 U407 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U408 ( .A(n349), .B(n348), .Z(n351) );
  NAND2_X1 U409 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n364) );
  XOR2_X1 U411 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n353) );
  XNOR2_X1 U412 ( .A(KEYINPUT30), .B(KEYINPUT67), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U414 ( .A(KEYINPUT29), .B(KEYINPUT68), .Z(n355) );
  XNOR2_X1 U415 ( .A(G169GAT), .B(G8GAT), .ZN(n354) );
  XNOR2_X1 U416 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U417 ( .A(n357), .B(n356), .Z(n362) );
  XOR2_X1 U418 ( .A(G29GAT), .B(G43GAT), .Z(n359) );
  XNOR2_X1 U419 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n393) );
  XNOR2_X1 U421 ( .A(n393), .B(n360), .ZN(n361) );
  XNOR2_X1 U422 ( .A(n362), .B(n361), .ZN(n363) );
  XOR2_X1 U423 ( .A(G64GAT), .B(G92GAT), .Z(n366) );
  XNOR2_X1 U424 ( .A(G176GAT), .B(G204GAT), .ZN(n365) );
  XNOR2_X1 U425 ( .A(n366), .B(n365), .ZN(n428) );
  XOR2_X1 U426 ( .A(G99GAT), .B(G85GAT), .Z(n388) );
  XOR2_X1 U427 ( .A(n428), .B(n388), .Z(n370) );
  NAND2_X1 U428 ( .A1(G230GAT), .A2(G233GAT), .ZN(n368) );
  INV_X1 U429 ( .A(KEYINPUT75), .ZN(n367) );
  XNOR2_X1 U430 ( .A(n371), .B(KEYINPUT76), .ZN(n372) );
  XNOR2_X1 U431 ( .A(n373), .B(n372), .ZN(n381) );
  XOR2_X1 U432 ( .A(n375), .B(n374), .Z(n379) );
  XOR2_X1 U433 ( .A(KEYINPUT33), .B(KEYINPUT32), .Z(n377) );
  XNOR2_X1 U434 ( .A(KEYINPUT73), .B(KEYINPUT31), .ZN(n376) );
  XNOR2_X1 U435 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U436 ( .A(n413), .B(KEYINPUT41), .ZN(n551) );
  AND2_X1 U437 ( .A1(n570), .A2(n551), .ZN(n383) );
  XOR2_X1 U438 ( .A(KEYINPUT111), .B(KEYINPUT46), .Z(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  NOR2_X1 U440 ( .A1(n579), .A2(n384), .ZN(n385) );
  XNOR2_X1 U441 ( .A(n385), .B(KEYINPUT112), .ZN(n406) );
  XOR2_X1 U442 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n387) );
  XNOR2_X1 U443 ( .A(G92GAT), .B(KEYINPUT65), .ZN(n386) );
  XNOR2_X1 U444 ( .A(n387), .B(n386), .ZN(n389) );
  XOR2_X1 U445 ( .A(n389), .B(n388), .Z(n391) );
  XNOR2_X1 U446 ( .A(G218GAT), .B(G106GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n392) );
  XOR2_X1 U448 ( .A(n392), .B(KEYINPUT78), .Z(n395) );
  XNOR2_X1 U449 ( .A(n393), .B(G134GAT), .ZN(n394) );
  XNOR2_X1 U450 ( .A(n395), .B(n394), .ZN(n405) );
  XOR2_X1 U451 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n397) );
  XNOR2_X1 U452 ( .A(KEYINPUT10), .B(KEYINPUT77), .ZN(n396) );
  XNOR2_X1 U453 ( .A(n397), .B(n396), .ZN(n403) );
  XNOR2_X1 U454 ( .A(G36GAT), .B(G190GAT), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n398), .B(KEYINPUT81), .ZN(n421) );
  XOR2_X1 U456 ( .A(n421), .B(n399), .Z(n401) );
  NAND2_X1 U457 ( .A1(G232GAT), .A2(G233GAT), .ZN(n400) );
  XNOR2_X1 U458 ( .A(n401), .B(n400), .ZN(n402) );
  XOR2_X1 U459 ( .A(n403), .B(n402), .Z(n404) );
  XNOR2_X1 U460 ( .A(n405), .B(n404), .ZN(n542) );
  NAND2_X1 U461 ( .A1(n406), .A2(n542), .ZN(n409) );
  INV_X1 U462 ( .A(KEYINPUT47), .ZN(n407) );
  XNOR2_X1 U463 ( .A(KEYINPUT36), .B(KEYINPUT107), .ZN(n410) );
  XNOR2_X1 U464 ( .A(n410), .B(n542), .ZN(n582) );
  NAND2_X1 U465 ( .A1(n579), .A2(n582), .ZN(n412) );
  XOR2_X1 U466 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n411) );
  XNOR2_X1 U467 ( .A(n412), .B(n411), .ZN(n414) );
  NAND2_X1 U468 ( .A1(n414), .A2(n413), .ZN(n415) );
  NOR2_X1 U469 ( .A1(n570), .A2(n415), .ZN(n416) );
  XNOR2_X1 U470 ( .A(KEYINPUT114), .B(n416), .ZN(n417) );
  NOR2_X1 U471 ( .A1(n418), .A2(n417), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n530) );
  XOR2_X1 U473 ( .A(n421), .B(KEYINPUT99), .Z(n423) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n423), .B(n422), .ZN(n427) );
  XNOR2_X1 U476 ( .A(n424), .B(KEYINPUT100), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n425), .B(KEYINPUT98), .ZN(n426) );
  XOR2_X1 U478 ( .A(n427), .B(n426), .Z(n431) );
  XNOR2_X1 U479 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U480 ( .A(n431), .B(n430), .ZN(n434) );
  INV_X1 U481 ( .A(n432), .ZN(n433) );
  XOR2_X1 U482 ( .A(n434), .B(n433), .Z(n501) );
  INV_X1 U483 ( .A(n501), .ZN(n521) );
  NAND2_X1 U484 ( .A1(n530), .A2(n521), .ZN(n435) );
  XNOR2_X1 U485 ( .A(n436), .B(KEYINPUT54), .ZN(n457) );
  XOR2_X1 U486 ( .A(KEYINPUT96), .B(KEYINPUT97), .Z(n438) );
  XNOR2_X1 U487 ( .A(KEYINPUT1), .B(KEYINPUT4), .ZN(n437) );
  XNOR2_X1 U488 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U489 ( .A(KEYINPUT5), .B(n439), .Z(n441) );
  NAND2_X1 U490 ( .A1(G225GAT), .A2(G233GAT), .ZN(n440) );
  XNOR2_X1 U491 ( .A(n441), .B(n440), .ZN(n442) );
  XOR2_X1 U492 ( .A(n442), .B(KEYINPUT6), .Z(n445) );
  XNOR2_X1 U493 ( .A(n443), .B(KEYINPUT95), .ZN(n444) );
  XNOR2_X1 U494 ( .A(n445), .B(n444), .ZN(n449) );
  XOR2_X1 U495 ( .A(G85GAT), .B(G162GAT), .Z(n447) );
  XNOR2_X1 U496 ( .A(G29GAT), .B(G141GAT), .ZN(n446) );
  XNOR2_X1 U497 ( .A(n447), .B(n446), .ZN(n448) );
  XOR2_X1 U498 ( .A(n449), .B(n448), .Z(n456) );
  INV_X1 U499 ( .A(n450), .ZN(n454) );
  XOR2_X1 U500 ( .A(G57GAT), .B(G148GAT), .Z(n452) );
  XNOR2_X1 U501 ( .A(G1GAT), .B(G120GAT), .ZN(n451) );
  XNOR2_X1 U502 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U503 ( .A(n454), .B(n453), .ZN(n455) );
  XNOR2_X1 U504 ( .A(n456), .B(n455), .ZN(n498) );
  NAND2_X1 U505 ( .A1(n457), .A2(n498), .ZN(n458) );
  XNOR2_X1 U506 ( .A(n458), .B(KEYINPUT64), .ZN(n569) );
  NOR2_X1 U507 ( .A1(n468), .A2(n569), .ZN(n459) );
  XNOR2_X1 U508 ( .A(n459), .B(KEYINPUT55), .ZN(n460) );
  NOR2_X2 U509 ( .A1(n532), .A2(n460), .ZN(n565) );
  NAND2_X1 U510 ( .A1(n565), .A2(n551), .ZN(n464) );
  XOR2_X1 U511 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n462) );
  XNOR2_X1 U512 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n461) );
  XNOR2_X1 U513 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n482) );
  INV_X1 U514 ( .A(n498), .ZN(n546) );
  NAND2_X1 U515 ( .A1(n413), .A2(n570), .ZN(n495) );
  XOR2_X1 U516 ( .A(n468), .B(KEYINPUT28), .Z(n506) );
  XNOR2_X1 U517 ( .A(n521), .B(KEYINPUT27), .ZN(n470) );
  NAND2_X1 U518 ( .A1(n506), .A2(n470), .ZN(n465) );
  NOR2_X1 U519 ( .A1(n498), .A2(n465), .ZN(n531) );
  NAND2_X1 U520 ( .A1(n531), .A2(n532), .ZN(n475) );
  NOR2_X1 U521 ( .A1(n532), .A2(n501), .ZN(n466) );
  NOR2_X1 U522 ( .A1(n468), .A2(n466), .ZN(n467) );
  XNOR2_X1 U523 ( .A(KEYINPUT25), .B(n467), .ZN(n472) );
  NAND2_X1 U524 ( .A1(n468), .A2(n532), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT26), .ZN(n568) );
  INV_X1 U526 ( .A(n568), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n548) );
  NAND2_X1 U528 ( .A1(n472), .A2(n548), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n473), .A2(n498), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n476) );
  XNOR2_X1 U531 ( .A(n476), .B(KEYINPUT101), .ZN(n492) );
  XOR2_X1 U532 ( .A(KEYINPUT87), .B(KEYINPUT16), .Z(n478) );
  NAND2_X1 U533 ( .A1(n579), .A2(n542), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(n479) );
  OR2_X1 U535 ( .A1(n492), .A2(n479), .ZN(n509) );
  NOR2_X1 U536 ( .A1(n495), .A2(n509), .ZN(n480) );
  XNOR2_X1 U537 ( .A(KEYINPUT102), .B(n480), .ZN(n488) );
  NAND2_X1 U538 ( .A1(n546), .A2(n488), .ZN(n481) );
  XNOR2_X1 U539 ( .A(n482), .B(n481), .ZN(G1324GAT) );
  XOR2_X1 U540 ( .A(G8GAT), .B(KEYINPUT103), .Z(n484) );
  NAND2_X1 U541 ( .A1(n521), .A2(n488), .ZN(n483) );
  XNOR2_X1 U542 ( .A(n484), .B(n483), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(KEYINPUT104), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U544 ( .A1(n488), .A2(n524), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(n487), .ZN(G1326GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n490) );
  INV_X1 U548 ( .A(n506), .ZN(n527) );
  NAND2_X1 U549 ( .A1(n488), .A2(n527), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n491), .ZN(G1327GAT) );
  NOR2_X1 U552 ( .A1(n579), .A2(n492), .ZN(n493) );
  NAND2_X1 U553 ( .A1(n582), .A2(n493), .ZN(n494) );
  XOR2_X1 U554 ( .A(KEYINPUT37), .B(n494), .Z(n519) );
  NOR2_X1 U555 ( .A1(n519), .A2(n495), .ZN(n497) );
  XOR2_X1 U556 ( .A(KEYINPUT108), .B(KEYINPUT38), .Z(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(n505) );
  NOR2_X1 U558 ( .A1(n498), .A2(n505), .ZN(n500) );
  XNOR2_X1 U559 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U561 ( .A1(n501), .A2(n505), .ZN(n502) );
  XOR2_X1 U562 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U563 ( .A1(n532), .A2(n505), .ZN(n503) );
  XOR2_X1 U564 ( .A(KEYINPUT40), .B(n503), .Z(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NOR2_X1 U566 ( .A1(n506), .A2(n505), .ZN(n507) );
  XOR2_X1 U567 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  XNOR2_X1 U568 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n511) );
  INV_X1 U569 ( .A(n570), .ZN(n508) );
  NAND2_X1 U570 ( .A1(n508), .A2(n551), .ZN(n518) );
  NOR2_X1 U571 ( .A1(n509), .A2(n518), .ZN(n514) );
  NAND2_X1 U572 ( .A1(n514), .A2(n546), .ZN(n510) );
  XNOR2_X1 U573 ( .A(n511), .B(n510), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n514), .A2(n521), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U576 ( .A1(n524), .A2(n514), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U578 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n516) );
  NAND2_X1 U579 ( .A1(n514), .A2(n527), .ZN(n515) );
  XNOR2_X1 U580 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U581 ( .A(G78GAT), .B(n517), .Z(G1335GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n518), .ZN(n526) );
  NAND2_X1 U583 ( .A1(n526), .A2(n546), .ZN(n520) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n520), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n526), .A2(n521), .ZN(n522) );
  XNOR2_X1 U586 ( .A(n522), .B(KEYINPUT110), .ZN(n523) );
  XNOR2_X1 U587 ( .A(G92GAT), .B(n523), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n526), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U590 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U591 ( .A(n528), .B(KEYINPUT44), .ZN(n529) );
  XNOR2_X1 U592 ( .A(G106GAT), .B(n529), .ZN(G1339GAT) );
  XOR2_X1 U593 ( .A(G113GAT), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U594 ( .A1(n530), .A2(n531), .ZN(n533) );
  NOR2_X1 U595 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(KEYINPUT116), .ZN(n543) );
  NAND2_X1 U597 ( .A1(n543), .A2(n570), .ZN(n535) );
  XNOR2_X1 U598 ( .A(n536), .B(n535), .ZN(G1340GAT) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U600 ( .A1(n543), .A2(n551), .ZN(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n540) );
  NAND2_X1 U603 ( .A1(n579), .A2(n543), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(n541) );
  XOR2_X1 U605 ( .A(G127GAT), .B(n541), .Z(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  INV_X1 U607 ( .A(n542), .ZN(n564) );
  NAND2_X1 U608 ( .A1(n564), .A2(n543), .ZN(n544) );
  XNOR2_X1 U609 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  XOR2_X1 U610 ( .A(G141GAT), .B(KEYINPUT119), .Z(n550) );
  NAND2_X1 U611 ( .A1(n530), .A2(n546), .ZN(n547) );
  NOR2_X1 U612 ( .A1(n548), .A2(n547), .ZN(n557) );
  NAND2_X1 U613 ( .A1(n557), .A2(n570), .ZN(n549) );
  XNOR2_X1 U614 ( .A(n550), .B(n549), .ZN(G1344GAT) );
  XOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U616 ( .A1(n557), .A2(n551), .ZN(n552) );
  XNOR2_X1 U617 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U618 ( .A(G148GAT), .B(n554), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n557), .A2(n579), .ZN(n555) );
  XNOR2_X1 U620 ( .A(n555), .B(KEYINPUT120), .ZN(n556) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n556), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n557), .A2(n564), .ZN(n558) );
  XNOR2_X1 U623 ( .A(n558), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n565), .A2(n570), .ZN(n559) );
  XNOR2_X1 U625 ( .A(n559), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U626 ( .A(G183GAT), .B(KEYINPUT123), .Z(n561) );
  NAND2_X1 U627 ( .A1(n565), .A2(n579), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1350GAT) );
  XNOR2_X1 U629 ( .A(G190GAT), .B(KEYINPUT125), .ZN(n562) );
  XNOR2_X1 U630 ( .A(n562), .B(KEYINPUT124), .ZN(n563) );
  XOR2_X1 U631 ( .A(KEYINPUT58), .B(n563), .Z(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1351GAT) );
  NAND2_X1 U634 ( .A1(n570), .A2(n581), .ZN(n574) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n577) );
  INV_X1 U640 ( .A(n413), .ZN(n575) );
  NAND2_X1 U641 ( .A1(n581), .A2(n575), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U643 ( .A(G204GAT), .B(n578), .Z(G1353GAT) );
  NAND2_X1 U644 ( .A1(n581), .A2(n579), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(n583), .B(KEYINPUT62), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

