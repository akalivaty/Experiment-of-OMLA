//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 0 1 0 1 0 0 0 1 0 1 1 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n873, new_n874, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n1000, new_n1001;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  NAND2_X1  g005(.A1(G229gat), .A2(G233gat), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT13), .Z(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT89), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n212));
  AOI22_X1  g011(.A1(new_n210), .A2(new_n211), .B1(new_n212), .B2(new_n209), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT89), .A3(G1gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT90), .ZN(new_n215));
  INV_X1    g014(.A(G8gat), .ZN(new_n216));
  AOI22_X1  g015(.A1(new_n213), .A2(new_n214), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n217), .B1(new_n215), .B2(new_n216), .ZN(new_n218));
  NAND4_X1  g017(.A1(new_n213), .A2(KEYINPUT90), .A3(G8gat), .A4(new_n214), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n218), .A2(KEYINPUT91), .A3(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT91), .B1(new_n218), .B2(new_n219), .ZN(new_n222));
  XNOR2_X1  g021(.A(KEYINPUT88), .B(G36gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G29gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT14), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n225), .B1(G29gat), .B2(G36gat), .ZN(new_n226));
  OR3_X1    g025(.A1(new_n225), .A2(G29gat), .A3(G36gat), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n224), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT15), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n224), .A2(KEYINPUT15), .A3(new_n226), .A4(new_n227), .ZN(new_n231));
  XNOR2_X1  g030(.A(G43gat), .B(G50gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n230), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n231), .A2(new_n232), .ZN(new_n234));
  AND2_X1   g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NOR3_X1   g034(.A1(new_n221), .A2(new_n222), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n233), .A2(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n218), .A2(new_n219), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT91), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n237), .B1(new_n240), .B2(new_n220), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n208), .B1(new_n236), .B2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT92), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n237), .A3(new_n220), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n237), .A2(KEYINPUT17), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT17), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n246), .B1(new_n233), .B2(new_n234), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n238), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n244), .A2(new_n207), .A3(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT18), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n206), .B1(new_n243), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n240), .A2(new_n220), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(new_n235), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n254), .A2(new_n244), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n255), .A2(KEYINPUT92), .A3(new_n208), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT92), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n242), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n249), .B(KEYINPUT18), .ZN(new_n260));
  INV_X1    g059(.A(new_n206), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(KEYINPUT71), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT71), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT1), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(G127gat), .B(G134gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(G113gat), .B(G120gat), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n268), .B(new_n269), .C1(new_n270), .C2(KEYINPUT70), .ZN(new_n271));
  INV_X1    g070(.A(G113gat), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(G120gat), .ZN(new_n273));
  INV_X1    g072(.A(G120gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n274), .A2(G113gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT70), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(G127gat), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT69), .B(G134gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(new_n278), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n270), .A2(KEYINPUT1), .ZN(new_n283));
  OAI22_X1  g082(.A1(new_n271), .A2(new_n277), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G169gat), .ZN(new_n286));
  INV_X1    g085(.A(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT26), .ZN(new_n289));
  NAND2_X1  g088(.A1(G169gat), .A2(G176gat), .ZN(new_n290));
  AND3_X1   g089(.A1(new_n288), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G183gat), .A2(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n292), .B1(new_n288), .B2(new_n289), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n291), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT67), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(G190gat), .ZN(new_n298));
  AND2_X1   g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  XNOR2_X1  g098(.A(KEYINPUT27), .B(G183gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n299), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n299), .A2(new_n300), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n304));
  OAI211_X1 g103(.A(new_n294), .B(new_n302), .C1(new_n303), .C2(new_n304), .ZN(new_n305));
  AND2_X1   g104(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n306));
  NOR2_X1   g105(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n288), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI211_X1 g109(.A(new_n288), .B(KEYINPUT66), .C1(new_n306), .C2(new_n307), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n290), .B1(new_n288), .B2(new_n313), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT64), .B1(G183gat), .B2(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  NOR3_X1   g115(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n292), .A2(KEYINPUT24), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT24), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n320), .A2(G183gat), .A3(G190gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n314), .B1(new_n318), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT25), .B1(new_n312), .B2(new_n323), .ZN(new_n324));
  OAI211_X1 g123(.A(KEYINPUT25), .B(new_n290), .C1(new_n288), .C2(new_n313), .ZN(new_n325));
  INV_X1    g124(.A(G183gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n296), .A2(new_n298), .A3(new_n326), .ZN(new_n327));
  AOI221_X4 g126(.A(new_n325), .B1(new_n322), .B2(new_n327), .C1(new_n310), .C2(new_n311), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n285), .B(new_n305), .C1(new_n324), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n329), .A2(KEYINPUT72), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT25), .ZN(new_n331));
  INV_X1    g130(.A(new_n311), .ZN(new_n332));
  XNOR2_X1  g131(.A(KEYINPUT65), .B(KEYINPUT23), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT66), .B1(new_n333), .B2(new_n288), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(new_n317), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n322), .A2(new_n336), .A3(new_n315), .ZN(new_n337));
  INV_X1    g136(.A(new_n314), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n331), .B1(new_n335), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n325), .B1(new_n322), .B2(new_n327), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n341), .A2(new_n312), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT72), .ZN(new_n344));
  NAND4_X1  g143(.A1(new_n343), .A2(new_n344), .A3(new_n285), .A4(new_n305), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n305), .B1(new_n324), .B2(new_n328), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(new_n284), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n330), .A2(new_n345), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT73), .ZN(new_n349));
  NAND2_X1  g148(.A1(G227gat), .A2(G233gat), .ZN(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  AND3_X1   g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(new_n349), .B1(new_n348), .B2(new_n351), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT32), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT33), .ZN(new_n355));
  OAI21_X1  g154(.A(new_n355), .B1(new_n352), .B2(new_n353), .ZN(new_n356));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT74), .ZN(new_n358));
  XNOR2_X1  g157(.A(G71gat), .B(G99gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n354), .A2(new_n356), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(KEYINPUT33), .ZN(new_n362));
  OAI211_X1 g161(.A(KEYINPUT32), .B(new_n362), .C1(new_n352), .C2(new_n353), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n330), .A2(new_n345), .A3(new_n347), .A4(new_n350), .ZN(new_n364));
  XOR2_X1   g163(.A(new_n364), .B(KEYINPUT34), .Z(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n354), .A2(new_n356), .A3(new_n360), .ZN(new_n368));
  AOI21_X1  g167(.A(new_n365), .B1(new_n368), .B2(new_n363), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT36), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n365), .ZN(new_n371));
  INV_X1    g170(.A(new_n363), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n371), .B1(new_n361), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT36), .ZN(new_n374));
  INV_X1    g173(.A(new_n366), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(new_n368), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(G155gat), .B(G162gat), .ZN(new_n378));
  INV_X1    g177(.A(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G141gat), .ZN(new_n380));
  INV_X1    g179(.A(G148gat), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT2), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n383), .A2(KEYINPUT77), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT77), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT2), .ZN(new_n386));
  NAND2_X1  g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387));
  NAND4_X1  g186(.A1(new_n382), .A2(new_n384), .A3(new_n386), .A4(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n379), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(G155gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n390), .A2(KEYINPUT78), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(G155gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n391), .A2(new_n393), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n383), .B1(new_n394), .B2(G162gat), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n378), .A2(new_n382), .A3(new_n387), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n389), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n284), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT80), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n270), .A2(KEYINPUT70), .ZN(new_n400));
  OAI21_X1  g199(.A(new_n276), .B1(new_n273), .B2(new_n275), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n400), .A2(new_n401), .A3(new_n269), .A4(new_n268), .ZN(new_n402));
  XNOR2_X1  g201(.A(KEYINPUT78), .B(G155gat), .ZN(new_n403));
  INV_X1    g202(.A(G162gat), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT2), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(G155gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n390), .A2(G162gat), .ZN(new_n407));
  AND4_X1   g206(.A1(new_n406), .A2(new_n382), .A3(new_n407), .A4(new_n387), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n405), .A2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n264), .B1(new_n273), .B2(new_n275), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT69), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n411), .A2(G134gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n279), .A2(KEYINPUT69), .ZN(new_n413));
  OAI21_X1  g212(.A(G127gat), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n414), .A3(new_n280), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n402), .A2(new_n409), .A3(new_n415), .A4(new_n389), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n398), .A2(new_n399), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(G225gat), .A2(G233gat), .ZN(new_n418));
  INV_X1    g217(.A(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n284), .A2(new_n397), .A3(KEYINPUT80), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n417), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT81), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  AOI22_X1  g222(.A1(new_n397), .A2(KEYINPUT3), .B1(new_n402), .B2(new_n415), .ZN(new_n424));
  AOI22_X1  g223(.A1(new_n405), .A2(new_n408), .B1(new_n379), .B2(new_n388), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT3), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n419), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(KEYINPUT4), .B1(new_n284), .B2(new_n397), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT4), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n425), .A2(new_n430), .A3(new_n415), .A4(new_n402), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(KEYINPUT79), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n433), .A3(KEYINPUT4), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n428), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n417), .A2(KEYINPUT81), .A3(new_n419), .A4(new_n420), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n423), .A2(KEYINPUT5), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT5), .B1(new_n429), .B2(new_n431), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n428), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XOR2_X1   g239(.A(G1gat), .B(G29gat), .Z(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G57gat), .B(G85gat), .ZN(new_n444));
  XNOR2_X1  g243(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n440), .A2(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n446), .B1(new_n438), .B2(new_n428), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n437), .A2(KEYINPUT83), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n447), .B1(new_n449), .B2(KEYINPUT6), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT6), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n445), .B1(new_n437), .B2(new_n439), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT83), .B1(new_n437), .B2(new_n448), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n451), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT37), .ZN(new_n456));
  NAND2_X1  g255(.A1(G226gat), .A2(G233gat), .ZN(new_n457));
  XOR2_X1   g256(.A(new_n457), .B(KEYINPUT75), .Z(new_n458));
  INV_X1    g257(.A(KEYINPUT29), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n458), .B1(new_n346), .B2(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(new_n457), .B1(new_n343), .B2(new_n305), .ZN(new_n461));
  OR2_X1    g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G197gat), .B(G204gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(G211gat), .A2(G218gat), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT22), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n463), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G211gat), .B(G218gat), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n467), .B(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n456), .B1(new_n462), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n470), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n346), .A2(new_n458), .ZN(new_n473));
  AOI21_X1  g272(.A(KEYINPUT29), .B1(new_n343), .B2(new_n305), .ZN(new_n474));
  INV_X1    g273(.A(new_n457), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n472), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT38), .B1(new_n471), .B2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(G64gat), .B(G92gat), .ZN(new_n479));
  XOR2_X1   g278(.A(new_n478), .B(new_n479), .Z(new_n480));
  OAI21_X1  g279(.A(new_n472), .B1(new_n460), .B2(new_n461), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n470), .B(new_n473), .C1(new_n474), .C2(new_n475), .ZN(new_n482));
  AND2_X1   g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n480), .B1(new_n483), .B2(new_n456), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n477), .A2(new_n484), .B1(new_n483), .B2(new_n480), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n480), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  NOR2_X1   g285(.A1(new_n480), .A2(new_n456), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n483), .A2(new_n456), .ZN(new_n489));
  OAI21_X1  g288(.A(KEYINPUT38), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n455), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G78gat), .B(G106gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(G22gat), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n470), .A2(new_n459), .A3(new_n397), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n397), .A2(KEYINPUT3), .ZN(new_n496));
  INV_X1    g295(.A(G228gat), .ZN(new_n497));
  INV_X1    g296(.A(G233gat), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n495), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n470), .B1(new_n427), .B2(new_n459), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT85), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n397), .A2(KEYINPUT3), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n472), .B1(new_n503), .B2(KEYINPUT29), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n496), .A2(new_n499), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT85), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .A4(new_n495), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n467), .A2(new_n469), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n468), .B1(new_n466), .B2(new_n463), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n459), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT84), .ZN(new_n512));
  AOI21_X1  g311(.A(KEYINPUT3), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n470), .A2(KEYINPUT84), .A3(new_n459), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n425), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI22_X1  g314(.A1(new_n515), .A2(new_n501), .B1(new_n497), .B2(new_n498), .ZN(new_n516));
  XOR2_X1   g315(.A(KEYINPUT31), .B(G50gat), .Z(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n508), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n508), .B2(new_n516), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n494), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(new_n521), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n523), .A2(new_n493), .A3(new_n519), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n429), .A2(new_n431), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n424), .A2(new_n427), .ZN(new_n527));
  AOI21_X1  g326(.A(new_n418), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n419), .B1(new_n417), .B2(new_n420), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT39), .ZN(new_n530));
  OR3_X1    g329(.A1(new_n528), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n446), .B1(new_n528), .B2(new_n530), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n533), .B1(KEYINPUT86), .B2(KEYINPUT40), .ZN(new_n534));
  NOR2_X1   g333(.A1(KEYINPUT86), .A2(KEYINPUT40), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n531), .A2(new_n535), .A3(new_n532), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n452), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT30), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n481), .A2(new_n482), .A3(new_n480), .ZN(new_n539));
  AOI21_X1  g338(.A(new_n486), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n481), .A2(new_n482), .A3(KEYINPUT30), .A4(new_n480), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT76), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n541), .A2(new_n542), .ZN(new_n544));
  OAI21_X1  g343(.A(new_n540), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n537), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n491), .A2(new_n525), .A3(new_n546), .ZN(new_n547));
  OR2_X1    g346(.A1(new_n541), .A2(new_n542), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n541), .A2(new_n542), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g349(.A1(new_n550), .A2(new_n450), .A3(new_n454), .A4(new_n540), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n522), .A2(new_n524), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  AND4_X1   g352(.A1(new_n370), .A2(new_n377), .A3(new_n547), .A4(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n455), .A2(new_n545), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT35), .B1(new_n556), .B2(KEYINPUT87), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n525), .B1(new_n361), .B2(new_n366), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(new_n369), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT87), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n560), .B1(new_n455), .B2(new_n545), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n552), .B1(new_n375), .B2(new_n368), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n563), .A2(new_n373), .A3(new_n556), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(KEYINPUT35), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n263), .B1(new_n555), .B2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G190gat), .B(G218gat), .Z(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT7), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(G85gat), .A3(G92gat), .A4(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  OAI211_X1 g374(.A(new_n569), .B(new_n570), .C1(new_n574), .C2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G99gat), .A2(G106gat), .ZN(new_n577));
  AOI22_X1  g376(.A1(KEYINPUT8), .A2(new_n577), .B1(new_n574), .B2(new_n575), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  XNOR2_X1  g378(.A(G99gat), .B(G106gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  XNOR2_X1  g380(.A(new_n579), .B(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n582), .B1(new_n233), .B2(new_n234), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  AND2_X1   g383(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT96), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NOR3_X1   g386(.A1(new_n583), .A2(KEYINPUT96), .A3(new_n585), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n582), .B1(new_n245), .B2(new_n247), .ZN(new_n589));
  OAI22_X1  g388(.A1(new_n587), .A2(new_n588), .B1(new_n589), .B2(KEYINPUT95), .ZN(new_n590));
  XNOR2_X1  g389(.A(new_n579), .B(new_n580), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n235), .A2(new_n246), .ZN(new_n592));
  INV_X1    g391(.A(new_n247), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n591), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT95), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n568), .B1(new_n590), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n598));
  XNOR2_X1  g397(.A(G134gat), .B(G162gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(new_n588), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n586), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n594), .A2(new_n595), .ZN(new_n603));
  INV_X1    g402(.A(new_n568), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n589), .A2(KEYINPUT95), .ZN(new_n605));
  NAND4_X1  g404(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n597), .A2(new_n600), .A3(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n600), .B1(new_n597), .B2(new_n606), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  XOR2_X1   g409(.A(G71gat), .B(G78gat), .Z(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT9), .ZN(new_n613));
  INV_X1    g412(.A(G71gat), .ZN(new_n614));
  INV_X1    g413(.A(G78gat), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n613), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  XOR2_X1   g415(.A(G57gat), .B(G64gat), .Z(new_n617));
  NAND3_X1  g416(.A1(new_n612), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n616), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(new_n611), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n622), .A2(KEYINPUT21), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n253), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT93), .B(KEYINPUT19), .ZN(new_n626));
  OR2_X1    g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OAI211_X1 g428(.A(G231gat), .B(G233gat), .C1(new_n622), .C2(KEYINPUT21), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT21), .ZN(new_n631));
  INV_X1    g430(.A(G231gat), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n621), .B(new_n631), .C1(new_n632), .C2(new_n498), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G127gat), .B(G155gat), .ZN(new_n635));
  XOR2_X1   g434(.A(new_n635), .B(KEYINPUT20), .Z(new_n636));
  OR2_X1    g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n634), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G183gat), .B(G211gat), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n637), .A2(new_n642), .A3(new_n638), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n627), .A2(new_n628), .A3(new_n641), .A4(new_n643), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G230gat), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n648), .A2(new_n498), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT97), .ZN(new_n650));
  OAI211_X1 g449(.A(new_n591), .B(new_n622), .C1(new_n650), .C2(new_n580), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n580), .A2(new_n650), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n582), .B1(new_n621), .B2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT10), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n651), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n591), .A2(new_n622), .A3(KEYINPUT10), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n649), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n651), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n649), .ZN(new_n660));
  XNOR2_X1  g459(.A(G120gat), .B(G148gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(G176gat), .B(G204gat), .ZN(new_n662));
  XOR2_X1   g461(.A(new_n661), .B(new_n662), .Z(new_n663));
  NAND3_X1  g462(.A1(new_n658), .A2(new_n660), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n658), .B2(new_n660), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n610), .A2(new_n647), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n567), .A2(new_n669), .ZN(new_n670));
  AND2_X1   g469(.A1(new_n450), .A2(new_n454), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT98), .B(G1gat), .Z(new_n673));
  XNOR2_X1  g472(.A(new_n672), .B(new_n673), .ZN(G1324gat));
  AND2_X1   g473(.A1(new_n567), .A2(new_n669), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n545), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n676), .A2(KEYINPUT99), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(KEYINPUT99), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n677), .A2(G8gat), .A3(new_n678), .ZN(new_n679));
  XOR2_X1   g478(.A(KEYINPUT16), .B(G8gat), .Z(new_n680));
  NAND4_X1  g479(.A1(new_n675), .A2(KEYINPUT42), .A3(new_n545), .A4(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n680), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n682), .B1(new_n677), .B2(new_n678), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n679), .B(new_n681), .C1(new_n683), .C2(KEYINPUT42), .ZN(G1325gat));
  AND2_X1   g483(.A1(new_n377), .A2(new_n370), .ZN(new_n685));
  OAI21_X1  g484(.A(G15gat), .B1(new_n670), .B2(new_n685), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n367), .A2(new_n369), .ZN(new_n687));
  INV_X1    g486(.A(new_n647), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n597), .A2(new_n606), .ZN(new_n689));
  INV_X1    g488(.A(new_n600), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n607), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n688), .A2(new_n692), .A3(new_n667), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(G15gat), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n567), .A2(new_n687), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n686), .A2(new_n695), .ZN(G1326gat));
  OR3_X1    g495(.A1(new_n670), .A2(KEYINPUT100), .A3(new_n525), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT100), .B1(new_n670), .B2(new_n525), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT43), .B(G22gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  INV_X1    g500(.A(KEYINPUT35), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n551), .B2(new_n560), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n539), .A2(new_n538), .ZN(new_n704));
  INV_X1    g503(.A(new_n486), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n706), .B1(new_n549), .B2(new_n548), .ZN(new_n707));
  AOI21_X1  g506(.A(KEYINPUT87), .B1(new_n671), .B2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n709), .A2(new_n559), .B1(KEYINPUT35), .B2(new_n564), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n610), .B1(new_n710), .B2(new_n554), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n647), .A2(new_n667), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n711), .A2(new_n263), .A3(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(G29gat), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n713), .A2(new_n714), .A3(new_n455), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT45), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n562), .A2(new_n717), .A3(new_n565), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n717), .B1(new_n562), .B2(new_n565), .ZN(new_n719));
  OAI21_X1  g518(.A(new_n555), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n721));
  NOR3_X1   g520(.A1(new_n608), .A2(new_n609), .A3(new_n721), .ZN(new_n722));
  AOI21_X1  g521(.A(KEYINPUT102), .B1(new_n691), .B2(new_n607), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n724), .A2(KEYINPUT44), .ZN(new_n725));
  AOI22_X1  g524(.A1(new_n720), .A2(new_n725), .B1(KEYINPUT44), .B2(new_n711), .ZN(new_n726));
  NOR4_X1   g525(.A1(new_n726), .A2(new_n671), .A3(new_n263), .A4(new_n712), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n716), .B1(new_n714), .B2(new_n727), .ZN(G1328gat));
  NOR2_X1   g527(.A1(new_n707), .A2(new_n223), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n713), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g529(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n731));
  OR2_X1    g530(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n731), .B2(new_n730), .ZN(new_n734));
  INV_X1    g533(.A(new_n726), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n263), .A2(new_n712), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n735), .A2(new_n545), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n223), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n737), .A2(KEYINPUT104), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(G1329gat));
  NOR3_X1   g540(.A1(new_n712), .A2(new_n692), .A3(G43gat), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n567), .A2(new_n687), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n743), .B1(new_n744), .B2(KEYINPUT47), .ZN(new_n745));
  INV_X1    g544(.A(new_n685), .ZN(new_n746));
  AND2_X1   g545(.A1(new_n720), .A2(new_n725), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n711), .A2(KEYINPUT44), .ZN(new_n748));
  OAI211_X1 g547(.A(new_n746), .B(new_n736), .C1(new_n747), .C2(new_n748), .ZN(new_n749));
  AOI21_X1  g548(.A(new_n745), .B1(new_n749), .B2(G43gat), .ZN(new_n750));
  AND2_X1   g549(.A1(new_n744), .A2(KEYINPUT47), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1330gat));
  INV_X1    g551(.A(new_n711), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n525), .A2(G50gat), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n753), .A2(new_n736), .A3(new_n754), .ZN(new_n755));
  OAI21_X1  g554(.A(new_n755), .B1(KEYINPUT106), .B2(KEYINPUT48), .ZN(new_n756));
  OAI211_X1 g555(.A(new_n552), .B(new_n736), .C1(new_n747), .C2(new_n748), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n756), .B1(new_n757), .B2(G50gat), .ZN(new_n758));
  AND2_X1   g557(.A1(KEYINPUT106), .A2(KEYINPUT48), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1331gat));
  NAND3_X1  g559(.A1(new_n671), .A2(KEYINPUT87), .A3(new_n707), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n702), .A3(new_n561), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n563), .A2(new_n373), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n702), .B1(new_n559), .B2(new_n556), .ZN(new_n765));
  OAI21_X1  g564(.A(KEYINPUT101), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n562), .A2(new_n717), .A3(new_n565), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n554), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n263), .A2(new_n688), .A3(new_n692), .A4(new_n668), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n455), .B(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g573(.A1(new_n770), .A2(new_n545), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n775), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n776));
  XOR2_X1   g575(.A(KEYINPUT49), .B(G64gat), .Z(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n775), .B2(new_n777), .ZN(G1333gat));
  AOI21_X1  g577(.A(new_n614), .B1(new_n770), .B2(new_n746), .ZN(new_n779));
  INV_X1    g578(.A(new_n687), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(G71gat), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n779), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  XNOR2_X1  g581(.A(new_n782), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g582(.A1(new_n770), .A2(new_n552), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g584(.A1(new_n263), .A2(new_n647), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n667), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n735), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(G85gat), .B1(new_n788), .B2(new_n671), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT51), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n263), .A2(new_n647), .A3(new_n610), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n790), .B1(new_n768), .B2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(new_n791), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n720), .A2(KEYINPUT51), .A3(new_n793), .ZN(new_n794));
  AND2_X1   g593(.A1(new_n792), .A2(new_n794), .ZN(new_n795));
  NAND3_X1  g594(.A1(new_n455), .A2(new_n668), .A3(new_n574), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n789), .B1(new_n795), .B2(new_n796), .ZN(G1336gat));
  INV_X1    g596(.A(new_n787), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n726), .A2(new_n707), .A3(new_n798), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n668), .A2(new_n545), .A3(new_n575), .ZN(new_n800));
  XOR2_X1   g599(.A(new_n800), .B(KEYINPUT108), .Z(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n792), .B2(new_n794), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT109), .ZN(new_n803));
  OAI22_X1  g602(.A1(new_n799), .A2(new_n575), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT52), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n545), .B(new_n787), .C1(new_n747), .C2(new_n748), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT52), .B1(new_n807), .B2(G92gat), .ZN(new_n808));
  OAI21_X1  g607(.A(KEYINPUT110), .B1(new_n795), .B2(new_n801), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n802), .A2(new_n810), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n808), .A2(new_n809), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n806), .A2(new_n812), .ZN(G1337gat));
  OAI21_X1  g612(.A(G99gat), .B1(new_n788), .B2(new_n685), .ZN(new_n814));
  OR3_X1    g613(.A1(new_n780), .A2(G99gat), .A3(new_n667), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n814), .B1(new_n795), .B2(new_n815), .ZN(G1338gat));
  OAI211_X1 g615(.A(new_n552), .B(new_n787), .C1(new_n747), .C2(new_n748), .ZN(new_n817));
  XNOR2_X1  g616(.A(KEYINPUT111), .B(G106gat), .ZN(new_n818));
  INV_X1    g617(.A(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n525), .A2(G106gat), .A3(new_n667), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n795), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT53), .B1(new_n820), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n817), .A2(new_n819), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n824), .B(new_n825), .C1(new_n795), .C2(new_n821), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n823), .A2(new_n826), .ZN(G1339gat));
  XNOR2_X1  g626(.A(new_n455), .B(KEYINPUT107), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n655), .A2(new_n649), .A3(new_n656), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n658), .A2(KEYINPUT54), .A3(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT54), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n663), .B1(new_n657), .B2(new_n831), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n830), .A2(KEYINPUT55), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT113), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n830), .A2(new_n832), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT55), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n834), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI211_X1 g636(.A(KEYINPUT113), .B(KEYINPUT55), .C1(new_n830), .C2(new_n832), .ZN(new_n838));
  OAI211_X1 g637(.A(new_n664), .B(new_n833), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT114), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n255), .A2(new_n208), .ZN(new_n842));
  AOI21_X1  g641(.A(new_n207), .B1(new_n244), .B2(new_n248), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n205), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  AND3_X1   g643(.A1(new_n262), .A2(new_n841), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n841), .B1(new_n262), .B2(new_n844), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n840), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n724), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n722), .A2(new_n723), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n252), .A2(new_n262), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n840), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n262), .A2(new_n668), .A3(new_n844), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n849), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n647), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT112), .B1(new_n669), .B2(new_n263), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n693), .A2(new_n850), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n828), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n559), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n860), .A2(new_n545), .ZN(new_n861));
  AOI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n850), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n839), .B1(new_n252), .B2(new_n262), .ZN(new_n863));
  INV_X1    g662(.A(new_n852), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n724), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI211_X1 g664(.A(new_n849), .B(new_n840), .C1(new_n846), .C2(new_n845), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n688), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n855), .A2(new_n857), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n525), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  OR4_X1    g668(.A1(new_n671), .A2(new_n869), .A3(new_n545), .A4(new_n780), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n870), .A2(new_n272), .A3(new_n263), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n862), .A2(new_n871), .ZN(G1340gat));
  AOI21_X1  g671(.A(G120gat), .B1(new_n861), .B2(new_n668), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n870), .A2(new_n274), .A3(new_n667), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n873), .A2(new_n874), .ZN(G1341gat));
  OAI21_X1  g674(.A(G127gat), .B1(new_n870), .B2(new_n647), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n278), .A3(new_n688), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1342gat));
  NOR2_X1   g677(.A1(new_n692), .A2(new_n545), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT115), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n860), .A2(new_n412), .A3(new_n413), .A4(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n882));
  OR2_X1    g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G134gat), .B1(new_n870), .B2(new_n692), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n881), .A2(new_n882), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n883), .A2(new_n884), .A3(new_n885), .ZN(G1343gat));
  NOR2_X1   g685(.A1(new_n746), .A2(new_n525), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n859), .A2(new_n707), .A3(new_n850), .A4(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  AOI22_X1  g688(.A1(new_n888), .A2(new_n380), .B1(KEYINPUT117), .B2(new_n889), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n552), .B1(new_n867), .B2(new_n868), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n835), .A2(new_n836), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n664), .A3(new_n833), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n894), .B1(new_n252), .B2(new_n262), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n692), .B1(new_n895), .B2(new_n864), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n688), .B1(new_n866), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n552), .B1(new_n897), .B2(new_n868), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(KEYINPUT57), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n746), .A2(new_n671), .A3(new_n545), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n263), .A2(new_n380), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n892), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n890), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n889), .A2(KEYINPUT117), .ZN(new_n904));
  INV_X1    g703(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n903), .B(new_n905), .ZN(G1344gat));
  NAND2_X1  g705(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n669), .A2(new_n263), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT118), .ZN(new_n909));
  OAI211_X1 g708(.A(new_n610), .B(new_n840), .C1(new_n845), .C2(new_n846), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n896), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n647), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n909), .A2(new_n912), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n525), .A2(KEYINPUT57), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n900), .A2(new_n668), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n907), .A2(new_n915), .A3(KEYINPUT119), .A4(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G148gat), .ZN(new_n918));
  AOI22_X1  g717(.A1(new_n891), .A2(KEYINPUT57), .B1(new_n913), .B2(new_n914), .ZN(new_n919));
  AOI21_X1  g718(.A(KEYINPUT119), .B1(new_n919), .B2(new_n916), .ZN(new_n920));
  OAI21_X1  g719(.A(KEYINPUT59), .B1(new_n918), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g720(.A1(new_n381), .A2(KEYINPUT59), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n892), .A2(new_n899), .A3(new_n900), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(new_n667), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n921), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n854), .A2(new_n858), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n772), .A3(new_n887), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n928), .A2(new_n381), .A3(new_n707), .A4(new_n668), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n925), .A2(new_n929), .ZN(G1345gat));
  NOR3_X1   g729(.A1(new_n923), .A2(new_n403), .A3(new_n647), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n927), .A2(new_n545), .A3(new_n647), .ZN(new_n932));
  XNOR2_X1  g731(.A(new_n932), .B(KEYINPUT120), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n931), .B1(new_n933), .B2(new_n403), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n923), .B2(new_n724), .ZN(new_n935));
  OR2_X1    g734(.A1(new_n880), .A2(G162gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n927), .B2(new_n936), .ZN(G1347gat));
  AOI21_X1  g736(.A(new_n455), .B1(new_n854), .B2(new_n858), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n763), .A2(new_n707), .ZN(new_n939));
  AND4_X1   g738(.A1(new_n286), .A2(new_n938), .A3(new_n850), .A4(new_n939), .ZN(new_n940));
  XOR2_X1   g739(.A(new_n940), .B(KEYINPUT121), .Z(new_n941));
  INV_X1    g740(.A(KEYINPUT122), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n828), .A2(new_n545), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n942), .B1(new_n943), .B2(new_n780), .ZN(new_n944));
  NAND4_X1  g743(.A1(new_n828), .A2(KEYINPUT122), .A3(new_n687), .A4(new_n545), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g745(.A(KEYINPUT123), .B1(new_n869), .B2(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT123), .ZN(new_n948));
  INV_X1    g747(.A(new_n946), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n926), .A2(new_n948), .A3(new_n525), .A4(new_n949), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n947), .A2(new_n950), .A3(new_n850), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n941), .B1(new_n286), .B2(new_n951), .ZN(G1348gat));
  AND3_X1   g751(.A1(new_n947), .A2(new_n950), .A3(new_n668), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n938), .A2(new_n939), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n668), .A2(new_n287), .ZN(new_n955));
  OAI22_X1  g754(.A1(new_n953), .A2(new_n287), .B1(new_n954), .B2(new_n955), .ZN(G1349gat));
  NAND3_X1  g755(.A1(new_n947), .A2(new_n950), .A3(new_n688), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G183gat), .ZN(new_n958));
  NAND4_X1  g757(.A1(new_n938), .A2(new_n300), .A3(new_n688), .A4(new_n939), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(KEYINPUT124), .B(KEYINPUT60), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n958), .A2(new_n959), .A3(new_n961), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(G1350gat));
  NAND3_X1  g764(.A1(new_n947), .A2(new_n950), .A3(new_n610), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G190gat), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT125), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n966), .A2(KEYINPUT125), .A3(G190gat), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(KEYINPUT61), .A3(new_n970), .ZN(new_n971));
  AND4_X1   g770(.A1(new_n299), .A2(new_n938), .A3(new_n849), .A4(new_n939), .ZN(new_n972));
  AOI21_X1  g771(.A(KEYINPUT125), .B1(new_n966), .B2(G190gat), .ZN(new_n973));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n974));
  AOI21_X1  g773(.A(new_n972), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n971), .A2(new_n975), .ZN(G1351gat));
  NOR2_X1   g775(.A1(new_n746), .A2(new_n943), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n919), .A2(G197gat), .A3(new_n850), .A4(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(G197gat), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n746), .A2(new_n707), .A3(new_n525), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n938), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n979), .B1(new_n981), .B2(new_n263), .ZN(new_n982));
  AND2_X1   g781(.A1(new_n978), .A2(new_n982), .ZN(G1352gat));
  XOR2_X1   g782(.A(KEYINPUT126), .B(G204gat), .Z(new_n984));
  INV_X1    g783(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n919), .A2(new_n977), .ZN(new_n986));
  OAI21_X1  g785(.A(new_n985), .B1(new_n986), .B2(new_n667), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n667), .A2(new_n985), .ZN(new_n988));
  INV_X1    g787(.A(new_n988), .ZN(new_n989));
  OAI21_X1  g788(.A(KEYINPUT62), .B1(new_n981), .B2(new_n989), .ZN(new_n990));
  OR3_X1    g789(.A1(new_n981), .A2(KEYINPUT62), .A3(new_n989), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n987), .A2(new_n990), .A3(new_n991), .ZN(G1353gat));
  OR3_X1    g791(.A1(new_n981), .A2(G211gat), .A3(new_n647), .ZN(new_n993));
  NAND3_X1  g792(.A1(new_n919), .A2(new_n688), .A3(new_n977), .ZN(new_n994));
  AND4_X1   g793(.A1(KEYINPUT127), .A2(new_n994), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n995));
  OAI21_X1  g794(.A(G211gat), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n996));
  INV_X1    g795(.A(new_n996), .ZN(new_n997));
  AOI22_X1  g796(.A1(new_n994), .A2(new_n997), .B1(KEYINPUT127), .B2(KEYINPUT63), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n993), .B1(new_n995), .B2(new_n998), .ZN(G1354gat));
  OAI21_X1  g798(.A(G218gat), .B1(new_n986), .B2(new_n692), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n724), .A2(G218gat), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1000), .B1(new_n981), .B2(new_n1001), .ZN(G1355gat));
endmodule


