

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n742), .A2(n741), .ZN(n744) );
  BUF_X1 U553 ( .A(n688), .Z(n566) );
  AND2_X2 U554 ( .A1(n521), .A2(G2104), .ZN(n892) );
  NOR2_X2 U555 ( .A1(n530), .A2(n529), .ZN(G160) );
  XNOR2_X1 U556 ( .A(n744), .B(n743), .ZN(n752) );
  NOR2_X2 U557 ( .A1(G2104), .A2(n521), .ZN(n567) );
  XOR2_X1 U558 ( .A(n734), .B(n733), .Z(n517) );
  XOR2_X1 U559 ( .A(n771), .B(KEYINPUT97), .Z(n518) );
  OR2_X1 U560 ( .A1(n778), .A2(n777), .ZN(n519) );
  OR2_X1 U561 ( .A1(n725), .A2(n724), .ZN(n520) );
  NOR2_X1 U562 ( .A1(n735), .A2(n950), .ZN(n696) );
  AND2_X1 U563 ( .A1(n700), .A2(n699), .ZN(n703) );
  INV_X1 U564 ( .A(KEYINPUT92), .ZN(n701) );
  XNOR2_X1 U565 ( .A(KEYINPUT94), .B(KEYINPUT32), .ZN(n743) );
  NAND2_X1 U566 ( .A1(n779), .A2(n519), .ZN(n780) );
  OR2_X1 U567 ( .A1(n518), .A2(n780), .ZN(n796) );
  XNOR2_X1 U568 ( .A(n578), .B(KEYINPUT13), .ZN(n579) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n527) );
  XNOR2_X1 U570 ( .A(n580), .B(n579), .ZN(n583) );
  NOR2_X1 U571 ( .A1(G651), .A2(n658), .ZN(n653) );
  NAND2_X1 U572 ( .A1(n585), .A2(n584), .ZN(n970) );
  INV_X1 U573 ( .A(G2105), .ZN(n521) );
  NAND2_X1 U574 ( .A1(n567), .A2(G125), .ZN(n526) );
  AND2_X1 U575 ( .A1(G2105), .A2(G2104), .ZN(n786) );
  NAND2_X1 U576 ( .A1(n786), .A2(G113), .ZN(n524) );
  NAND2_X1 U577 ( .A1(G101), .A2(n892), .ZN(n522) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n522), .Z(n523) );
  AND2_X1 U579 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U580 ( .A1(n526), .A2(n525), .ZN(n530) );
  XOR2_X1 U581 ( .A(n527), .B(KEYINPUT17), .Z(n528) );
  XNOR2_X1 U582 ( .A(n528), .B(KEYINPUT66), .ZN(n688) );
  AND2_X1 U583 ( .A1(G137), .A2(n688), .ZN(n529) );
  XOR2_X1 U584 ( .A(G2446), .B(G2430), .Z(n532) );
  XNOR2_X1 U585 ( .A(G2451), .B(G2454), .ZN(n531) );
  XNOR2_X1 U586 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U587 ( .A(n533), .B(G2427), .Z(n535) );
  XNOR2_X1 U588 ( .A(G1348), .B(G1341), .ZN(n534) );
  XNOR2_X1 U589 ( .A(n535), .B(n534), .ZN(n539) );
  XOR2_X1 U590 ( .A(G2443), .B(KEYINPUT100), .Z(n537) );
  XNOR2_X1 U591 ( .A(G2438), .B(G2435), .ZN(n536) );
  XNOR2_X1 U592 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U593 ( .A(n539), .B(n538), .Z(n540) );
  AND2_X1 U594 ( .A1(G14), .A2(n540), .ZN(G401) );
  AND2_X1 U595 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U596 ( .A(G57), .ZN(G237) );
  INV_X1 U597 ( .A(G69), .ZN(G235) );
  INV_X1 U598 ( .A(G108), .ZN(G238) );
  INV_X1 U599 ( .A(G120), .ZN(G236) );
  INV_X1 U600 ( .A(G132), .ZN(G219) );
  XOR2_X1 U601 ( .A(G543), .B(KEYINPUT0), .Z(n658) );
  NAND2_X1 U602 ( .A1(G52), .A2(n653), .ZN(n541) );
  XOR2_X1 U603 ( .A(KEYINPUT68), .B(n541), .Z(n551) );
  NOR2_X1 U604 ( .A1(G651), .A2(G543), .ZN(n542) );
  XOR2_X2 U605 ( .A(KEYINPUT65), .B(n542), .Z(n645) );
  NAND2_X1 U606 ( .A1(G90), .A2(n645), .ZN(n544) );
  INV_X1 U607 ( .A(G651), .ZN(n546) );
  NOR2_X1 U608 ( .A1(n658), .A2(n546), .ZN(n643) );
  NAND2_X1 U609 ( .A1(G77), .A2(n643), .ZN(n543) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  XNOR2_X1 U611 ( .A(n545), .B(KEYINPUT9), .ZN(n549) );
  NOR2_X1 U612 ( .A1(G543), .A2(n546), .ZN(n547) );
  XOR2_X1 U613 ( .A(KEYINPUT1), .B(n547), .Z(n657) );
  NAND2_X1 U614 ( .A1(G64), .A2(n657), .ZN(n548) );
  NAND2_X1 U615 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U616 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U617 ( .A1(n653), .A2(G51), .ZN(n552) );
  XOR2_X1 U618 ( .A(KEYINPUT73), .B(n552), .Z(n554) );
  NAND2_X1 U619 ( .A1(n657), .A2(G63), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT6), .B(n555), .ZN(n562) );
  NAND2_X1 U622 ( .A1(G89), .A2(n645), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT4), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n557), .B(KEYINPUT72), .ZN(n559) );
  NAND2_X1 U625 ( .A1(G76), .A2(n643), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U627 ( .A(n560), .B(KEYINPUT5), .Z(n561) );
  NOR2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U629 ( .A(KEYINPUT74), .B(n563), .Z(n564) );
  XNOR2_X1 U630 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  XNOR2_X1 U631 ( .A(KEYINPUT75), .B(KEYINPUT8), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G168), .ZN(G286) );
  AND2_X1 U633 ( .A1(G138), .A2(n566), .ZN(n572) );
  NAND2_X1 U634 ( .A1(G102), .A2(n892), .ZN(n571) );
  NAND2_X1 U635 ( .A1(G114), .A2(n786), .ZN(n569) );
  NAND2_X1 U636 ( .A1(G126), .A2(n567), .ZN(n568) );
  AND2_X1 U637 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n689) );
  NOR2_X1 U639 ( .A1(n572), .A2(n689), .ZN(G164) );
  NAND2_X1 U640 ( .A1(G7), .A2(G661), .ZN(n573) );
  XNOR2_X1 U641 ( .A(n573), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U642 ( .A(G223), .ZN(n835) );
  NAND2_X1 U643 ( .A1(n835), .A2(G567), .ZN(n574) );
  XOR2_X1 U644 ( .A(KEYINPUT11), .B(n574), .Z(G234) );
  NAND2_X1 U645 ( .A1(n645), .A2(G81), .ZN(n575) );
  XNOR2_X1 U646 ( .A(n575), .B(KEYINPUT12), .ZN(n577) );
  NAND2_X1 U647 ( .A1(G68), .A2(n643), .ZN(n576) );
  NAND2_X1 U648 ( .A1(n577), .A2(n576), .ZN(n580) );
  XNOR2_X1 U649 ( .A(KEYINPUT70), .B(KEYINPUT71), .ZN(n578) );
  NAND2_X1 U650 ( .A1(n657), .A2(G56), .ZN(n581) );
  XOR2_X1 U651 ( .A(KEYINPUT14), .B(n581), .Z(n582) );
  NOR2_X1 U652 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U653 ( .A1(n653), .A2(G43), .ZN(n584) );
  INV_X1 U654 ( .A(G860), .ZN(n626) );
  OR2_X1 U655 ( .A1(n970), .A2(n626), .ZN(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G92), .A2(n645), .ZN(n587) );
  NAND2_X1 U659 ( .A1(G79), .A2(n643), .ZN(n586) );
  NAND2_X1 U660 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U661 ( .A1(G66), .A2(n657), .ZN(n589) );
  NAND2_X1 U662 ( .A1(G54), .A2(n653), .ZN(n588) );
  NAND2_X1 U663 ( .A1(n589), .A2(n588), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U665 ( .A(KEYINPUT15), .B(n592), .Z(n976) );
  OR2_X1 U666 ( .A1(n976), .A2(G868), .ZN(n593) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U668 ( .A1(G65), .A2(n657), .ZN(n596) );
  NAND2_X1 U669 ( .A1(G53), .A2(n653), .ZN(n595) );
  NAND2_X1 U670 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U671 ( .A1(G91), .A2(n645), .ZN(n598) );
  NAND2_X1 U672 ( .A1(G78), .A2(n643), .ZN(n597) );
  NAND2_X1 U673 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U674 ( .A1(n600), .A2(n599), .ZN(n980) );
  INV_X1 U675 ( .A(n980), .ZN(G299) );
  XOR2_X1 U676 ( .A(KEYINPUT76), .B(G868), .Z(n601) );
  NOR2_X1 U677 ( .A1(G286), .A2(n601), .ZN(n603) );
  NOR2_X1 U678 ( .A1(G868), .A2(G299), .ZN(n602) );
  NOR2_X1 U679 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U680 ( .A1(n626), .A2(G559), .ZN(n604) );
  NAND2_X1 U681 ( .A1(n604), .A2(n976), .ZN(n605) );
  XNOR2_X1 U682 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U683 ( .A1(G868), .A2(n970), .ZN(n608) );
  NAND2_X1 U684 ( .A1(G868), .A2(n976), .ZN(n606) );
  NOR2_X1 U685 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U686 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U687 ( .A1(G123), .A2(n567), .ZN(n609) );
  XNOR2_X1 U688 ( .A(n609), .B(KEYINPUT18), .ZN(n612) );
  NAND2_X1 U689 ( .A1(G111), .A2(n786), .ZN(n610) );
  XOR2_X1 U690 ( .A(KEYINPUT77), .B(n610), .Z(n611) );
  NAND2_X1 U691 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G99), .A2(n892), .ZN(n614) );
  NAND2_X1 U693 ( .A1(G135), .A2(n566), .ZN(n613) );
  NAND2_X1 U694 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U695 ( .A1(n616), .A2(n615), .ZN(n921) );
  XNOR2_X1 U696 ( .A(G2096), .B(n921), .ZN(n618) );
  INV_X1 U697 ( .A(G2100), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(G156) );
  NAND2_X1 U699 ( .A1(G93), .A2(n645), .ZN(n620) );
  NAND2_X1 U700 ( .A1(G80), .A2(n643), .ZN(n619) );
  NAND2_X1 U701 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U702 ( .A1(G67), .A2(n657), .ZN(n622) );
  NAND2_X1 U703 ( .A1(G55), .A2(n653), .ZN(n621) );
  NAND2_X1 U704 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U705 ( .A1(n624), .A2(n623), .ZN(n669) );
  XOR2_X1 U706 ( .A(n669), .B(KEYINPUT78), .Z(n628) );
  NAND2_X1 U707 ( .A1(G559), .A2(n976), .ZN(n625) );
  XOR2_X1 U708 ( .A(n970), .B(n625), .Z(n667) );
  NAND2_X1 U709 ( .A1(n667), .A2(n626), .ZN(n627) );
  XNOR2_X1 U710 ( .A(n628), .B(n627), .ZN(G145) );
  NAND2_X1 U711 ( .A1(G88), .A2(n645), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G75), .A2(n643), .ZN(n629) );
  NAND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U714 ( .A1(n657), .A2(G62), .ZN(n631) );
  XOR2_X1 U715 ( .A(KEYINPUT80), .B(n631), .Z(n632) );
  NOR2_X1 U716 ( .A1(n633), .A2(n632), .ZN(n635) );
  NAND2_X1 U717 ( .A1(n653), .A2(G50), .ZN(n634) );
  NAND2_X1 U718 ( .A1(n635), .A2(n634), .ZN(G303) );
  INV_X1 U719 ( .A(G303), .ZN(G166) );
  NAND2_X1 U720 ( .A1(G72), .A2(n643), .ZN(n637) );
  NAND2_X1 U721 ( .A1(G47), .A2(n653), .ZN(n636) );
  NAND2_X1 U722 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U723 ( .A1(G85), .A2(n645), .ZN(n638) );
  XNOR2_X1 U724 ( .A(KEYINPUT67), .B(n638), .ZN(n639) );
  NOR2_X1 U725 ( .A1(n640), .A2(n639), .ZN(n642) );
  NAND2_X1 U726 ( .A1(n657), .A2(G60), .ZN(n641) );
  NAND2_X1 U727 ( .A1(n642), .A2(n641), .ZN(G290) );
  NAND2_X1 U728 ( .A1(G73), .A2(n643), .ZN(n644) );
  XNOR2_X1 U729 ( .A(n644), .B(KEYINPUT2), .ZN(n652) );
  NAND2_X1 U730 ( .A1(G86), .A2(n645), .ZN(n647) );
  NAND2_X1 U731 ( .A1(G48), .A2(n653), .ZN(n646) );
  NAND2_X1 U732 ( .A1(n647), .A2(n646), .ZN(n650) );
  NAND2_X1 U733 ( .A1(G61), .A2(n657), .ZN(n648) );
  XNOR2_X1 U734 ( .A(KEYINPUT79), .B(n648), .ZN(n649) );
  NOR2_X1 U735 ( .A1(n650), .A2(n649), .ZN(n651) );
  NAND2_X1 U736 ( .A1(n652), .A2(n651), .ZN(G305) );
  NAND2_X1 U737 ( .A1(G49), .A2(n653), .ZN(n655) );
  NAND2_X1 U738 ( .A1(G74), .A2(G651), .ZN(n654) );
  NAND2_X1 U739 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U740 ( .A1(n657), .A2(n656), .ZN(n660) );
  NAND2_X1 U741 ( .A1(n658), .A2(G87), .ZN(n659) );
  NAND2_X1 U742 ( .A1(n660), .A2(n659), .ZN(G288) );
  XNOR2_X1 U743 ( .A(G166), .B(G290), .ZN(n661) );
  XNOR2_X1 U744 ( .A(n661), .B(G305), .ZN(n664) );
  XOR2_X1 U745 ( .A(KEYINPUT81), .B(KEYINPUT19), .Z(n662) );
  XNOR2_X1 U746 ( .A(G288), .B(n662), .ZN(n663) );
  XOR2_X1 U747 ( .A(n664), .B(n663), .Z(n666) );
  XNOR2_X1 U748 ( .A(n980), .B(n669), .ZN(n665) );
  XNOR2_X1 U749 ( .A(n666), .B(n665), .ZN(n905) );
  XNOR2_X1 U750 ( .A(n667), .B(n905), .ZN(n668) );
  NAND2_X1 U751 ( .A1(n668), .A2(G868), .ZN(n671) );
  OR2_X1 U752 ( .A1(G868), .A2(n669), .ZN(n670) );
  NAND2_X1 U753 ( .A1(n671), .A2(n670), .ZN(G295) );
  XOR2_X1 U754 ( .A(KEYINPUT20), .B(KEYINPUT82), .Z(n673) );
  NAND2_X1 U755 ( .A1(G2084), .A2(G2078), .ZN(n672) );
  XNOR2_X1 U756 ( .A(n673), .B(n672), .ZN(n674) );
  NAND2_X1 U757 ( .A1(G2090), .A2(n674), .ZN(n675) );
  XNOR2_X1 U758 ( .A(KEYINPUT21), .B(n675), .ZN(n676) );
  NAND2_X1 U759 ( .A1(n676), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U760 ( .A(KEYINPUT69), .B(G82), .ZN(G220) );
  XNOR2_X1 U761 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U762 ( .A1(G219), .A2(G220), .ZN(n678) );
  XNOR2_X1 U763 ( .A(KEYINPUT83), .B(KEYINPUT22), .ZN(n677) );
  XNOR2_X1 U764 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U765 ( .A1(n679), .A2(G218), .ZN(n680) );
  NAND2_X1 U766 ( .A1(G96), .A2(n680), .ZN(n841) );
  NAND2_X1 U767 ( .A1(n841), .A2(G2106), .ZN(n685) );
  NOR2_X1 U768 ( .A1(G236), .A2(G238), .ZN(n682) );
  NOR2_X1 U769 ( .A1(G235), .A2(G237), .ZN(n681) );
  NAND2_X1 U770 ( .A1(n682), .A2(n681), .ZN(n683) );
  XNOR2_X1 U771 ( .A(KEYINPUT84), .B(n683), .ZN(n842) );
  NAND2_X1 U772 ( .A1(n842), .A2(G567), .ZN(n684) );
  NAND2_X1 U773 ( .A1(n685), .A2(n684), .ZN(n843) );
  NAND2_X1 U774 ( .A1(G661), .A2(G483), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n843), .A2(n686), .ZN(n840) );
  NAND2_X1 U776 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U777 ( .A(G1384), .ZN(n690) );
  AND2_X1 U778 ( .A1(G138), .A2(n690), .ZN(n687) );
  NAND2_X1 U779 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U780 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U781 ( .A1(n692), .A2(n691), .ZN(n693) );
  XNOR2_X1 U782 ( .A(n693), .B(KEYINPUT64), .ZN(n781) );
  INV_X1 U783 ( .A(n781), .ZN(n694) );
  NAND2_X1 U784 ( .A1(G160), .A2(G40), .ZN(n782) );
  NOR2_X2 U785 ( .A1(n694), .A2(n782), .ZN(n721) );
  INV_X1 U786 ( .A(n721), .ZN(n735) );
  INV_X1 U787 ( .A(G1996), .ZN(n950) );
  INV_X1 U788 ( .A(KEYINPUT26), .ZN(n695) );
  XNOR2_X1 U789 ( .A(n696), .B(n695), .ZN(n698) );
  NAND2_X1 U790 ( .A1(n735), .A2(G1341), .ZN(n697) );
  AND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n700) );
  INV_X1 U792 ( .A(n970), .ZN(n699) );
  NOR2_X1 U793 ( .A1(n703), .A2(n976), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n702), .B(n701), .ZN(n709) );
  NAND2_X1 U795 ( .A1(n703), .A2(n976), .ZN(n707) );
  NOR2_X1 U796 ( .A1(n721), .A2(G1348), .ZN(n705) );
  NOR2_X1 U797 ( .A1(G2067), .A2(n735), .ZN(n704) );
  NOR2_X1 U798 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U799 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U800 ( .A1(n709), .A2(n708), .ZN(n715) );
  NAND2_X1 U801 ( .A1(n735), .A2(G1956), .ZN(n712) );
  NAND2_X1 U802 ( .A1(n721), .A2(G2072), .ZN(n710) );
  XOR2_X1 U803 ( .A(KEYINPUT27), .B(n710), .Z(n711) );
  NAND2_X1 U804 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U805 ( .A(n713), .B(KEYINPUT91), .ZN(n716) );
  NAND2_X1 U806 ( .A1(n980), .A2(n716), .ZN(n714) );
  NAND2_X1 U807 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U808 ( .A1(n980), .A2(n716), .ZN(n717) );
  XOR2_X1 U809 ( .A(n717), .B(KEYINPUT28), .Z(n718) );
  NAND2_X1 U810 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U811 ( .A(n720), .B(KEYINPUT29), .ZN(n725) );
  NAND2_X1 U812 ( .A1(G1961), .A2(n735), .ZN(n723) );
  XOR2_X1 U813 ( .A(KEYINPUT25), .B(G2078), .Z(n957) );
  NAND2_X1 U814 ( .A1(n721), .A2(n957), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n729) );
  NOR2_X1 U816 ( .A1(G301), .A2(n729), .ZN(n724) );
  INV_X1 U817 ( .A(KEYINPUT31), .ZN(n734) );
  NAND2_X1 U818 ( .A1(G8), .A2(n735), .ZN(n778) );
  NOR2_X1 U819 ( .A1(G1966), .A2(n778), .ZN(n748) );
  NOR2_X1 U820 ( .A1(G2084), .A2(n735), .ZN(n745) );
  NOR2_X1 U821 ( .A1(n748), .A2(n745), .ZN(n726) );
  NAND2_X1 U822 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U823 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U824 ( .A1(G168), .A2(n728), .ZN(n731) );
  AND2_X1 U825 ( .A1(G301), .A2(n729), .ZN(n730) );
  NOR2_X1 U826 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U827 ( .A(n732), .B(KEYINPUT93), .ZN(n733) );
  NAND2_X1 U828 ( .A1(n520), .A2(n517), .ZN(n746) );
  NAND2_X1 U829 ( .A1(n746), .A2(G286), .ZN(n742) );
  INV_X1 U830 ( .A(G8), .ZN(n740) );
  NOR2_X1 U831 ( .A1(G1971), .A2(n778), .ZN(n737) );
  NOR2_X1 U832 ( .A1(G2090), .A2(n735), .ZN(n736) );
  NOR2_X1 U833 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U834 ( .A1(n738), .A2(G303), .ZN(n739) );
  OR2_X1 U835 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U836 ( .A1(n745), .A2(G8), .ZN(n750) );
  INV_X1 U837 ( .A(n746), .ZN(n747) );
  NOR2_X1 U838 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n774) );
  NOR2_X1 U841 ( .A1(G1976), .A2(G288), .ZN(n753) );
  XNOR2_X1 U842 ( .A(KEYINPUT95), .B(n753), .ZN(n986) );
  NAND2_X1 U843 ( .A1(n774), .A2(n986), .ZN(n762) );
  NOR2_X1 U844 ( .A1(G1971), .A2(G303), .ZN(n760) );
  XNOR2_X1 U845 ( .A(G1981), .B(G305), .ZN(n972) );
  INV_X1 U846 ( .A(KEYINPUT33), .ZN(n756) );
  OR2_X1 U847 ( .A1(n778), .A2(n986), .ZN(n754) );
  NOR2_X1 U848 ( .A1(n756), .A2(n754), .ZN(n755) );
  XOR2_X1 U849 ( .A(n755), .B(KEYINPUT96), .Z(n763) );
  INV_X1 U850 ( .A(n763), .ZN(n757) );
  OR2_X1 U851 ( .A1(n757), .A2(n756), .ZN(n758) );
  OR2_X1 U852 ( .A1(n972), .A2(n758), .ZN(n768) );
  INV_X1 U853 ( .A(n768), .ZN(n759) );
  OR2_X1 U854 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n770) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n981) );
  AND2_X1 U857 ( .A1(n981), .A2(n763), .ZN(n765) );
  INV_X1 U858 ( .A(n972), .ZN(n764) );
  NAND2_X1 U859 ( .A1(n765), .A2(n764), .ZN(n766) );
  OR2_X1 U860 ( .A1(n766), .A2(n778), .ZN(n767) );
  AND2_X1 U861 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U862 ( .A1(n770), .A2(n769), .ZN(n771) );
  NOR2_X1 U863 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U864 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n775), .A2(n778), .ZN(n779) );
  NOR2_X1 U867 ( .A1(G1981), .A2(G305), .ZN(n776) );
  XOR2_X1 U868 ( .A(n776), .B(KEYINPUT24), .Z(n777) );
  NOR2_X1 U869 ( .A1(n781), .A2(n782), .ZN(n829) );
  NAND2_X1 U870 ( .A1(G104), .A2(n892), .ZN(n784) );
  NAND2_X1 U871 ( .A1(G140), .A2(n566), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U873 ( .A(KEYINPUT34), .B(n785), .ZN(n793) );
  XNOR2_X1 U874 ( .A(KEYINPUT86), .B(KEYINPUT35), .ZN(n791) );
  NAND2_X1 U875 ( .A1(n567), .A2(G128), .ZN(n789) );
  NAND2_X1 U876 ( .A1(n786), .A2(G116), .ZN(n787) );
  XOR2_X1 U877 ( .A(KEYINPUT85), .B(n787), .Z(n788) );
  NAND2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U879 ( .A(n791), .B(n790), .Z(n792) );
  NOR2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n794) );
  XOR2_X1 U881 ( .A(n794), .B(KEYINPUT36), .Z(n795) );
  XNOR2_X1 U882 ( .A(KEYINPUT87), .B(n795), .ZN(n900) );
  XNOR2_X1 U883 ( .A(G2067), .B(KEYINPUT37), .ZN(n819) );
  NOR2_X1 U884 ( .A1(n900), .A2(n819), .ZN(n926) );
  NAND2_X1 U885 ( .A1(n829), .A2(n926), .ZN(n826) );
  NAND2_X1 U886 ( .A1(n796), .A2(n826), .ZN(n816) );
  NAND2_X1 U887 ( .A1(G107), .A2(n786), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G119), .A2(n567), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n892), .A2(G95), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT88), .B(n799), .Z(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G131), .A2(n566), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n881) );
  AND2_X1 U895 ( .A1(n881), .A2(G1991), .ZN(n813) );
  NAND2_X1 U896 ( .A1(G105), .A2(n892), .ZN(n804) );
  XOR2_X1 U897 ( .A(KEYINPUT38), .B(n804), .Z(n809) );
  NAND2_X1 U898 ( .A1(G117), .A2(n786), .ZN(n806) );
  NAND2_X1 U899 ( .A1(G129), .A2(n567), .ZN(n805) );
  NAND2_X1 U900 ( .A1(n806), .A2(n805), .ZN(n807) );
  XOR2_X1 U901 ( .A(KEYINPUT89), .B(n807), .Z(n808) );
  NOR2_X1 U902 ( .A1(n809), .A2(n808), .ZN(n811) );
  NAND2_X1 U903 ( .A1(G141), .A2(n566), .ZN(n810) );
  NAND2_X1 U904 ( .A1(n811), .A2(n810), .ZN(n878) );
  AND2_X1 U905 ( .A1(n878), .A2(G1996), .ZN(n812) );
  NOR2_X1 U906 ( .A1(n813), .A2(n812), .ZN(n923) );
  INV_X1 U907 ( .A(n829), .ZN(n814) );
  NOR2_X1 U908 ( .A1(n923), .A2(n814), .ZN(n822) );
  XNOR2_X1 U909 ( .A(KEYINPUT90), .B(n822), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n816), .A2(n815), .ZN(n818) );
  XNOR2_X1 U911 ( .A(G1986), .B(G290), .ZN(n988) );
  NAND2_X1 U912 ( .A1(n988), .A2(n829), .ZN(n817) );
  NAND2_X1 U913 ( .A1(n818), .A2(n817), .ZN(n832) );
  NAND2_X1 U914 ( .A1(n900), .A2(n819), .ZN(n933) );
  NOR2_X1 U915 ( .A1(G1996), .A2(n878), .ZN(n918) );
  NOR2_X1 U916 ( .A1(G1991), .A2(n881), .ZN(n922) );
  NOR2_X1 U917 ( .A1(G1986), .A2(G290), .ZN(n820) );
  NOR2_X1 U918 ( .A1(n922), .A2(n820), .ZN(n821) );
  NOR2_X1 U919 ( .A1(n822), .A2(n821), .ZN(n823) );
  NOR2_X1 U920 ( .A1(n918), .A2(n823), .ZN(n824) );
  XNOR2_X1 U921 ( .A(KEYINPUT39), .B(n824), .ZN(n825) );
  XNOR2_X1 U922 ( .A(n825), .B(KEYINPUT98), .ZN(n827) );
  NAND2_X1 U923 ( .A1(n827), .A2(n826), .ZN(n828) );
  NAND2_X1 U924 ( .A1(n933), .A2(n828), .ZN(n830) );
  NAND2_X1 U925 ( .A1(n830), .A2(n829), .ZN(n831) );
  NAND2_X1 U926 ( .A1(n832), .A2(n831), .ZN(n834) );
  XOR2_X1 U927 ( .A(KEYINPUT99), .B(KEYINPUT40), .Z(n833) );
  XNOR2_X1 U928 ( .A(n834), .B(n833), .ZN(G329) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n835), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n836) );
  XNOR2_X1 U931 ( .A(KEYINPUT101), .B(n836), .ZN(n837) );
  NAND2_X1 U932 ( .A1(n837), .A2(G661), .ZN(n838) );
  XNOR2_X1 U933 ( .A(KEYINPUT102), .B(n838), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(G188) );
  INV_X1 U937 ( .A(G96), .ZN(G221) );
  NOR2_X1 U938 ( .A1(n842), .A2(n841), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n843), .ZN(G319) );
  XOR2_X1 U941 ( .A(KEYINPUT42), .B(G2072), .Z(n845) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2078), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U944 ( .A(n846), .B(G2096), .Z(n848) );
  XNOR2_X1 U945 ( .A(G2090), .B(G2084), .ZN(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U947 ( .A(KEYINPUT43), .B(G2678), .Z(n850) );
  XNOR2_X1 U948 ( .A(KEYINPUT103), .B(G2100), .ZN(n849) );
  XNOR2_X1 U949 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U950 ( .A(n852), .B(n851), .Z(G227) );
  XNOR2_X1 U951 ( .A(G1966), .B(KEYINPUT41), .ZN(n862) );
  XOR2_X1 U952 ( .A(G1981), .B(G1956), .Z(n854) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1961), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n858) );
  XOR2_X1 U955 ( .A(G1976), .B(G1971), .Z(n856) );
  XNOR2_X1 U956 ( .A(G1996), .B(G1991), .ZN(n855) );
  XNOR2_X1 U957 ( .A(n856), .B(n855), .ZN(n857) );
  XOR2_X1 U958 ( .A(n858), .B(n857), .Z(n860) );
  XNOR2_X1 U959 ( .A(KEYINPUT104), .B(G2474), .ZN(n859) );
  XNOR2_X1 U960 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U961 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U962 ( .A1(G100), .A2(n892), .ZN(n864) );
  NAND2_X1 U963 ( .A1(G112), .A2(n786), .ZN(n863) );
  NAND2_X1 U964 ( .A1(n864), .A2(n863), .ZN(n865) );
  XNOR2_X1 U965 ( .A(n865), .B(KEYINPUT105), .ZN(n867) );
  NAND2_X1 U966 ( .A1(G136), .A2(n566), .ZN(n866) );
  NAND2_X1 U967 ( .A1(n867), .A2(n866), .ZN(n870) );
  NAND2_X1 U968 ( .A1(n567), .A2(G124), .ZN(n868) );
  XOR2_X1 U969 ( .A(KEYINPUT44), .B(n868), .Z(n869) );
  NOR2_X1 U970 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G103), .A2(n892), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G139), .A2(n566), .ZN(n871) );
  NAND2_X1 U973 ( .A1(n872), .A2(n871), .ZN(n877) );
  NAND2_X1 U974 ( .A1(G115), .A2(n786), .ZN(n874) );
  NAND2_X1 U975 ( .A1(G127), .A2(n567), .ZN(n873) );
  NAND2_X1 U976 ( .A1(n874), .A2(n873), .ZN(n875) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n875), .Z(n876) );
  NOR2_X1 U978 ( .A1(n877), .A2(n876), .ZN(n937) );
  XOR2_X1 U979 ( .A(n937), .B(n921), .Z(n880) );
  XOR2_X1 U980 ( .A(n878), .B(G162), .Z(n879) );
  XNOR2_X1 U981 ( .A(n880), .B(n879), .ZN(n884) );
  XNOR2_X1 U982 ( .A(G160), .B(G164), .ZN(n882) );
  XOR2_X1 U983 ( .A(n882), .B(n881), .Z(n883) );
  XOR2_X1 U984 ( .A(n884), .B(n883), .Z(n889) );
  XOR2_X1 U985 ( .A(KEYINPUT106), .B(KEYINPUT48), .Z(n886) );
  XNOR2_X1 U986 ( .A(KEYINPUT46), .B(KEYINPUT108), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n886), .B(n885), .ZN(n887) );
  XNOR2_X1 U988 ( .A(KEYINPUT107), .B(n887), .ZN(n888) );
  XNOR2_X1 U989 ( .A(n889), .B(n888), .ZN(n899) );
  NAND2_X1 U990 ( .A1(G118), .A2(n786), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G130), .A2(n567), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n897) );
  NAND2_X1 U993 ( .A1(G106), .A2(n892), .ZN(n894) );
  NAND2_X1 U994 ( .A1(G142), .A2(n566), .ZN(n893) );
  NAND2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U996 ( .A(n895), .B(KEYINPUT45), .Z(n896) );
  NOR2_X1 U997 ( .A1(n897), .A2(n896), .ZN(n898) );
  XOR2_X1 U998 ( .A(n899), .B(n898), .Z(n901) );
  XOR2_X1 U999 ( .A(n901), .B(n900), .Z(n902) );
  NOR2_X1 U1000 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U1001 ( .A(n970), .B(KEYINPUT109), .ZN(n904) );
  XNOR2_X1 U1002 ( .A(G171), .B(n976), .ZN(n903) );
  XNOR2_X1 U1003 ( .A(n904), .B(n903), .ZN(n907) );
  XOR2_X1 U1004 ( .A(G286), .B(n905), .Z(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n908), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(KEYINPUT110), .B(n909), .ZN(G397) );
  XNOR2_X1 U1008 ( .A(KEYINPUT111), .B(KEYINPUT49), .ZN(n911) );
  NOR2_X1 U1009 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1010 ( .A(n911), .B(n910), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(G395), .A2(G397), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(n912), .B(KEYINPUT112), .ZN(n913) );
  NAND2_X1 U1013 ( .A1(n914), .A2(n913), .ZN(n915) );
  NOR2_X1 U1014 ( .A1(G401), .A2(n915), .ZN(n916) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n916), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1017 ( .A(G2090), .B(G162), .Z(n917) );
  NOR2_X1 U1018 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1019 ( .A(KEYINPUT51), .B(n919), .Z(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT114), .B(n920), .ZN(n931) );
  NOR2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(n928) );
  XNOR2_X1 U1022 ( .A(G160), .B(G2084), .ZN(n924) );
  NAND2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1025 ( .A1(n928), .A2(n927), .ZN(n929) );
  XNOR2_X1 U1026 ( .A(KEYINPUT113), .B(n929), .ZN(n930) );
  NAND2_X1 U1027 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(n932), .B(KEYINPUT115), .ZN(n934) );
  NAND2_X1 U1029 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1030 ( .A(KEYINPUT116), .B(n935), .ZN(n942) );
  XNOR2_X1 U1031 ( .A(G164), .B(G2078), .ZN(n936) );
  XNOR2_X1 U1032 ( .A(n936), .B(KEYINPUT117), .ZN(n939) );
  XOR2_X1 U1033 ( .A(G2072), .B(n937), .Z(n938) );
  NOR2_X1 U1034 ( .A1(n939), .A2(n938), .ZN(n940) );
  XOR2_X1 U1035 ( .A(KEYINPUT50), .B(n940), .Z(n941) );
  NOR2_X1 U1036 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1037 ( .A(KEYINPUT52), .B(n943), .ZN(n945) );
  INV_X1 U1038 ( .A(KEYINPUT55), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n946), .A2(G29), .ZN(n1027) );
  XOR2_X1 U1041 ( .A(G29), .B(KEYINPUT120), .Z(n968) );
  XNOR2_X1 U1042 ( .A(G2084), .B(G34), .ZN(n947) );
  XNOR2_X1 U1043 ( .A(n947), .B(KEYINPUT54), .ZN(n965) );
  XNOR2_X1 U1044 ( .A(G2090), .B(G35), .ZN(n962) );
  XNOR2_X1 U1045 ( .A(G2067), .B(G26), .ZN(n949) );
  XNOR2_X1 U1046 ( .A(G1991), .B(G25), .ZN(n948) );
  NOR2_X1 U1047 ( .A1(n949), .A2(n948), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(G32), .B(n950), .ZN(n951) );
  NAND2_X1 U1049 ( .A1(n951), .A2(G28), .ZN(n954) );
  XNOR2_X1 U1050 ( .A(KEYINPUT118), .B(G2072), .ZN(n952) );
  XNOR2_X1 U1051 ( .A(G33), .B(n952), .ZN(n953) );
  NOR2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n955) );
  NAND2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n959) );
  XNOR2_X1 U1054 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1056 ( .A(KEYINPUT53), .B(n960), .ZN(n961) );
  NOR2_X1 U1057 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1058 ( .A(n963), .B(KEYINPUT119), .ZN(n964) );
  NOR2_X1 U1059 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1060 ( .A(n966), .B(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(G11), .A2(n969), .ZN(n1025) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n996) );
  XNOR2_X1 U1064 ( .A(n970), .B(G1341), .ZN(n975) );
  XOR2_X1 U1065 ( .A(G1966), .B(G168), .Z(n971) );
  NOR2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1067 ( .A(KEYINPUT57), .B(n973), .ZN(n974) );
  NOR2_X1 U1068 ( .A1(n975), .A2(n974), .ZN(n994) );
  XOR2_X1 U1069 ( .A(G1348), .B(n976), .Z(n977) );
  XNOR2_X1 U1070 ( .A(KEYINPUT121), .B(n977), .ZN(n979) );
  XNOR2_X1 U1071 ( .A(G171), .B(G1961), .ZN(n978) );
  NAND2_X1 U1072 ( .A1(n979), .A2(n978), .ZN(n992) );
  XNOR2_X1 U1073 ( .A(n980), .B(G1956), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n985) );
  XOR2_X1 U1075 ( .A(G1971), .B(G166), .Z(n983) );
  XNOR2_X1 U1076 ( .A(KEYINPUT122), .B(n983), .ZN(n984) );
  NOR2_X1 U1077 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n989) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1080 ( .A(KEYINPUT123), .B(n990), .ZN(n991) );
  NOR2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n1023) );
  INV_X1 U1084 ( .A(G16), .ZN(n1021) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n997) );
  XNOR2_X1 U1086 ( .A(G4), .B(n997), .ZN(n1005) );
  XNOR2_X1 U1087 ( .A(G1341), .B(G19), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G6), .B(G1981), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  XOR2_X1 U1090 ( .A(KEYINPUT124), .B(n1000), .Z(n1002) );
  XNOR2_X1 U1091 ( .A(G1956), .B(G20), .ZN(n1001) );
  NOR2_X1 U1092 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1093 ( .A(n1003), .B(KEYINPUT125), .ZN(n1004) );
  NOR2_X1 U1094 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XNOR2_X1 U1095 ( .A(KEYINPUT60), .B(n1006), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(n1007), .B(KEYINPUT126), .ZN(n1011) );
  XNOR2_X1 U1097 ( .A(G1961), .B(G5), .ZN(n1009) );
  XNOR2_X1 U1098 ( .A(G1966), .B(G21), .ZN(n1008) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1018) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1013) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1012) );
  NOR2_X1 U1103 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1107 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(KEYINPUT61), .B(n1019), .ZN(n1020) );
  NAND2_X1 U1109 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  NAND2_X1 U1110 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NOR2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XNOR2_X1 U1113 ( .A(n1028), .B(KEYINPUT62), .ZN(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT127), .B(n1029), .ZN(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

