

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757;

  XNOR2_X1 U374 ( .A(n429), .B(n505), .ZN(n724) );
  INV_X1 U375 ( .A(G953), .ZN(n748) );
  AND2_X2 U376 ( .A1(n374), .A2(n373), .ZN(n372) );
  NOR2_X2 U377 ( .A1(n676), .A2(n405), .ZN(n605) );
  NOR2_X2 U378 ( .A1(n593), .A2(n592), .ZN(n745) );
  XNOR2_X2 U379 ( .A(n448), .B(KEYINPUT19), .ZN(n597) );
  XNOR2_X2 U380 ( .A(n428), .B(G101), .ZN(n523) );
  NOR2_X1 U381 ( .A1(n663), .A2(n368), .ZN(n456) );
  INV_X1 U382 ( .A(n601), .ZN(n682) );
  XNOR2_X1 U383 ( .A(n381), .B(KEYINPUT45), .ZN(n726) );
  AND2_X1 U384 ( .A1(n468), .A2(n466), .ZN(n580) );
  XNOR2_X1 U385 ( .A(n436), .B(G125), .ZN(n504) );
  NOR2_X1 U386 ( .A1(n628), .A2(n725), .ZN(n629) );
  NOR2_X1 U387 ( .A1(n633), .A2(n725), .ZN(n422) );
  NAND2_X1 U388 ( .A1(n726), .A2(n745), .ZN(n363) );
  NAND2_X1 U389 ( .A1(n618), .A2(n352), .ZN(n381) );
  XNOR2_X1 U390 ( .A(n421), .B(n420), .ZN(n618) );
  XNOR2_X1 U391 ( .A(n452), .B(n451), .ZN(n752) );
  AND2_X1 U392 ( .A1(n617), .A2(n449), .ZN(n643) );
  NOR2_X1 U393 ( .A1(n616), .A2(n615), .ZN(n452) );
  XNOR2_X1 U394 ( .A(n571), .B(n353), .ZN(n405) );
  XNOR2_X1 U395 ( .A(n527), .B(G472), .ZN(n601) );
  XNOR2_X1 U396 ( .A(n719), .B(n718), .ZN(n720) );
  INV_X1 U397 ( .A(n679), .ZN(n440) );
  XOR2_X1 U398 ( .A(n624), .B(KEYINPUT59), .Z(n625) );
  XNOR2_X1 U399 ( .A(n740), .B(n507), .ZN(n429) );
  XNOR2_X1 U400 ( .A(G134), .B(n519), .ZN(n537) );
  XNOR2_X1 U401 ( .A(n524), .B(n488), .ZN(n731) );
  XNOR2_X1 U402 ( .A(n547), .B(n556), .ZN(n740) );
  XNOR2_X1 U403 ( .A(n504), .B(n503), .ZN(n547) );
  NAND2_X1 U404 ( .A1(n475), .A2(n432), .ZN(n519) );
  XNOR2_X1 U405 ( .A(n472), .B(n471), .ZN(n620) );
  INV_X1 U406 ( .A(n425), .ZN(n486) );
  INV_X1 U407 ( .A(G146), .ZN(n436) );
  XNOR2_X1 U408 ( .A(G119), .B(KEYINPUT3), .ZN(n485) );
  XNOR2_X1 U409 ( .A(KEYINPUT87), .B(G902), .ZN(n472) );
  XNOR2_X1 U410 ( .A(G113), .B(G116), .ZN(n425) );
  INV_X1 U411 ( .A(KEYINPUT68), .ZN(n428) );
  XOR2_X1 U412 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n502) );
  XNOR2_X2 U413 ( .A(n497), .B(n496), .ZN(n448) );
  XNOR2_X1 U414 ( .A(n489), .B(G107), .ZN(n732) );
  XNOR2_X1 U415 ( .A(n741), .B(G146), .ZN(n558) );
  XNOR2_X1 U416 ( .A(n500), .B(n499), .ZN(n679) );
  XNOR2_X1 U417 ( .A(n537), .B(n520), .ZN(n741) );
  XNOR2_X1 U418 ( .A(KEYINPUT4), .B(G131), .ZN(n520) );
  XNOR2_X1 U419 ( .A(n490), .B(n732), .ZN(n407) );
  XNOR2_X1 U420 ( .A(n523), .B(KEYINPUT71), .ZN(n490) );
  NAND2_X1 U421 ( .A1(n444), .A2(n443), .ZN(n442) );
  NOR2_X1 U422 ( .A1(n447), .A2(G902), .ZN(n444) );
  NOR2_X1 U423 ( .A1(G902), .A2(n712), .ZN(n559) );
  AND2_X1 U424 ( .A1(n621), .A2(KEYINPUT2), .ZN(n453) );
  XNOR2_X1 U425 ( .A(n470), .B(n498), .ZN(n510) );
  XOR2_X1 U426 ( .A(KEYINPUT20), .B(KEYINPUT91), .Z(n498) );
  NAND2_X1 U427 ( .A1(n620), .A2(G234), .ZN(n470) );
  XOR2_X1 U428 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n509) );
  NAND2_X1 U429 ( .A1(n412), .A2(n416), .ZN(n411) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n495) );
  XNOR2_X1 U431 ( .A(n521), .B(KEYINPUT73), .ZN(n388) );
  XOR2_X1 U432 ( .A(G137), .B(KEYINPUT5), .Z(n522) );
  NOR2_X1 U433 ( .A1(n577), .A2(n464), .ZN(n463) );
  INV_X1 U434 ( .A(n756), .ZN(n464) );
  NAND2_X1 U435 ( .A1(n394), .A2(n393), .ZN(n392) );
  NOR2_X1 U436 ( .A1(n384), .A2(n643), .ZN(n394) );
  NAND2_X1 U437 ( .A1(n396), .A2(n395), .ZN(n384) );
  AND2_X1 U438 ( .A1(n399), .A2(n398), .ZN(n397) );
  NAND2_X1 U439 ( .A1(n371), .A2(n370), .ZN(n369) );
  NAND2_X1 U440 ( .A1(n380), .A2(n377), .ZN(n370) );
  AND2_X1 U441 ( .A1(n376), .A2(KEYINPUT65), .ZN(n371) );
  NAND2_X1 U442 ( .A1(n605), .A2(n682), .ZN(n685) );
  INV_X1 U443 ( .A(KEYINPUT105), .ZN(n469) );
  AND2_X1 U444 ( .A1(n438), .A2(n442), .ZN(n427) );
  NOR2_X1 U445 ( .A1(G953), .A2(G237), .ZN(n548) );
  XNOR2_X1 U446 ( .A(KEYINPUT10), .B(KEYINPUT70), .ZN(n503) );
  XNOR2_X1 U447 ( .A(n544), .B(n433), .ZN(n546) );
  XNOR2_X1 U448 ( .A(n545), .B(n434), .ZN(n433) );
  INV_X1 U449 ( .A(KEYINPUT96), .ZN(n434) );
  XNOR2_X1 U450 ( .A(G113), .B(G140), .ZN(n540) );
  XOR2_X1 U451 ( .A(G122), .B(G104), .Z(n541) );
  XNOR2_X1 U452 ( .A(n558), .B(n457), .ZN(n712) );
  XNOR2_X1 U453 ( .A(n557), .B(n459), .ZN(n458) );
  XNOR2_X1 U454 ( .A(n569), .B(KEYINPUT41), .ZN(n688) );
  XNOR2_X1 U455 ( .A(n575), .B(KEYINPUT39), .ZN(n591) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n616) );
  INV_X1 U457 ( .A(KEYINPUT22), .ZN(n400) );
  NAND2_X1 U458 ( .A1(n667), .A2(n440), .ZN(n402) );
  NOR2_X1 U459 ( .A1(n571), .A2(n564), .ZN(n570) );
  AND2_X1 U460 ( .A1(n682), .A2(n562), .ZN(n563) );
  NAND2_X1 U461 ( .A1(n445), .A2(n442), .ZN(n461) );
  NOR2_X1 U462 ( .A1(n441), .A2(n389), .ZN(n445) );
  AND2_X1 U463 ( .A1(n526), .A2(n630), .ZN(n527) );
  NOR2_X1 U464 ( .A1(n616), .A2(n610), .ZN(n617) );
  XNOR2_X1 U465 ( .A(KEYINPUT86), .B(n627), .ZN(n725) );
  INV_X1 U466 ( .A(KEYINPUT15), .ZN(n471) );
  NAND2_X1 U467 ( .A1(n363), .A2(n358), .ZN(n376) );
  NAND2_X1 U468 ( .A1(n379), .A2(n378), .ZN(n377) );
  NAND2_X1 U469 ( .A1(n622), .A2(n360), .ZN(n378) );
  NAND2_X1 U470 ( .A1(n453), .A2(n619), .ZN(n379) );
  XNOR2_X1 U471 ( .A(n477), .B(n476), .ZN(n478) );
  INV_X1 U472 ( .A(KEYINPUT18), .ZN(n476) );
  XNOR2_X1 U473 ( .A(n406), .B(n511), .ZN(n447) );
  NAND2_X1 U474 ( .A1(n510), .A2(G217), .ZN(n406) );
  XNOR2_X1 U475 ( .A(KEYINPUT76), .B(KEYINPUT92), .ZN(n508) );
  INV_X1 U476 ( .A(KEYINPUT84), .ZN(n420) );
  XNOR2_X1 U477 ( .A(KEYINPUT98), .B(KEYINPUT12), .ZN(n542) );
  XNOR2_X1 U478 ( .A(G143), .B(G131), .ZN(n545) );
  XOR2_X1 U479 ( .A(G137), .B(G140), .Z(n556) );
  XNOR2_X1 U480 ( .A(n555), .B(n460), .ZN(n459) );
  INV_X1 U481 ( .A(KEYINPUT77), .ZN(n460) );
  XNOR2_X1 U482 ( .A(n366), .B(n365), .ZN(n665) );
  INV_X1 U483 ( .A(KEYINPUT108), .ZN(n365) );
  NAND2_X1 U484 ( .A1(n669), .A2(n668), .ZN(n366) );
  XNOR2_X1 U485 ( .A(n568), .B(n367), .ZN(n669) );
  INV_X1 U486 ( .A(KEYINPUT38), .ZN(n367) );
  NAND2_X1 U487 ( .A1(n605), .A2(n612), .ZN(n607) );
  NOR2_X1 U488 ( .A1(n579), .A2(n578), .ZN(n667) );
  NOR2_X1 U489 ( .A1(n679), .A2(n518), .ZN(n562) );
  NAND2_X1 U490 ( .A1(n447), .A2(G902), .ZN(n446) );
  AND2_X1 U491 ( .A1(n724), .A2(n447), .ZN(n441) );
  INV_X1 U492 ( .A(G902), .ZN(n526) );
  XNOR2_X1 U493 ( .A(n558), .B(n386), .ZN(n630) );
  XNOR2_X1 U494 ( .A(n525), .B(n387), .ZN(n386) );
  XNOR2_X1 U495 ( .A(n388), .B(n522), .ZN(n387) );
  XNOR2_X1 U496 ( .A(G104), .B(G110), .ZN(n489) );
  XNOR2_X1 U497 ( .A(n487), .B(KEYINPUT16), .ZN(n488) );
  INV_X1 U498 ( .A(G122), .ZN(n487) );
  XOR2_X1 U499 ( .A(G128), .B(G119), .Z(n506) );
  XNOR2_X1 U500 ( .A(G122), .B(KEYINPUT99), .ZN(n530) );
  XOR2_X1 U501 ( .A(KEYINPUT100), .B(KEYINPUT9), .Z(n531) );
  XNOR2_X1 U502 ( .A(G116), .B(G107), .ZN(n529) );
  XNOR2_X1 U503 ( .A(n431), .B(n430), .ZN(n534) );
  INV_X1 U504 ( .A(KEYINPUT8), .ZN(n430) );
  NAND2_X1 U505 ( .A1(n748), .A2(G234), .ZN(n431) );
  INV_X1 U506 ( .A(KEYINPUT85), .ZN(n496) );
  XNOR2_X1 U507 ( .A(n599), .B(KEYINPUT31), .ZN(n600) );
  INV_X1 U508 ( .A(KEYINPUT94), .ZN(n599) );
  INV_X1 U509 ( .A(n572), .ZN(n467) );
  INV_X1 U510 ( .A(n568), .ZN(n590) );
  XOR2_X1 U511 ( .A(n630), .B(KEYINPUT62), .Z(n631) );
  XNOR2_X1 U512 ( .A(n549), .B(n435), .ZN(n624) );
  XNOR2_X1 U513 ( .A(n550), .B(n354), .ZN(n435) );
  XNOR2_X1 U514 ( .A(n710), .B(n357), .ZN(n424) );
  NAND2_X1 U515 ( .A1(n362), .A2(G210), .ZN(n710) );
  INV_X1 U516 ( .A(n725), .ZN(n423) );
  INV_X2 U517 ( .A(n363), .ZN(n380) );
  XNOR2_X1 U518 ( .A(n391), .B(KEYINPUT42), .ZN(n753) );
  XNOR2_X1 U519 ( .A(n390), .B(n355), .ZN(n754) );
  INV_X1 U520 ( .A(KEYINPUT35), .ZN(n385) );
  INV_X1 U521 ( .A(n608), .ZN(n454) );
  XNOR2_X1 U522 ( .A(KEYINPUT66), .B(KEYINPUT32), .ZN(n451) );
  NOR2_X1 U523 ( .A1(n682), .A2(n450), .ZN(n449) );
  INV_X1 U524 ( .A(n461), .ZN(n450) );
  NOR2_X1 U525 ( .A1(n578), .A2(n561), .ZN(n651) );
  XNOR2_X1 U526 ( .A(n723), .B(n724), .ZN(n417) );
  XNOR2_X1 U527 ( .A(n716), .B(n717), .ZN(n364) );
  INV_X1 U528 ( .A(n405), .ZN(n610) );
  AND2_X1 U529 ( .A1(n392), .A2(n397), .ZN(n352) );
  XOR2_X1 U530 ( .A(KEYINPUT1), .B(KEYINPUT67), .Z(n353) );
  NOR2_X1 U531 ( .A1(n651), .A2(n653), .ZN(n664) );
  INV_X1 U532 ( .A(n664), .ZN(n416) );
  AND2_X1 U533 ( .A1(G214), .A2(n548), .ZN(n354) );
  AND2_X1 U534 ( .A1(n617), .A2(n418), .ZN(n635) );
  XOR2_X1 U535 ( .A(KEYINPUT107), .B(KEYINPUT40), .Z(n355) );
  XOR2_X1 U536 ( .A(KEYINPUT46), .B(KEYINPUT64), .Z(n356) );
  XOR2_X1 U537 ( .A(n709), .B(n708), .Z(n357) );
  AND2_X1 U538 ( .A1(n453), .A2(KEYINPUT74), .ZN(n358) );
  AND2_X1 U539 ( .A1(n377), .A2(n623), .ZN(n359) );
  INV_X1 U540 ( .A(KEYINPUT44), .ZN(n395) );
  XOR2_X1 U541 ( .A(KEYINPUT74), .B(KEYINPUT2), .Z(n360) );
  XOR2_X1 U542 ( .A(n711), .B(KEYINPUT56), .Z(n361) );
  INV_X1 U543 ( .A(KEYINPUT65), .ZN(n623) );
  NAND2_X1 U544 ( .A1(n372), .A2(n369), .ZN(n362) );
  NAND2_X1 U545 ( .A1(n372), .A2(n369), .ZN(n715) );
  AND2_X1 U546 ( .A1(n380), .A2(n360), .ZN(n703) );
  XNOR2_X1 U547 ( .A(n380), .B(n619), .ZN(n408) );
  NAND2_X1 U548 ( .A1(n380), .A2(n359), .ZN(n373) );
  NOR2_X1 U549 ( .A1(n364), .A2(n725), .ZN(G54) );
  NAND2_X1 U550 ( .A1(n424), .A2(n423), .ZN(n419) );
  NOR2_X2 U551 ( .A1(n368), .A2(n685), .ZN(n437) );
  NOR2_X1 U552 ( .A1(n368), .A2(n402), .ZN(n401) );
  NOR2_X1 U553 ( .A1(n368), .A2(n603), .ZN(n638) );
  XNOR2_X2 U554 ( .A(n598), .B(KEYINPUT0), .ZN(n368) );
  NAND2_X1 U555 ( .A1(n375), .A2(n623), .ZN(n374) );
  INV_X1 U556 ( .A(n376), .ZN(n375) );
  BUF_X1 U557 ( .A(n654), .Z(n382) );
  NAND2_X1 U558 ( .A1(n383), .A2(n609), .ZN(n421) );
  NOR2_X1 U559 ( .A1(n403), .A2(n635), .ZN(n383) );
  NOR2_X1 U560 ( .A1(n396), .A2(n395), .ZN(n403) );
  XNOR2_X2 U561 ( .A(n404), .B(n385), .ZN(n396) );
  XNOR2_X1 U562 ( .A(n396), .B(G122), .ZN(G24) );
  INV_X1 U563 ( .A(n446), .ZN(n389) );
  NAND2_X1 U564 ( .A1(n753), .A2(n754), .ZN(n576) );
  NAND2_X1 U565 ( .A1(n591), .A2(n651), .ZN(n390) );
  NAND2_X1 U566 ( .A1(n688), .A2(n570), .ZN(n391) );
  INV_X1 U567 ( .A(n752), .ZN(n393) );
  NAND2_X1 U568 ( .A1(n643), .A2(KEYINPUT44), .ZN(n398) );
  NAND2_X1 U569 ( .A1(n752), .A2(KEYINPUT44), .ZN(n399) );
  NAND2_X1 U570 ( .A1(n455), .A2(n454), .ZN(n404) );
  XNOR2_X2 U571 ( .A(n559), .B(G469), .ZN(n571) );
  XNOR2_X2 U572 ( .A(n427), .B(KEYINPUT69), .ZN(n676) );
  XNOR2_X1 U573 ( .A(n407), .B(n731), .ZN(n491) );
  XNOR2_X1 U574 ( .A(n407), .B(n458), .ZN(n457) );
  AND2_X1 U575 ( .A1(n408), .A2(KEYINPUT2), .ZN(n697) );
  NAND2_X1 U576 ( .A1(n410), .A2(n409), .ZN(n415) );
  NOR2_X1 U577 ( .A1(n638), .A2(KEYINPUT95), .ZN(n409) );
  INV_X1 U578 ( .A(n654), .ZN(n410) );
  XNOR2_X2 U579 ( .A(n437), .B(n600), .ZN(n654) );
  NOR2_X2 U580 ( .A1(n413), .A2(n411), .ZN(n604) );
  NAND2_X1 U581 ( .A1(n638), .A2(KEYINPUT95), .ZN(n412) );
  NAND2_X1 U582 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U583 ( .A1(n654), .A2(KEYINPUT95), .ZN(n414) );
  XNOR2_X1 U584 ( .A(n576), .B(n356), .ZN(n465) );
  XNOR2_X1 U585 ( .A(n602), .B(n469), .ZN(n468) );
  NOR2_X1 U586 ( .A1(n417), .A2(n725), .ZN(G66) );
  NOR2_X1 U587 ( .A1(n678), .A2(n612), .ZN(n418) );
  XNOR2_X1 U588 ( .A(n419), .B(n361), .ZN(G51) );
  XNOR2_X1 U589 ( .A(n422), .B(n634), .ZN(G57) );
  XNOR2_X1 U590 ( .A(n426), .B(n504), .ZN(n479) );
  INV_X1 U591 ( .A(n519), .ZN(n426) );
  NAND2_X1 U592 ( .A1(n465), .A2(n463), .ZN(n462) );
  XNOR2_X1 U593 ( .A(n462), .B(n583), .ZN(n593) );
  NAND2_X1 U594 ( .A1(n473), .A2(G143), .ZN(n432) );
  NOR2_X1 U595 ( .A1(n441), .A2(n439), .ZN(n438) );
  NAND2_X1 U596 ( .A1(n446), .A2(n440), .ZN(n439) );
  INV_X1 U597 ( .A(n724), .ZN(n443) );
  NOR2_X1 U598 ( .A1(n584), .A2(n448), .ZN(n554) );
  XNOR2_X1 U599 ( .A(n456), .B(KEYINPUT34), .ZN(n455) );
  NAND2_X1 U600 ( .A1(n461), .A2(n572), .ZN(n518) );
  XNOR2_X1 U601 ( .A(n461), .B(KEYINPUT102), .ZN(n678) );
  NOR2_X1 U602 ( .A1(n574), .A2(n467), .ZN(n466) );
  NOR2_X2 U603 ( .A1(n676), .A2(n571), .ZN(n602) );
  XNOR2_X2 U604 ( .A(n486), .B(n485), .ZN(n524) );
  INV_X1 U605 ( .A(n556), .ZN(n557) );
  INV_X1 U606 ( .A(KEYINPUT74), .ZN(n619) );
  XNOR2_X1 U607 ( .A(n607), .B(n606), .ZN(n663) );
  BUF_X1 U608 ( .A(n567), .Z(n568) );
  XNOR2_X1 U609 ( .A(n721), .B(n720), .ZN(n722) );
  XOR2_X1 U610 ( .A(KEYINPUT48), .B(KEYINPUT83), .Z(n583) );
  INV_X1 U611 ( .A(G128), .ZN(n473) );
  INV_X1 U612 ( .A(G143), .ZN(n474) );
  NAND2_X1 U613 ( .A1(n474), .A2(G128), .ZN(n475) );
  NAND2_X1 U614 ( .A1(G224), .A2(n748), .ZN(n477) );
  XNOR2_X1 U615 ( .A(n479), .B(n478), .ZN(n484) );
  XOR2_X1 U616 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n481) );
  XNOR2_X1 U617 ( .A(KEYINPUT78), .B(KEYINPUT17), .ZN(n480) );
  XNOR2_X1 U618 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U619 ( .A(KEYINPUT4), .B(n482), .ZN(n483) );
  XNOR2_X1 U620 ( .A(n484), .B(n483), .ZN(n492) );
  XNOR2_X1 U621 ( .A(n491), .B(n492), .ZN(n706) );
  INV_X1 U622 ( .A(n620), .ZN(n622) );
  NOR2_X1 U623 ( .A1(n706), .A2(n622), .ZN(n494) );
  NAND2_X1 U624 ( .A1(G210), .A2(n495), .ZN(n493) );
  XNOR2_X1 U625 ( .A(n494), .B(n493), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G214), .A2(n495), .ZN(n668) );
  NAND2_X1 U627 ( .A1(n567), .A2(n668), .ZN(n497) );
  XOR2_X1 U628 ( .A(KEYINPUT21), .B(KEYINPUT93), .Z(n500) );
  NAND2_X1 U629 ( .A1(G221), .A2(n510), .ZN(n499) );
  NAND2_X1 U630 ( .A1(G221), .A2(n534), .ZN(n501) );
  XNOR2_X1 U631 ( .A(n502), .B(n501), .ZN(n505) );
  XNOR2_X1 U632 ( .A(G110), .B(n506), .ZN(n507) );
  XNOR2_X1 U633 ( .A(n509), .B(n508), .ZN(n511) );
  NAND2_X1 U634 ( .A1(G234), .A2(G237), .ZN(n512) );
  XNOR2_X1 U635 ( .A(n512), .B(KEYINPUT14), .ZN(n662) );
  NAND2_X1 U636 ( .A1(G953), .A2(n526), .ZN(n513) );
  NAND2_X1 U637 ( .A1(n662), .A2(n513), .ZN(n515) );
  NOR2_X1 U638 ( .A1(G953), .A2(G952), .ZN(n514) );
  NOR2_X1 U639 ( .A1(n515), .A2(n514), .ZN(n595) );
  NAND2_X1 U640 ( .A1(G953), .A2(G900), .ZN(n516) );
  NAND2_X1 U641 ( .A1(n595), .A2(n516), .ZN(n517) );
  XOR2_X1 U642 ( .A(KEYINPUT80), .B(n517), .Z(n572) );
  NAND2_X1 U643 ( .A1(n548), .A2(G210), .ZN(n521) );
  XNOR2_X1 U644 ( .A(n523), .B(n524), .ZN(n525) );
  XNOR2_X1 U645 ( .A(KEYINPUT6), .B(n601), .ZN(n612) );
  NAND2_X1 U646 ( .A1(n562), .A2(n612), .ZN(n528) );
  XNOR2_X1 U647 ( .A(KEYINPUT103), .B(n528), .ZN(n553) );
  XNOR2_X1 U648 ( .A(n529), .B(KEYINPUT7), .ZN(n533) );
  XNOR2_X1 U649 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U650 ( .A(n533), .B(n532), .Z(n536) );
  NAND2_X1 U651 ( .A1(G217), .A2(n534), .ZN(n535) );
  XNOR2_X1 U652 ( .A(n536), .B(n535), .ZN(n538) );
  XNOR2_X1 U653 ( .A(n538), .B(n537), .ZN(n719) );
  NOR2_X1 U654 ( .A1(G902), .A2(n719), .ZN(n539) );
  XOR2_X1 U655 ( .A(G478), .B(n539), .Z(n578) );
  XNOR2_X1 U656 ( .A(KEYINPUT13), .B(G475), .ZN(n552) );
  XNOR2_X1 U657 ( .A(n541), .B(n540), .ZN(n550) );
  XOR2_X1 U658 ( .A(KEYINPUT97), .B(KEYINPUT11), .Z(n543) );
  XNOR2_X1 U659 ( .A(n543), .B(n542), .ZN(n544) );
  XOR2_X1 U660 ( .A(n547), .B(n546), .Z(n549) );
  NOR2_X1 U661 ( .A1(G902), .A2(n624), .ZN(n551) );
  XNOR2_X1 U662 ( .A(n552), .B(n551), .ZN(n579) );
  INV_X1 U663 ( .A(n579), .ZN(n561) );
  NAND2_X1 U664 ( .A1(n553), .A2(n651), .ZN(n584) );
  XNOR2_X1 U665 ( .A(n554), .B(KEYINPUT36), .ZN(n560) );
  NAND2_X1 U666 ( .A1(G227), .A2(n748), .ZN(n555) );
  NAND2_X1 U667 ( .A1(n560), .A2(n610), .ZN(n656) );
  NAND2_X1 U668 ( .A1(n561), .A2(n578), .ZN(n644) );
  INV_X1 U669 ( .A(n644), .ZN(n653) );
  XOR2_X1 U670 ( .A(KEYINPUT28), .B(n563), .Z(n564) );
  NAND2_X1 U671 ( .A1(n570), .A2(n597), .ZN(n647) );
  NOR2_X1 U672 ( .A1(n664), .A2(n647), .ZN(n565) );
  XNOR2_X1 U673 ( .A(n565), .B(KEYINPUT47), .ZN(n566) );
  NAND2_X1 U674 ( .A1(n656), .A2(n566), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n665), .A2(n667), .ZN(n569) );
  NAND2_X1 U676 ( .A1(n682), .A2(n668), .ZN(n573) );
  XNOR2_X1 U677 ( .A(KEYINPUT30), .B(n573), .ZN(n574) );
  NAND2_X1 U678 ( .A1(n580), .A2(n669), .ZN(n575) );
  NAND2_X1 U679 ( .A1(n579), .A2(n578), .ZN(n608) );
  NOR2_X1 U680 ( .A1(n590), .A2(n608), .ZN(n581) );
  NAND2_X1 U681 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U682 ( .A(n582), .B(KEYINPUT106), .ZN(n756) );
  INV_X1 U683 ( .A(n584), .ZN(n585) );
  NAND2_X1 U684 ( .A1(n585), .A2(n668), .ZN(n586) );
  NOR2_X1 U685 ( .A1(n610), .A2(n586), .ZN(n588) );
  XOR2_X1 U686 ( .A(KEYINPUT43), .B(KEYINPUT104), .Z(n587) );
  XNOR2_X1 U687 ( .A(n588), .B(n587), .ZN(n589) );
  NAND2_X1 U688 ( .A1(n590), .A2(n589), .ZN(n660) );
  NAND2_X1 U689 ( .A1(n591), .A2(n653), .ZN(n659) );
  NAND2_X1 U690 ( .A1(n660), .A2(n659), .ZN(n592) );
  XNOR2_X1 U691 ( .A(G898), .B(KEYINPUT90), .ZN(n735) );
  NAND2_X1 U692 ( .A1(n735), .A2(G953), .ZN(n594) );
  AND2_X1 U693 ( .A1(n595), .A2(n594), .ZN(n596) );
  NAND2_X1 U694 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n602), .A2(n601), .ZN(n603) );
  XNOR2_X1 U696 ( .A(n604), .B(KEYINPUT101), .ZN(n609) );
  INV_X1 U697 ( .A(n678), .ZN(n611) );
  XOR2_X1 U698 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n606) );
  OR2_X1 U699 ( .A1(n612), .A2(n611), .ZN(n613) );
  NOR2_X1 U700 ( .A1(n405), .A2(n613), .ZN(n614) );
  XNOR2_X1 U701 ( .A(n614), .B(KEYINPUT79), .ZN(n615) );
  XNOR2_X1 U702 ( .A(n620), .B(KEYINPUT81), .ZN(n621) );
  NAND2_X1 U703 ( .A1(n715), .A2(G475), .ZN(n626) );
  XNOR2_X1 U704 ( .A(n626), .B(n625), .ZN(n628) );
  NOR2_X1 U705 ( .A1(G952), .A2(n748), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U707 ( .A(KEYINPUT63), .ZN(n634) );
  NAND2_X1 U708 ( .A1(n715), .A2(G472), .ZN(n632) );
  XNOR2_X1 U709 ( .A(n632), .B(n631), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n635), .B(G101), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT109), .ZN(G3) );
  NAND2_X1 U712 ( .A1(n638), .A2(n651), .ZN(n637) );
  XNOR2_X1 U713 ( .A(n637), .B(G104), .ZN(G6) );
  XNOR2_X1 U714 ( .A(G107), .B(KEYINPUT27), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT110), .B(KEYINPUT26), .Z(n640) );
  NAND2_X1 U716 ( .A1(n638), .A2(n653), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n640), .B(n639), .ZN(n641) );
  XNOR2_X1 U718 ( .A(n642), .B(n641), .ZN(G9) );
  XOR2_X1 U719 ( .A(G110), .B(n643), .Z(G12) );
  NOR2_X1 U720 ( .A1(n644), .A2(n647), .ZN(n646) );
  XNOR2_X1 U721 ( .A(G128), .B(KEYINPUT29), .ZN(n645) );
  XNOR2_X1 U722 ( .A(n646), .B(n645), .ZN(G30) );
  INV_X1 U723 ( .A(n651), .ZN(n648) );
  NOR2_X1 U724 ( .A1(n648), .A2(n647), .ZN(n649) );
  XOR2_X1 U725 ( .A(KEYINPUT112), .B(n649), .Z(n650) );
  XNOR2_X1 U726 ( .A(G146), .B(n650), .ZN(G48) );
  NAND2_X1 U727 ( .A1(n382), .A2(n651), .ZN(n652) );
  XNOR2_X1 U728 ( .A(n652), .B(G113), .ZN(G15) );
  NAND2_X1 U729 ( .A1(n382), .A2(n653), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n655), .B(G116), .ZN(G18) );
  XNOR2_X1 U731 ( .A(KEYINPUT37), .B(KEYINPUT113), .ZN(n657) );
  XNOR2_X1 U732 ( .A(n657), .B(n656), .ZN(n658) );
  XNOR2_X1 U733 ( .A(G125), .B(n658), .ZN(G27) );
  XNOR2_X1 U734 ( .A(G134), .B(n659), .ZN(G36) );
  XNOR2_X1 U735 ( .A(G140), .B(KEYINPUT114), .ZN(n661) );
  XNOR2_X1 U736 ( .A(n661), .B(n660), .ZN(G42) );
  XNOR2_X1 U737 ( .A(KEYINPUT118), .B(KEYINPUT53), .ZN(n705) );
  NAND2_X1 U738 ( .A1(G952), .A2(n662), .ZN(n694) );
  NAND2_X1 U739 ( .A1(n665), .A2(n416), .ZN(n666) );
  XOR2_X1 U740 ( .A(KEYINPUT116), .B(n666), .Z(n674) );
  INV_X1 U741 ( .A(n667), .ZN(n671) );
  NOR2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U744 ( .A(KEYINPUT115), .B(n672), .Z(n673) );
  NOR2_X1 U745 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U746 ( .A1(n663), .A2(n675), .ZN(n691) );
  NAND2_X1 U747 ( .A1(n405), .A2(n676), .ZN(n677) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT50), .ZN(n684) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  XNOR2_X1 U750 ( .A(KEYINPUT49), .B(n680), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n686) );
  NAND2_X1 U753 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U754 ( .A(KEYINPUT51), .B(n687), .ZN(n689) );
  INV_X1 U755 ( .A(n688), .ZN(n698) );
  NOR2_X1 U756 ( .A1(n689), .A2(n698), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n692) );
  XNOR2_X1 U758 ( .A(n692), .B(KEYINPUT52), .ZN(n693) );
  NOR2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U760 ( .A(KEYINPUT117), .B(n695), .Z(n696) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n701) );
  NOR2_X1 U762 ( .A1(n663), .A2(n698), .ZN(n699) );
  NOR2_X1 U763 ( .A1(G953), .A2(n699), .ZN(n700) );
  NAND2_X1 U764 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n705), .B(n704), .ZN(G75) );
  XNOR2_X1 U767 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n709) );
  BUF_X1 U768 ( .A(n706), .Z(n707) );
  XNOR2_X1 U769 ( .A(n707), .B(KEYINPUT55), .ZN(n708) );
  XNOR2_X1 U770 ( .A(KEYINPUT82), .B(KEYINPUT120), .ZN(n711) );
  XNOR2_X1 U771 ( .A(KEYINPUT58), .B(KEYINPUT121), .ZN(n714) );
  XNOR2_X1 U772 ( .A(n712), .B(KEYINPUT57), .ZN(n713) );
  XNOR2_X1 U773 ( .A(n714), .B(n713), .ZN(n717) );
  NAND2_X1 U774 ( .A1(n362), .A2(G469), .ZN(n716) );
  NAND2_X1 U775 ( .A1(n362), .A2(G478), .ZN(n721) );
  XOR2_X1 U776 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n718) );
  NOR2_X1 U777 ( .A1(n725), .A2(n722), .ZN(G63) );
  NAND2_X1 U778 ( .A1(G217), .A2(n362), .ZN(n723) );
  NAND2_X1 U779 ( .A1(n748), .A2(n726), .ZN(n730) );
  NAND2_X1 U780 ( .A1(G953), .A2(G224), .ZN(n727) );
  XNOR2_X1 U781 ( .A(n727), .B(KEYINPUT61), .ZN(n728) );
  NAND2_X1 U782 ( .A1(n728), .A2(n735), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n730), .A2(n729), .ZN(n739) );
  XNOR2_X1 U784 ( .A(n731), .B(KEYINPUT124), .ZN(n734) );
  XNOR2_X1 U785 ( .A(G101), .B(n732), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n734), .B(n733), .ZN(n737) );
  NOR2_X1 U787 ( .A1(n735), .A2(n748), .ZN(n736) );
  NOR2_X1 U788 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U789 ( .A(n739), .B(n738), .ZN(G69) );
  XNOR2_X1 U790 ( .A(n741), .B(n740), .ZN(n746) );
  XNOR2_X1 U791 ( .A(G227), .B(n746), .ZN(n742) );
  NAND2_X1 U792 ( .A1(n742), .A2(G900), .ZN(n743) );
  NAND2_X1 U793 ( .A1(G953), .A2(n743), .ZN(n744) );
  XNOR2_X1 U794 ( .A(n744), .B(KEYINPUT126), .ZN(n751) );
  XNOR2_X1 U795 ( .A(KEYINPUT125), .B(n745), .ZN(n747) );
  XNOR2_X1 U796 ( .A(n747), .B(n746), .ZN(n749) );
  NAND2_X1 U797 ( .A1(n749), .A2(n748), .ZN(n750) );
  NAND2_X1 U798 ( .A1(n751), .A2(n750), .ZN(G72) );
  XOR2_X1 U799 ( .A(n752), .B(G119), .Z(G21) );
  XNOR2_X1 U800 ( .A(G137), .B(n753), .ZN(G39) );
  XOR2_X1 U801 ( .A(G131), .B(n754), .Z(n755) );
  XNOR2_X1 U802 ( .A(KEYINPUT127), .B(n755), .ZN(G33) );
  XOR2_X1 U803 ( .A(G143), .B(n756), .Z(n757) );
  XNOR2_X1 U804 ( .A(KEYINPUT111), .B(n757), .ZN(G45) );
endmodule

