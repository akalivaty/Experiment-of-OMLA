//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 1 0 0 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n681, new_n682, new_n683, new_n684, new_n685, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n792, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n876,
    new_n877, new_n879, new_n880, new_n881, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n997, new_n998, new_n999, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1006, new_n1007;
  NAND2_X1  g000(.A1(G228gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(new_n202), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT77), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G155gat), .B2(G162gat), .ZN(new_n205));
  OR2_X1    g004(.A1(G141gat), .A2(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(G141gat), .A2(G148gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT2), .ZN(new_n209));
  AOI21_X1  g008(.A(new_n209), .B1(G155gat), .B2(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n205), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  AND2_X1   g010(.A1(G155gat), .A2(G162gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(G155gat), .A2(G162gat), .ZN(new_n213));
  NOR2_X1   g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(new_n214), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n206), .B(new_n207), .C1(new_n212), .C2(new_n209), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(new_n217), .A3(new_n205), .ZN(new_n218));
  AND2_X1   g017(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT75), .ZN(new_n221));
  AND2_X1   g020(.A1(G211gat), .A2(G218gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G211gat), .A2(G218gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G211gat), .ZN(new_n225));
  INV_X1    g024(.A(G218gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G211gat), .A2(G218gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT75), .A3(new_n228), .ZN(new_n229));
  AND2_X1   g028(.A1(new_n224), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT74), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n231), .B1(new_n222), .B2(KEYINPUT22), .ZN(new_n232));
  XNOR2_X1  g031(.A(G197gat), .B(G204gat), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT22), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n228), .A2(KEYINPUT74), .A3(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT76), .ZN(new_n237));
  NOR3_X1   g036(.A1(new_n230), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n235), .ZN(new_n239));
  AND2_X1   g038(.A1(G197gat), .A2(G204gat), .ZN(new_n240));
  NOR2_X1   g039(.A1(G197gat), .A2(G204gat), .ZN(new_n241));
  NOR2_X1   g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT74), .B1(new_n228), .B2(new_n234), .ZN(new_n243));
  NOR3_X1   g042(.A1(new_n239), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n224), .A2(new_n229), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT76), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n238), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT79), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n248), .B1(new_n244), .B2(new_n245), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n230), .A2(KEYINPUT79), .A3(new_n236), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(KEYINPUT80), .B(new_n220), .C1(new_n247), .C2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  OAI211_X1 g053(.A(new_n249), .B(new_n250), .C1(new_n238), .C2(new_n246), .ZN(new_n255));
  AOI21_X1  g054(.A(KEYINPUT80), .B1(new_n255), .B2(new_n220), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n219), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  OAI22_X1  g056(.A1(new_n238), .A2(new_n246), .B1(new_n245), .B2(new_n244), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n215), .A2(new_n218), .ZN(new_n259));
  AOI21_X1  g058(.A(KEYINPUT29), .B1(new_n259), .B2(new_n253), .ZN(new_n260));
  NOR2_X1   g059(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n203), .B1(new_n257), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT81), .B1(new_n258), .B2(new_n260), .ZN(new_n264));
  AND2_X1   g063(.A1(new_n264), .A2(new_n203), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n258), .A2(new_n220), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(new_n253), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n267), .A2(new_n219), .ZN(new_n268));
  OR3_X1    g067(.A1(new_n258), .A2(new_n260), .A3(KEYINPUT81), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  OAI21_X1  g069(.A(G22gat), .B1(new_n263), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n265), .A2(new_n268), .A3(new_n269), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n220), .B1(new_n247), .B2(new_n251), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT80), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n276), .A2(new_n253), .A3(new_n252), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n261), .B1(new_n277), .B2(new_n219), .ZN(new_n278));
  OAI211_X1 g077(.A(new_n272), .B(new_n273), .C1(new_n278), .C2(new_n203), .ZN(new_n279));
  XNOR2_X1  g078(.A(G78gat), .B(G106gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT31), .B(G50gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n280), .B(new_n281), .Z(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n271), .A2(new_n279), .A3(new_n283), .ZN(new_n284));
  AND3_X1   g083(.A1(new_n271), .A2(KEYINPUT82), .A3(new_n279), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT82), .ZN(new_n286));
  OAI211_X1 g085(.A(new_n286), .B(G22gat), .C1(new_n263), .C2(new_n270), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(new_n282), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n285), .A2(KEYINPUT83), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT83), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n287), .A2(new_n282), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n271), .A2(KEYINPUT82), .A3(new_n279), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n284), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(G183gat), .A2(G190gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT27), .B(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n300));
  AOI21_X1  g099(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(G169gat), .ZN(new_n302));
  INV_X1    g101(.A(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT26), .ZN(new_n305));
  NAND2_X1  g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT66), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(G169gat), .B2(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n308), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n305), .B(new_n306), .C1(new_n311), .C2(KEYINPUT26), .ZN(new_n312));
  XNOR2_X1  g111(.A(KEYINPUT68), .B(KEYINPUT28), .ZN(new_n313));
  OAI211_X1 g112(.A(new_n301), .B(new_n312), .C1(new_n299), .C2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(KEYINPUT23), .A3(new_n310), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT25), .ZN(new_n316));
  OR2_X1    g115(.A1(G183gat), .A2(G190gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(KEYINPUT24), .A3(new_n295), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT23), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n296), .A2(new_n321), .ZN(new_n322));
  NAND4_X1  g121(.A1(new_n318), .A2(new_n320), .A3(new_n322), .A4(new_n306), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n316), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(KEYINPUT67), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT65), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT25), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n307), .A2(KEYINPUT23), .ZN(new_n328));
  XNOR2_X1  g127(.A(new_n328), .B(KEYINPUT64), .ZN(new_n329));
  OAI211_X1 g128(.A(new_n326), .B(new_n327), .C1(new_n329), .C2(new_n323), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT67), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n331), .B1(new_n316), .B2(new_n323), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n325), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n327), .B1(new_n329), .B2(new_n323), .ZN(new_n334));
  AND2_X1   g133(.A1(new_n334), .A2(KEYINPUT65), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n314), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G113gat), .ZN(new_n337));
  INV_X1    g136(.A(G120gat), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT1), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n339), .B1(new_n337), .B2(new_n338), .ZN(new_n340));
  XNOR2_X1  g139(.A(G127gat), .B(G134gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n341), .A2(new_n342), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n340), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT70), .B(G120gat), .Z(new_n346));
  OAI211_X1 g145(.A(new_n339), .B(new_n341), .C1(new_n346), .C2(new_n337), .ZN(new_n347));
  AND2_X1   g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n336), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT65), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n350), .A2(new_n330), .A3(new_n325), .A4(new_n332), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n345), .A2(new_n347), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n314), .ZN(new_n353));
  AND2_X1   g152(.A1(new_n349), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(G227gat), .A2(G233gat), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT72), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT34), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  OAI211_X1 g157(.A(KEYINPUT72), .B(KEYINPUT34), .C1(new_n354), .C2(new_n355), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n349), .A2(new_n355), .A3(new_n353), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT32), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT33), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n361), .A2(new_n363), .ZN(new_n364));
  XOR2_X1   g163(.A(G15gat), .B(G43gat), .Z(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT71), .ZN(new_n366));
  XOR2_X1   g165(.A(G71gat), .B(G99gat), .Z(new_n367));
  XOR2_X1   g166(.A(new_n366), .B(new_n367), .Z(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(new_n364), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n361), .B(KEYINPUT32), .C1(new_n363), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g172(.A1(new_n358), .A2(new_n369), .A3(new_n359), .A4(new_n371), .ZN(new_n374));
  AOI21_X1  g173(.A(KEYINPUT73), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n358), .A2(new_n369), .A3(new_n359), .A4(new_n371), .ZN(new_n376));
  AND2_X1   g175(.A1(new_n376), .A2(KEYINPUT73), .ZN(new_n377));
  NOR2_X1   g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n258), .ZN(new_n379));
  NAND2_X1  g178(.A1(G226gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n336), .B2(new_n220), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n380), .B1(new_n351), .B2(new_n314), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n336), .A2(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT29), .B1(new_n351), .B2(new_n314), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n385), .B(new_n258), .C1(new_n386), .C2(new_n381), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  XNOR2_X1  g187(.A(G8gat), .B(G36gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(G64gat), .B(G92gat), .ZN(new_n390));
  XOR2_X1   g189(.A(new_n389), .B(new_n390), .Z(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n388), .A2(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n384), .A2(new_n387), .A3(new_n391), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(KEYINPUT30), .A3(new_n394), .ZN(new_n395));
  OR3_X1    g194(.A1(new_n388), .A2(KEYINPUT30), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G1gat), .B(G29gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT0), .ZN(new_n399));
  XNOR2_X1  g198(.A(G57gat), .B(G85gat), .ZN(new_n400));
  XNOR2_X1  g199(.A(new_n399), .B(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n348), .A2(KEYINPUT4), .A3(new_n259), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n259), .A2(new_n345), .A3(new_n347), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT4), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n259), .A2(new_n253), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n215), .A2(KEYINPUT3), .A3(new_n218), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n408), .A2(new_n352), .A3(new_n409), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n404), .A2(new_n407), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n219), .A2(new_n352), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT78), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(new_n405), .ZN(new_n414));
  INV_X1    g213(.A(new_n403), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n219), .A2(new_n352), .A3(KEYINPUT78), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI22_X1  g216(.A1(new_n403), .A2(new_n411), .B1(new_n417), .B2(KEYINPUT5), .ZN(new_n418));
  NAND4_X1  g217(.A1(new_n404), .A2(new_n407), .A3(new_n410), .A4(new_n403), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT5), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n402), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(KEYINPUT5), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n419), .ZN(new_n424));
  INV_X1    g223(.A(new_n421), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n401), .B(KEYINPUT86), .ZN(new_n426));
  INV_X1    g225(.A(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n424), .A2(new_n425), .A3(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT6), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n422), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n424), .A2(new_n425), .A3(KEYINPUT6), .A4(new_n401), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT35), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n378), .A2(new_n397), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n424), .A2(new_n425), .A3(new_n401), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n422), .A2(new_n434), .A3(new_n429), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(new_n431), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n397), .A2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n373), .A2(new_n374), .ZN(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n294), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI22_X1  g240(.A1(new_n294), .A2(new_n433), .B1(new_n441), .B2(KEYINPUT35), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n384), .A2(KEYINPUT88), .A3(new_n387), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT88), .ZN(new_n444));
  OAI211_X1 g243(.A(new_n444), .B(new_n379), .C1(new_n382), .C2(new_n383), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n443), .A2(KEYINPUT37), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT38), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n447), .B(new_n392), .C1(new_n388), .C2(KEYINPUT37), .ZN(new_n448));
  OAI21_X1  g247(.A(KEYINPUT89), .B1(new_n446), .B2(new_n448), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n392), .A2(KEYINPUT37), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n393), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT89), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n443), .A2(KEYINPUT37), .A3(new_n445), .ZN(new_n453));
  NAND4_X1  g252(.A1(new_n451), .A2(new_n452), .A3(new_n447), .A4(new_n453), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n388), .A2(KEYINPUT37), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n392), .B1(new_n388), .B2(KEYINPUT37), .ZN(new_n456));
  OAI21_X1  g255(.A(KEYINPUT38), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n430), .A2(new_n431), .A3(new_n394), .ZN(new_n458));
  NAND4_X1  g257(.A1(new_n449), .A2(new_n454), .A3(new_n457), .A4(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT40), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n410), .A2(new_n404), .A3(new_n407), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n415), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT39), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n415), .B1(new_n414), .B2(new_n416), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n426), .B1(new_n462), .B2(KEYINPUT39), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n460), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT87), .ZN(new_n468));
  XNOR2_X1  g267(.A(new_n467), .B(new_n468), .ZN(new_n469));
  OR3_X1    g268(.A1(new_n465), .A2(new_n460), .A3(new_n466), .ZN(new_n470));
  AND2_X1   g269(.A1(new_n470), .A2(new_n428), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n469), .A2(new_n471), .A3(new_n396), .A4(new_n395), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n459), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n284), .ZN(new_n474));
  OAI21_X1  g273(.A(KEYINPUT83), .B1(new_n285), .B2(new_n288), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n291), .A2(new_n290), .A3(new_n292), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n473), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n294), .A2(KEYINPUT84), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT84), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n437), .A3(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT36), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n375), .B2(new_n377), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n440), .A2(KEYINPUT36), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n482), .A2(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT85), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n478), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n482), .A2(KEYINPUT85), .A3(new_n486), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n442), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G15gat), .B(G22gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n492), .B(KEYINPUT92), .ZN(new_n493));
  INV_X1    g292(.A(G1gat), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n494), .A2(KEYINPUT16), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n492), .B(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n494), .ZN(new_n499));
  INV_X1    g298(.A(G8gat), .ZN(new_n500));
  AND3_X1   g299(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n500), .B1(new_n496), .B2(new_n499), .ZN(new_n502));
  NOR2_X1   g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g302(.A(G43gat), .B(G50gat), .ZN(new_n504));
  INV_X1    g303(.A(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT14), .ZN(new_n506));
  INV_X1    g305(.A(G29gat), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n509));
  AOI21_X1  g308(.A(G36gat), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(G36gat), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n506), .A2(new_n511), .A3(G29gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G50gat), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT91), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT15), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n505), .B1(new_n513), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n517), .ZN(new_n519));
  OAI211_X1 g318(.A(new_n519), .B(new_n504), .C1(new_n510), .C2(new_n512), .ZN(new_n520));
  OR3_X1    g319(.A1(new_n510), .A2(KEYINPUT15), .A3(new_n512), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n518), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT17), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n518), .A2(KEYINPUT17), .A3(new_n520), .A4(new_n521), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n503), .A2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(G229gat), .A2(G233gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n522), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n501), .B2(new_n502), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT93), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n532), .A2(KEYINPUT18), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n502), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n496), .A2(new_n499), .A3(new_n500), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n522), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(KEYINPUT94), .A3(new_n530), .ZN(new_n538));
  XOR2_X1   g337(.A(new_n528), .B(KEYINPUT13), .Z(new_n539));
  INV_X1    g338(.A(KEYINPUT94), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n503), .A2(new_n540), .A3(new_n522), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(new_n533), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n527), .A2(new_n528), .A3(new_n530), .A4(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n534), .A2(new_n542), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G113gat), .B(G141gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(KEYINPUT90), .B(KEYINPUT11), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n546), .B(new_n547), .ZN(new_n548));
  XOR2_X1   g347(.A(G169gat), .B(G197gat), .Z(new_n549));
  XNOR2_X1  g348(.A(new_n548), .B(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(KEYINPUT12), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n545), .A2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n534), .A2(new_n542), .A3(new_n544), .A4(new_n551), .ZN(new_n554));
  NAND3_X1  g353(.A1(new_n553), .A2(KEYINPUT95), .A3(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT95), .B1(new_n553), .B2(new_n554), .ZN(new_n557));
  NOR2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT21), .ZN(new_n559));
  XOR2_X1   g358(.A(G57gat), .B(G64gat), .Z(new_n560));
  INV_X1    g359(.A(KEYINPUT9), .ZN(new_n561));
  INV_X1    g360(.A(G71gat), .ZN(new_n562));
  INV_X1    g361(.A(G78gat), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  XOR2_X1   g364(.A(G71gat), .B(G78gat), .Z(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n503), .B1(new_n559), .B2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G183gat), .B(G211gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(G231gat), .ZN(new_n571));
  INV_X1    g370(.A(G233gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n567), .A2(new_n559), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n574), .B1(new_n567), .B2(new_n559), .ZN(new_n577));
  OAI21_X1  g376(.A(G127gat), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g377(.A(new_n577), .ZN(new_n579));
  INV_X1    g378(.A(G127gat), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(new_n575), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n570), .B1(new_n578), .B2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  XNOR2_X1  g382(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n584));
  INV_X1    g383(.A(G155gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n584), .B(new_n585), .ZN(new_n586));
  NAND3_X1  g385(.A1(new_n578), .A2(new_n581), .A3(new_n570), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n583), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  INV_X1    g388(.A(new_n587), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n589), .B1(new_n590), .B2(new_n582), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n568), .B1(new_n588), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n588), .A2(new_n591), .A3(new_n568), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  INV_X1    g396(.A(new_n595), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n592), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G134gat), .B(G162gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G99gat), .A2(G106gat), .ZN(new_n602));
  INV_X1    g401(.A(G85gat), .ZN(new_n603));
  INV_X1    g402(.A(G92gat), .ZN(new_n604));
  AOI22_X1  g403(.A1(KEYINPUT8), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n603), .B2(new_n604), .ZN(new_n607));
  NAND3_X1  g406(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n605), .A2(new_n607), .A3(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(G99gat), .B(G106gat), .Z(new_n610));
  OR2_X1    g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT98), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n609), .A2(new_n610), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  OR3_X1    g413(.A1(new_n609), .A2(new_n612), .A3(new_n610), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n526), .A2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n619));
  AND2_X1   g418(.A1(G232gat), .A2(G233gat), .ZN(new_n620));
  AOI22_X1  g419(.A1(new_n616), .A2(new_n529), .B1(KEYINPUT41), .B2(new_n620), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n618), .A2(new_n619), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n619), .B1(new_n618), .B2(new_n621), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n601), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n621), .ZN(new_n626));
  AOI21_X1  g425(.A(new_n616), .B1(new_n524), .B2(new_n525), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT99), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n601), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n622), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n620), .A2(KEYINPUT41), .ZN(new_n632));
  XNOR2_X1  g431(.A(G190gat), .B(G218gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n625), .A2(new_n634), .A3(new_n630), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n566), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n565), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n641), .A2(new_n611), .A3(new_n613), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n642), .B1(new_n616), .B2(new_n641), .ZN(new_n643));
  NAND2_X1  g442(.A1(G230gat), .A2(G233gat), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(G120gat), .B(G148gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G176gat), .B(G204gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n647), .B(new_n648), .Z(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT10), .ZN(new_n651));
  OAI211_X1 g450(.A(new_n642), .B(new_n651), .C1(new_n616), .C2(new_n641), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n616), .A2(KEYINPUT10), .A3(new_n641), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT100), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n645), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n652), .A2(KEYINPUT100), .A3(new_n653), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n650), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n654), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n646), .B1(new_n660), .B2(new_n645), .ZN(new_n661));
  INV_X1    g460(.A(new_n649), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n600), .A2(new_n639), .A3(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n491), .A2(new_n558), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n436), .B(KEYINPUT101), .Z(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G1gat), .ZN(G1324gat));
  INV_X1    g469(.A(new_n397), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  XOR2_X1   g471(.A(KEYINPUT16), .B(G8gat), .Z(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n672), .A2(new_n500), .ZN(new_n675));
  OAI21_X1  g474(.A(KEYINPUT42), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n673), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT42), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(G1325gat));
  INV_X1    g479(.A(G15gat), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n667), .A2(new_n681), .A3(new_n378), .ZN(new_n682));
  INV_X1    g481(.A(new_n486), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n667), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n682), .B1(new_n684), .B2(new_n681), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT102), .ZN(G1326gat));
  NAND2_X1  g485(.A1(new_n475), .A2(new_n476), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n480), .B1(new_n687), .B2(new_n284), .ZN(new_n688));
  AOI211_X1 g487(.A(KEYINPUT84), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n667), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(KEYINPUT43), .B(G22gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NOR2_X1   g492(.A1(new_n491), .A2(new_n558), .ZN(new_n694));
  NOR3_X1   g493(.A1(new_n600), .A2(new_n639), .A3(new_n664), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n507), .A3(new_n668), .A4(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  INV_X1    g496(.A(new_n442), .ZN(new_n698));
  AND2_X1   g497(.A1(new_n459), .A2(new_n472), .ZN(new_n699));
  AOI22_X1  g498(.A1(new_n699), .A2(new_n294), .B1(new_n485), .B2(new_n484), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n482), .A2(new_n700), .A3(KEYINPUT103), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n482), .B2(new_n700), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n698), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(KEYINPUT104), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT103), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n688), .A2(new_n689), .A3(new_n438), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n486), .B1(new_n477), .B2(new_n473), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n482), .A2(new_n700), .A3(KEYINPUT103), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT104), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n710), .A2(new_n711), .A3(new_n698), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n636), .A2(KEYINPUT105), .A3(new_n637), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(KEYINPUT105), .B1(new_n636), .B2(new_n637), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n716), .A2(KEYINPUT44), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n704), .A2(new_n712), .A3(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT44), .B1(new_n491), .B2(new_n639), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n600), .A2(new_n664), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n553), .A2(new_n554), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n668), .ZN(new_n726));
  OAI21_X1  g525(.A(G29gat), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n697), .A2(new_n727), .ZN(G1328gat));
  INV_X1    g527(.A(KEYINPUT106), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n723), .B1(new_n718), .B2(new_n719), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n511), .B1(new_n730), .B2(new_n671), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n489), .A2(new_n490), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n698), .ZN(new_n733));
  INV_X1    g532(.A(new_n557), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n555), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n397), .A2(G36gat), .ZN(new_n736));
  NAND4_X1  g535(.A1(new_n733), .A2(new_n735), .A3(new_n695), .A4(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT46), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n729), .B1(new_n731), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT46), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n737), .B(new_n740), .ZN(new_n741));
  AOI211_X1 g540(.A(new_n397), .B(new_n723), .C1(new_n718), .C2(new_n719), .ZN(new_n742));
  OAI211_X1 g541(.A(new_n741), .B(KEYINPUT106), .C1(new_n742), .C2(new_n511), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n739), .A2(new_n743), .ZN(G1329gat));
  NAND3_X1  g543(.A1(new_n730), .A2(G43gat), .A3(new_n683), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n694), .A2(new_n695), .ZN(new_n746));
  INV_X1    g545(.A(new_n378), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n514), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n745), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(KEYINPUT47), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT47), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n745), .A2(new_n751), .A3(new_n748), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n750), .A2(new_n752), .ZN(G1330gat));
  OAI21_X1  g552(.A(G50gat), .B1(new_n725), .B2(new_n294), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT48), .ZN(new_n755));
  INV_X1    g554(.A(new_n746), .ZN(new_n756));
  INV_X1    g555(.A(new_n690), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n757), .A2(G50gat), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n755), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n754), .A2(new_n759), .ZN(new_n760));
  NOR3_X1   g559(.A1(new_n746), .A2(G50gat), .A3(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n730), .A2(new_n690), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n761), .B1(new_n762), .B2(G50gat), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n760), .B1(KEYINPUT48), .B2(new_n763), .ZN(G1331gat));
  AND2_X1   g563(.A1(new_n704), .A2(new_n712), .ZN(new_n765));
  INV_X1    g564(.A(new_n600), .ZN(new_n766));
  NOR4_X1   g565(.A1(new_n766), .A2(new_n722), .A3(new_n638), .A4(new_n665), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n726), .ZN(new_n769));
  XNOR2_X1  g568(.A(KEYINPUT107), .B(G57gat), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1332gat));
  XNOR2_X1  g570(.A(new_n397), .B(KEYINPUT108), .ZN(new_n772));
  INV_X1    g571(.A(new_n772), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n773), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n765), .A2(new_n767), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT109), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT109), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n765), .A2(new_n777), .A3(new_n767), .A4(new_n774), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  OR2_X1    g578(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n776), .A2(new_n782), .A3(new_n778), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n781), .A2(new_n783), .ZN(G1333gat));
  OAI21_X1  g583(.A(G71gat), .B1(new_n768), .B2(new_n486), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n765), .A2(new_n562), .A3(new_n378), .A4(new_n767), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT50), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n785), .A2(KEYINPUT50), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(G1334gat));
  NOR2_X1   g590(.A1(new_n768), .A2(new_n757), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(new_n563), .ZN(G1335gat));
  NOR2_X1   g592(.A1(new_n600), .A2(new_n722), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(new_n664), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n795), .B1(new_n718), .B2(new_n719), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  OAI21_X1  g596(.A(G85gat), .B1(new_n797), .B2(new_n726), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n794), .A2(new_n638), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n710), .B2(new_n698), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT51), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n664), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n668), .A2(new_n603), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n798), .B1(new_n802), .B2(new_n803), .ZN(G1336gat));
  AOI21_X1  g603(.A(new_n442), .B1(new_n708), .B2(new_n709), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT110), .B1(new_n805), .B2(new_n799), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT51), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT110), .ZN(new_n808));
  INV_X1    g607(.A(new_n799), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n703), .A2(new_n808), .A3(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n806), .A2(new_n807), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g610(.A(KEYINPUT111), .B1(new_n800), .B2(KEYINPUT51), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR3_X1   g612(.A1(new_n773), .A2(G92gat), .A3(new_n665), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n806), .A2(KEYINPUT111), .A3(new_n810), .A4(new_n807), .ZN(new_n815));
  AND3_X1   g614(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n604), .B1(new_n796), .B2(new_n671), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT52), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(KEYINPUT52), .B1(new_n801), .B2(new_n814), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n796), .A2(new_n772), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(new_n820), .B2(new_n604), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n818), .A2(new_n821), .ZN(G1337gat));
  OAI21_X1  g621(.A(G99gat), .B1(new_n797), .B2(new_n486), .ZN(new_n823));
  OR2_X1    g622(.A1(new_n747), .A2(G99gat), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n823), .B1(new_n802), .B2(new_n824), .ZN(G1338gat));
  NOR3_X1   g624(.A1(new_n294), .A2(G106gat), .A3(new_n665), .ZN(new_n826));
  AND3_X1   g625(.A1(new_n813), .A2(new_n815), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(G106gat), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n796), .B2(new_n690), .ZN(new_n829));
  OAI21_X1  g628(.A(KEYINPUT53), .B1(new_n827), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(KEYINPUT53), .B1(new_n801), .B2(new_n826), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n796), .A2(new_n477), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(new_n828), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n830), .A2(new_n833), .ZN(G1339gat));
  INV_X1    g633(.A(new_n722), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n600), .A2(new_n835), .A3(new_n639), .A4(new_n665), .ZN(new_n836));
  INV_X1    g635(.A(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n539), .B1(new_n538), .B2(new_n541), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n528), .B1(new_n527), .B2(new_n530), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n550), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AND2_X1   g639(.A1(new_n840), .A2(new_n554), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n841), .A2(new_n664), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT54), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n654), .A2(new_n843), .A3(new_n644), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n844), .A2(new_n662), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n656), .A2(new_n657), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n652), .A2(new_n645), .A3(new_n653), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT54), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT55), .B(new_n846), .C1(new_n847), .C2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(KEYINPUT55), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n849), .B1(new_n656), .B2(new_n657), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n852), .B2(new_n845), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n850), .A2(new_n853), .A3(new_n659), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n842), .B1(new_n854), .B2(new_n835), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT112), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT112), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n857), .B(new_n842), .C1(new_n854), .C2(new_n835), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n856), .A2(new_n716), .A3(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT105), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n638), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n713), .ZN(new_n862));
  INV_X1    g661(.A(new_n854), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n862), .A2(new_n863), .A3(new_n841), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n859), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n837), .B1(new_n865), .B2(new_n766), .ZN(new_n866));
  INV_X1    g665(.A(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n477), .A2(new_n439), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n867), .A2(new_n868), .A3(new_n668), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n869), .A2(new_n772), .ZN(new_n870));
  AOI21_X1  g669(.A(G113gat), .B1(new_n870), .B2(new_n722), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n866), .A2(new_n690), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n872), .A2(new_n378), .A3(new_n668), .A4(new_n773), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n873), .A2(new_n337), .A3(new_n558), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n871), .A2(new_n874), .ZN(G1340gat));
  NAND3_X1  g674(.A1(new_n870), .A2(new_n346), .A3(new_n664), .ZN(new_n876));
  OAI21_X1  g675(.A(G120gat), .B1(new_n873), .B2(new_n665), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n876), .A2(new_n877), .ZN(G1341gat));
  NAND3_X1  g677(.A1(new_n870), .A2(new_n580), .A3(new_n600), .ZN(new_n879));
  OAI21_X1  g678(.A(G127gat), .B1(new_n873), .B2(new_n766), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT113), .Z(G1342gat));
  OAI21_X1  g681(.A(G134gat), .B1(new_n873), .B2(new_n639), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT114), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n397), .A2(new_n638), .ZN(new_n885));
  NOR3_X1   g684(.A1(new_n869), .A2(G134gat), .A3(new_n885), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT56), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n884), .A2(new_n887), .ZN(G1343gat));
  INV_X1    g687(.A(KEYINPUT58), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT118), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n890), .B1(new_n867), .B2(new_n668), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n600), .B1(new_n859), .B2(new_n864), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n890), .B(new_n668), .C1(new_n892), .C2(new_n837), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n893), .A2(new_n477), .A3(new_n486), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n558), .A2(G141gat), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  NOR4_X1   g695(.A1(new_n891), .A2(new_n894), .A3(new_n772), .A4(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT57), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n898), .B1(new_n866), .B2(new_n294), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT116), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n852), .A2(new_n845), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n658), .B1(new_n901), .B2(KEYINPUT55), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT115), .B(new_n851), .C1(new_n852), .C2(new_n845), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n853), .A2(new_n904), .ZN(new_n905));
  AND3_X1   g704(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  AOI22_X1  g705(.A1(new_n906), .A2(new_n735), .B1(new_n664), .B2(new_n841), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n864), .B1(new_n907), .B2(new_n638), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n837), .B1(new_n908), .B2(new_n766), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n479), .A2(KEYINPUT57), .A3(new_n481), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n900), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n902), .A2(new_n841), .A3(new_n853), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n912), .B1(new_n861), .B2(new_n713), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n902), .A2(new_n903), .A3(new_n905), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n842), .B1(new_n558), .B2(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n915), .B2(new_n639), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n836), .B1(new_n916), .B2(new_n600), .ZN(new_n917));
  NAND4_X1  g716(.A1(new_n917), .A2(KEYINPUT116), .A3(KEYINPUT57), .A4(new_n690), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n899), .A2(new_n911), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g718(.A1(new_n683), .A2(new_n726), .A3(new_n772), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n919), .A2(new_n722), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(G141gat), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n897), .B1(new_n922), .B2(KEYINPUT117), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT117), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n921), .A2(new_n924), .A3(G141gat), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n889), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n919), .A2(new_n920), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n735), .ZN(new_n928));
  AOI211_X1 g727(.A(KEYINPUT58), .B(new_n897), .C1(new_n928), .C2(G141gat), .ZN(new_n929));
  OAI21_X1  g728(.A(KEYINPUT119), .B1(new_n926), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(G141gat), .ZN(new_n932));
  INV_X1    g731(.A(new_n897), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n932), .A2(new_n889), .A3(new_n933), .ZN(new_n934));
  AND3_X1   g733(.A1(new_n921), .A2(new_n924), .A3(G141gat), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n924), .B1(new_n921), .B2(G141gat), .ZN(new_n936));
  NOR3_X1   g735(.A1(new_n935), .A2(new_n936), .A3(new_n897), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n931), .B(new_n934), .C1(new_n937), .C2(new_n889), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n930), .A2(new_n938), .ZN(G1344gat));
  NOR3_X1   g738(.A1(new_n891), .A2(new_n894), .A3(new_n772), .ZN(new_n940));
  INV_X1    g739(.A(G148gat), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(new_n941), .A3(new_n664), .ZN(new_n942));
  XNOR2_X1  g741(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n867), .A2(KEYINPUT57), .A3(new_n477), .ZN(new_n944));
  OR2_X1    g743(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n666), .A2(new_n735), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n915), .A2(new_n639), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n947), .B1(new_n639), .B2(new_n912), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n946), .B1(new_n948), .B2(new_n766), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n898), .B1(new_n949), .B2(new_n757), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n944), .A2(KEYINPUT121), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n945), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n664), .A3(new_n920), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n943), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  AOI211_X1 g753(.A(KEYINPUT59), .B(new_n941), .C1(new_n927), .C2(new_n664), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n942), .B1(new_n954), .B2(new_n955), .ZN(G1345gat));
  NAND3_X1  g755(.A1(new_n940), .A2(new_n585), .A3(new_n600), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n927), .A2(new_n600), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n585), .ZN(G1346gat));
  OR4_X1    g758(.A1(G162gat), .A2(new_n891), .A3(new_n894), .A4(new_n885), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n927), .A2(new_n862), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G162gat), .ZN(new_n963));
  NOR2_X1   g762(.A1(new_n961), .A2(KEYINPUT122), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1347gat));
  NOR2_X1   g764(.A1(new_n866), .A2(new_n668), .ZN(new_n966));
  AND3_X1   g765(.A1(new_n966), .A2(new_n868), .A3(new_n772), .ZN(new_n967));
  AOI21_X1  g766(.A(G169gat), .B1(new_n967), .B2(new_n722), .ZN(new_n968));
  NAND4_X1  g767(.A1(new_n872), .A2(new_n671), .A3(new_n378), .A4(new_n726), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n302), .A3(new_n558), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n968), .A2(new_n970), .ZN(G1348gat));
  AOI21_X1  g770(.A(G176gat), .B1(new_n967), .B2(new_n664), .ZN(new_n972));
  XNOR2_X1  g771(.A(new_n972), .B(KEYINPUT123), .ZN(new_n973));
  NOR3_X1   g772(.A1(new_n969), .A2(new_n303), .A3(new_n665), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n973), .A2(new_n974), .ZN(G1349gat));
  NAND3_X1  g774(.A1(new_n967), .A2(new_n297), .A3(new_n600), .ZN(new_n976));
  OAI21_X1  g775(.A(G183gat), .B1(new_n969), .B2(new_n766), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g778(.A(G190gat), .B1(new_n969), .B2(new_n639), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n980), .A2(new_n981), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(KEYINPUT61), .A3(new_n983), .ZN(new_n984));
  NAND3_X1  g783(.A1(new_n967), .A2(new_n298), .A3(new_n862), .ZN(new_n985));
  OAI211_X1 g784(.A(new_n984), .B(new_n985), .C1(KEYINPUT61), .C2(new_n983), .ZN(G1351gat));
  XNOR2_X1  g785(.A(KEYINPUT126), .B(G197gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n486), .A2(new_n671), .A3(new_n726), .ZN(new_n988));
  XOR2_X1   g787(.A(new_n988), .B(KEYINPUT127), .Z(new_n989));
  NAND2_X1  g788(.A1(new_n952), .A2(new_n989), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n987), .B1(new_n990), .B2(new_n558), .ZN(new_n991));
  NAND4_X1  g790(.A1(new_n966), .A2(new_n477), .A3(new_n486), .A4(new_n772), .ZN(new_n992));
  XNOR2_X1  g791(.A(new_n992), .B(KEYINPUT125), .ZN(new_n993));
  NOR2_X1   g792(.A1(new_n835), .A2(new_n987), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n991), .A2(new_n995), .ZN(G1352gat));
  OAI21_X1  g795(.A(G204gat), .B1(new_n990), .B2(new_n665), .ZN(new_n997));
  NOR3_X1   g796(.A1(new_n992), .A2(G204gat), .A3(new_n665), .ZN(new_n998));
  XNOR2_X1  g797(.A(new_n998), .B(KEYINPUT62), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n997), .A2(new_n999), .ZN(G1353gat));
  NAND3_X1  g799(.A1(new_n993), .A2(new_n225), .A3(new_n600), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n952), .A2(new_n600), .A3(new_n989), .ZN(new_n1002));
  AND3_X1   g801(.A1(new_n1002), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1003));
  AOI21_X1  g802(.A(KEYINPUT63), .B1(new_n1002), .B2(G211gat), .ZN(new_n1004));
  OAI21_X1  g803(.A(new_n1001), .B1(new_n1003), .B2(new_n1004), .ZN(G1354gat));
  OAI21_X1  g804(.A(G218gat), .B1(new_n990), .B2(new_n639), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n993), .A2(new_n226), .A3(new_n862), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n1006), .A2(new_n1007), .ZN(G1355gat));
endmodule


