//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n457, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n540, new_n541, new_n542,
    new_n543, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n554, new_n556, new_n557, new_n559, new_n560, new_n561,
    new_n562, new_n563, new_n564, new_n565, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n600, new_n601, new_n604,
    new_n605, new_n607, new_n608, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT66), .Z(G217));
  NOR4_X1   g025(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  AOI22_X1  g030(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n453), .ZN(G319));
  NAND2_X1  g031(.A1(G101), .A2(G2104), .ZN(new_n457));
  INV_X1    g032(.A(G2104), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n458), .A2(KEYINPUT3), .ZN(new_n459));
  INV_X1    g034(.A(KEYINPUT3), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G137), .ZN(new_n463));
  OAI21_X1  g038(.A(new_n457), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n462), .A2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n459), .A2(new_n461), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n468), .B1(new_n472), .B2(G125), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  AOI211_X1 g049(.A(KEYINPUT68), .B(new_n474), .C1(new_n469), .C2(new_n471), .ZN(new_n475));
  INV_X1    g050(.A(G113), .ZN(new_n476));
  OAI22_X1  g051(.A1(new_n473), .A2(new_n475), .B1(new_n476), .B2(new_n458), .ZN(new_n477));
  AOI21_X1  g052(.A(new_n467), .B1(new_n477), .B2(G2105), .ZN(G160));
  NOR2_X1   g053(.A1(new_n462), .A2(new_n465), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n462), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n465), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n480), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  AOI211_X1 g064(.A(KEYINPUT4), .B(new_n489), .C1(new_n469), .C2(new_n471), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(new_n459), .A3(new_n461), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT69), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n488), .A2(new_n459), .A3(new_n461), .A4(KEYINPUT69), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n493), .A2(KEYINPUT4), .A3(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT70), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n493), .A2(KEYINPUT70), .A3(KEYINPUT4), .A4(new_n494), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n490), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n459), .A2(new_n461), .A3(G126), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n465), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n458), .A2(G2105), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G102), .ZN(new_n504));
  INV_X1    g079(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(new_n506), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n499), .A2(new_n507), .ZN(G164));
  INV_X1    g083(.A(G50), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT71), .ZN(new_n512));
  XNOR2_X1  g087(.A(new_n511), .B(new_n512), .ZN(new_n513));
  OR2_X1    g088(.A1(new_n510), .A2(KEYINPUT6), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n513), .A2(G543), .A3(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT5), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT5), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G543), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n513), .A2(new_n521), .A3(new_n514), .ZN(new_n522));
  INV_X1    g097(.A(G88), .ZN(new_n523));
  OAI22_X1  g098(.A1(new_n509), .A2(new_n515), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n521), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n526), .A2(new_n510), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n525), .A2(new_n527), .ZN(G303));
  INV_X1    g103(.A(G303), .ZN(G166));
  INV_X1    g104(.A(new_n522), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(G89), .ZN(new_n531));
  INV_X1    g106(.A(new_n515), .ZN(new_n532));
  XNOR2_X1  g107(.A(KEYINPUT73), .B(G51), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n521), .A2(G63), .A3(G651), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  NAND4_X1  g112(.A1(new_n531), .A2(new_n534), .A3(new_n535), .A4(new_n537), .ZN(G286));
  INV_X1    g113(.A(G286), .ZN(G168));
  NAND2_X1  g114(.A1(new_n530), .A2(G90), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n532), .A2(G52), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n521), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  NAND3_X1  g118(.A1(new_n540), .A2(new_n541), .A3(new_n543), .ZN(G301));
  INV_X1    g119(.A(G301), .ZN(G171));
  NAND2_X1  g120(.A1(new_n530), .A2(G81), .ZN(new_n546));
  XNOR2_X1  g121(.A(KEYINPUT74), .B(G43), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n532), .A2(new_n547), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n521), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n549));
  OR2_X1    g124(.A1(new_n549), .A2(new_n510), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n546), .A2(new_n548), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  AND3_X1   g128(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G36), .ZN(G176));
  NAND2_X1  g130(.A1(G1), .A2(G3), .ZN(new_n556));
  XNOR2_X1  g131(.A(new_n556), .B(KEYINPUT8), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(G188));
  NAND4_X1  g133(.A1(new_n513), .A2(G53), .A3(G543), .A4(new_n514), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT9), .ZN(new_n560));
  INV_X1    g135(.A(G65), .ZN(new_n561));
  INV_X1    g136(.A(G78), .ZN(new_n562));
  OAI22_X1  g137(.A1(new_n520), .A2(new_n561), .B1(new_n562), .B2(new_n516), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(KEYINPUT75), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT75), .ZN(new_n565));
  OAI221_X1 g140(.A(new_n565), .B1(new_n562), .B2(new_n516), .C1(new_n520), .C2(new_n561), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n564), .A2(G651), .A3(new_n566), .ZN(new_n567));
  NAND4_X1  g142(.A1(new_n513), .A2(G91), .A3(new_n521), .A4(new_n514), .ZN(new_n568));
  AND2_X1   g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n560), .A2(new_n569), .ZN(G299));
  NAND2_X1  g145(.A1(new_n532), .A2(G49), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n530), .A2(G87), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n521), .B2(G74), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n521), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n510), .ZN(new_n576));
  AOI21_X1  g151(.A(new_n576), .B1(new_n530), .B2(G86), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n532), .A2(G48), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n577), .A2(new_n578), .ZN(G305));
  NAND2_X1  g154(.A1(new_n532), .A2(G47), .ZN(new_n580));
  XOR2_X1   g155(.A(KEYINPUT76), .B(G85), .Z(new_n581));
  NAND2_X1  g156(.A1(new_n530), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g157(.A1(new_n521), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n583));
  OAI211_X1 g158(.A(new_n580), .B(new_n582), .C1(new_n510), .C2(new_n583), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  INV_X1    g160(.A(G92), .ZN(new_n586));
  OR3_X1    g161(.A1(new_n522), .A2(KEYINPUT77), .A3(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT77), .B1(new_n522), .B2(new_n586), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n587), .A2(KEYINPUT10), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g164(.A(KEYINPUT10), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  INV_X1    g167(.A(G66), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n520), .B2(new_n593), .ZN(new_n594));
  AOI22_X1  g169(.A1(new_n532), .A2(G54), .B1(G651), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g171(.A(new_n596), .B(KEYINPUT78), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G284));
  OAI21_X1  g173(.A(new_n585), .B1(new_n597), .B2(G868), .ZN(G321));
  NAND2_X1  g174(.A1(G286), .A2(G868), .ZN(new_n600));
  INV_X1    g175(.A(G299), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G297));
  OAI21_X1  g177(.A(new_n600), .B1(new_n601), .B2(G868), .ZN(G280));
  INV_X1    g178(.A(G559), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n597), .B1(new_n604), .B2(G860), .ZN(new_n605));
  XOR2_X1   g180(.A(new_n605), .B(KEYINPUT79), .Z(G148));
  INV_X1    g181(.A(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n551), .A2(new_n607), .ZN(new_n608));
  AND2_X1   g183(.A1(new_n597), .A2(new_n604), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(new_n607), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT80), .Z(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g187(.A1(new_n472), .A2(new_n503), .ZN(new_n613));
  XNOR2_X1  g188(.A(KEYINPUT81), .B(KEYINPUT12), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n615), .B(new_n617), .ZN(new_n618));
  NOR2_X1   g193(.A1(KEYINPUT82), .A2(G2100), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n479), .A2(G123), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n481), .A2(G135), .ZN(new_n621));
  NOR2_X1   g196(.A1(G99), .A2(G2105), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(new_n465), .B2(G111), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  AOI21_X1  g199(.A(new_n619), .B1(new_n624), .B2(G2096), .ZN(new_n625));
  OAI211_X1 g200(.A(new_n618), .B(new_n625), .C1(G2096), .C2(new_n624), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2435), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT83), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XOR2_X1   g207(.A(G2451), .B(G2454), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n632), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G1341), .B(G1348), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XNOR2_X1  g212(.A(G2443), .B(G2446), .ZN(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n637), .B(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n640), .A2(G14), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2072), .B(G2078), .Z(new_n643));
  XOR2_X1   g218(.A(G2067), .B(G2678), .Z(new_n644));
  INV_X1    g219(.A(new_n644), .ZN(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g222(.A(new_n643), .B1(new_n647), .B2(KEYINPUT18), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(G2096), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2100), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n647), .A2(KEYINPUT17), .ZN(new_n651));
  OR2_X1    g226(.A1(new_n645), .A2(new_n646), .ZN(new_n652));
  AOI21_X1  g227(.A(KEYINPUT18), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(new_n650), .B(new_n653), .Z(G227));
  XNOR2_X1  g229(.A(G1971), .B(G1976), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT84), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT19), .Z(new_n657));
  XNOR2_X1  g232(.A(G1956), .B(G2474), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n657), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(new_n663), .B1(new_n657), .B2(new_n664), .ZN(new_n665));
  OR3_X1    g240(.A1(new_n657), .A2(new_n661), .A3(new_n664), .ZN(new_n666));
  OAI211_X1 g241(.A(new_n665), .B(new_n666), .C1(new_n663), .C2(new_n662), .ZN(new_n667));
  XOR2_X1   g242(.A(KEYINPUT21), .B(G1986), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(G1991), .B(G1996), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(KEYINPUT22), .B(G1981), .ZN(new_n672));
  XOR2_X1   g247(.A(new_n671), .B(new_n672), .Z(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(G229));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G35), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G162), .B2(new_n675), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT95), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT29), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2090), .ZN(new_n680));
  NAND2_X1  g255(.A1(G171), .A2(G16), .ZN(new_n681));
  OAI21_X1  g256(.A(new_n681), .B1(G5), .B2(G16), .ZN(new_n682));
  INV_X1    g257(.A(G1961), .ZN(new_n683));
  AND2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n685), .A2(G19), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(new_n552), .B2(new_n685), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1341), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G21), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(G168), .B2(G16), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n690), .A2(G1966), .ZN(new_n691));
  NOR4_X1   g266(.A1(new_n680), .A2(new_n684), .A3(new_n688), .A4(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n481), .A2(G141), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n479), .A2(G129), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n503), .A2(G105), .ZN(new_n695));
  NAND3_X1  g270(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT26), .Z(new_n697));
  NAND4_X1  g272(.A1(new_n693), .A2(new_n694), .A3(new_n695), .A4(new_n697), .ZN(new_n698));
  MUX2_X1   g273(.A(G32), .B(new_n698), .S(G29), .Z(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(new_n624), .A2(new_n675), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT31), .B(G11), .Z(new_n703));
  INV_X1    g278(.A(KEYINPUT30), .ZN(new_n704));
  OR2_X1    g279(.A1(new_n704), .A2(G28), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(G28), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n705), .A2(new_n706), .A3(new_n675), .ZN(new_n707));
  OAI21_X1  g282(.A(new_n707), .B1(new_n682), .B2(new_n683), .ZN(new_n708));
  OR2_X1    g283(.A1(G29), .A2(G33), .ZN(new_n709));
  AOI22_X1  g284(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n710));
  NOR2_X1   g285(.A1(new_n710), .A2(new_n465), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT90), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n481), .A2(G139), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n503), .A2(G103), .ZN(new_n714));
  XOR2_X1   g289(.A(new_n714), .B(KEYINPUT25), .Z(new_n715));
  NAND3_X1  g290(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(new_n709), .B1(new_n716), .B2(new_n675), .ZN(new_n717));
  INV_X1    g292(.A(G2072), .ZN(new_n718));
  AOI211_X1 g293(.A(new_n703), .B(new_n708), .C1(new_n717), .C2(new_n718), .ZN(new_n719));
  NAND4_X1  g294(.A1(new_n692), .A2(new_n701), .A3(new_n702), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT91), .B(KEYINPUT24), .ZN(new_n721));
  INV_X1    g296(.A(G34), .ZN(new_n722));
  AOI21_X1  g297(.A(G29), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(KEYINPUT92), .Z(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(new_n722), .B2(new_n721), .ZN(new_n725));
  INV_X1    g300(.A(G160), .ZN(new_n726));
  OAI21_X1  g301(.A(new_n725), .B1(new_n726), .B2(new_n675), .ZN(new_n727));
  INV_X1    g302(.A(G2084), .ZN(new_n728));
  AND2_X1   g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n690), .A2(G1966), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT94), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n675), .A2(G27), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G164), .B2(new_n675), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n731), .B1(G2078), .B2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n675), .A2(G26), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n479), .A2(G128), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n481), .A2(G140), .ZN(new_n737));
  OR2_X1    g312(.A1(G104), .A2(G2105), .ZN(new_n738));
  OAI211_X1 g313(.A(new_n738), .B(G2104), .C1(G116), .C2(new_n465), .ZN(new_n739));
  NAND3_X1  g314(.A1(new_n736), .A2(new_n737), .A3(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(KEYINPUT89), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n735), .B1(new_n743), .B2(new_n675), .ZN(new_n744));
  MUX2_X1   g319(.A(new_n735), .B(new_n744), .S(KEYINPUT28), .Z(new_n745));
  AND2_X1   g320(.A1(new_n745), .A2(G2067), .ZN(new_n746));
  NOR2_X1   g321(.A1(new_n745), .A2(G2067), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n717), .A2(new_n718), .ZN(new_n748));
  NOR3_X1   g323(.A1(new_n746), .A2(new_n747), .A3(new_n748), .ZN(new_n749));
  OR2_X1    g324(.A1(new_n733), .A2(G2078), .ZN(new_n750));
  NOR2_X1   g325(.A1(new_n727), .A2(new_n728), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT93), .ZN(new_n752));
  NAND4_X1  g327(.A1(new_n734), .A2(new_n749), .A3(new_n750), .A4(new_n752), .ZN(new_n753));
  NOR3_X1   g328(.A1(new_n720), .A2(new_n729), .A3(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G4), .A2(G16), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(new_n597), .B2(G16), .ZN(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT88), .B(G1348), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n685), .A2(KEYINPUT23), .A3(G20), .ZN(new_n759));
  INV_X1    g334(.A(KEYINPUT23), .ZN(new_n760));
  INV_X1    g335(.A(G20), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n760), .B1(new_n761), .B2(G16), .ZN(new_n762));
  OAI211_X1 g337(.A(new_n759), .B(new_n762), .C1(new_n601), .C2(new_n685), .ZN(new_n763));
  INV_X1    g338(.A(G1956), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n754), .A2(new_n758), .A3(new_n765), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT96), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n685), .A2(G22), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G166), .B2(new_n685), .ZN(new_n769));
  INV_X1    g344(.A(G1971), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n769), .B(new_n770), .ZN(new_n771));
  NOR2_X1   g346(.A1(G16), .A2(G23), .ZN(new_n772));
  INV_X1    g347(.A(G288), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n772), .B1(new_n773), .B2(G16), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT33), .B(G1976), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  MUX2_X1   g351(.A(G6), .B(G305), .S(G16), .Z(new_n777));
  XOR2_X1   g352(.A(KEYINPUT32), .B(G1981), .Z(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  NAND3_X1  g354(.A1(new_n771), .A2(new_n776), .A3(new_n779), .ZN(new_n780));
  XOR2_X1   g355(.A(new_n780), .B(KEYINPUT34), .Z(new_n781));
  NOR2_X1   g356(.A1(G16), .A2(G24), .ZN(new_n782));
  XOR2_X1   g357(.A(G290), .B(KEYINPUT87), .Z(new_n783));
  AOI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(G16), .ZN(new_n784));
  INV_X1    g359(.A(G1986), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  AOI22_X1  g361(.A1(G119), .A2(new_n479), .B1(new_n481), .B2(G131), .ZN(new_n787));
  OAI21_X1  g362(.A(G2104), .B1(new_n465), .B2(G107), .ZN(new_n788));
  NOR2_X1   g363(.A1(G95), .A2(G2105), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT86), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n787), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  MUX2_X1   g366(.A(G25), .B(new_n791), .S(G29), .Z(new_n792));
  XNOR2_X1  g367(.A(KEYINPUT35), .B(G1991), .ZN(new_n793));
  INV_X1    g368(.A(new_n793), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n792), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n781), .A2(new_n786), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT36), .Z(new_n797));
  NOR2_X1   g372(.A1(new_n767), .A2(new_n797), .ZN(G311));
  INV_X1    g373(.A(KEYINPUT96), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n766), .B(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n797), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(new_n801), .ZN(G150));
  NAND2_X1  g377(.A1(new_n530), .A2(G93), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n532), .A2(G55), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n521), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n805), .A2(new_n510), .ZN(new_n806));
  NAND3_X1  g381(.A1(new_n803), .A2(new_n804), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n807), .A2(G860), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT99), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT37), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n597), .A2(G559), .ZN(new_n811));
  XNOR2_X1  g386(.A(new_n811), .B(KEYINPUT39), .ZN(new_n812));
  INV_X1    g387(.A(new_n807), .ZN(new_n813));
  OR2_X1    g388(.A1(new_n551), .A2(KEYINPUT98), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n551), .A2(KEYINPUT98), .ZN(new_n815));
  AOI21_X1  g390(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n814), .A2(new_n813), .A3(new_n815), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n812), .B(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n810), .B1(new_n822), .B2(G860), .ZN(G145));
  XNOR2_X1  g398(.A(new_n742), .B(new_n698), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n497), .A2(new_n498), .ZN(new_n825));
  INV_X1    g400(.A(new_n490), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT100), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n828), .B1(new_n502), .B2(new_n505), .ZN(new_n829));
  INV_X1    g404(.A(new_n501), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT3), .B(G2104), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(G126), .ZN(new_n832));
  OAI211_X1 g407(.A(KEYINPUT100), .B(new_n504), .C1(new_n832), .C2(new_n465), .ZN(new_n833));
  AND2_X1   g408(.A1(new_n829), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n827), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n824), .B(new_n836), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n837), .B1(KEYINPUT101), .B2(new_n716), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n716), .B(KEYINPUT101), .ZN(new_n839));
  AOI21_X1  g414(.A(new_n838), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n615), .B(new_n791), .Z(new_n841));
  AND2_X1   g416(.A1(new_n479), .A2(G130), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n481), .A2(G142), .ZN(new_n844));
  OAI21_X1  g419(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n845));
  OR2_X1    g420(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n845), .A2(KEYINPUT103), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n846), .B(new_n847), .C1(G118), .C2(new_n465), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n842), .A2(KEYINPUT102), .ZN(new_n849));
  NAND4_X1  g424(.A1(new_n843), .A2(new_n844), .A3(new_n848), .A4(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n841), .B(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n840), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(G160), .B(new_n624), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G162), .ZN(new_n854));
  OR2_X1    g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G37), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n854), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g434(.A1(new_n807), .A2(new_n607), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n609), .B(new_n819), .ZN(new_n861));
  INV_X1    g436(.A(new_n596), .ZN(new_n862));
  INV_X1    g437(.A(KEYINPUT104), .ZN(new_n863));
  NAND2_X1  g438(.A1(G299), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n601), .A2(KEYINPUT104), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n596), .A2(new_n863), .A3(G299), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(KEYINPUT41), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n866), .A2(KEYINPUT41), .A3(new_n867), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n861), .A2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(new_n868), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n873), .B1(new_n874), .B2(new_n861), .ZN(new_n875));
  XNOR2_X1  g450(.A(G290), .B(G288), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(KEYINPUT105), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(G303), .B(G305), .ZN(new_n880));
  INV_X1    g455(.A(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n878), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT42), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n875), .B(new_n885), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n860), .B1(new_n886), .B2(new_n607), .ZN(G295));
  OAI21_X1  g462(.A(new_n860), .B1(new_n886), .B2(new_n607), .ZN(G331));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n889));
  INV_X1    g464(.A(KEYINPUT43), .ZN(new_n890));
  XNOR2_X1  g465(.A(G286), .B(G301), .ZN(new_n891));
  INV_X1    g466(.A(new_n818), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(new_n892), .B2(new_n816), .ZN(new_n893));
  INV_X1    g468(.A(new_n891), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n817), .A2(new_n894), .A3(new_n818), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT106), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n893), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n819), .A2(KEYINPUT106), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(new_n874), .ZN(new_n900));
  INV_X1    g475(.A(new_n884), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n895), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n870), .A2(new_n871), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n904), .A2(new_n856), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n900), .A2(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n884), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n890), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n904), .A2(new_n856), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n870), .A2(new_n871), .A3(new_n898), .A4(new_n897), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n874), .A2(new_n895), .A3(new_n893), .ZN(new_n911));
  AOI21_X1  g486(.A(new_n901), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g487(.A1(new_n909), .A2(KEYINPUT43), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n889), .B1(new_n908), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n914), .A2(KEYINPUT107), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT107), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n916), .B(new_n889), .C1(new_n908), .C2(new_n913), .ZN(new_n917));
  OAI21_X1  g492(.A(KEYINPUT43), .B1(new_n909), .B2(new_n912), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT108), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n905), .A2(new_n890), .A3(new_n907), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT108), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(KEYINPUT43), .C1(new_n909), .C2(new_n912), .ZN(new_n922));
  NAND4_X1  g497(.A1(new_n919), .A2(KEYINPUT44), .A3(new_n920), .A4(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n915), .A2(new_n917), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT109), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n915), .A2(KEYINPUT109), .A3(new_n917), .A4(new_n923), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(G397));
  XNOR2_X1  g503(.A(KEYINPUT110), .B(G1384), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n836), .A2(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT111), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n932));
  INV_X1    g507(.A(G40), .ZN(new_n933));
  AOI211_X1 g508(.A(new_n933), .B(new_n467), .C1(new_n477), .C2(G2105), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n932), .A3(new_n934), .ZN(new_n935));
  NOR3_X1   g510(.A1(new_n935), .A2(G1986), .A3(G290), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n935), .A2(new_n785), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(G290), .B2(new_n937), .ZN(new_n938));
  XNOR2_X1  g513(.A(new_n938), .B(KEYINPUT112), .ZN(new_n939));
  INV_X1    g514(.A(G2067), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n742), .B(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(G1996), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n698), .B(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n791), .B(new_n794), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n935), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g522(.A1(new_n939), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(G8), .ZN(new_n949));
  INV_X1    g524(.A(G1384), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n950), .B1(new_n499), .B2(new_n834), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n951), .A2(KEYINPUT113), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n953));
  OAI211_X1 g528(.A(new_n953), .B(new_n950), .C1(new_n499), .C2(new_n834), .ZN(new_n954));
  AOI21_X1  g529(.A(KEYINPUT50), .B1(new_n952), .B2(new_n954), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n950), .B1(new_n499), .B2(new_n507), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT50), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n934), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n955), .A2(new_n958), .A3(G2090), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n836), .A2(KEYINPUT45), .A3(new_n929), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n956), .A2(new_n932), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(new_n934), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n770), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n949), .B1(new_n959), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(G303), .A2(G8), .ZN(new_n965));
  XNOR2_X1  g540(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n965), .B(new_n966), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n964), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n968), .B(KEYINPUT115), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n952), .A2(new_n954), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n949), .B1(new_n971), .B2(new_n934), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n773), .A2(G1976), .ZN(new_n973));
  AND2_X1   g548(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g549(.A(KEYINPUT116), .B(G1976), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT52), .B1(G288), .B2(new_n975), .ZN(new_n976));
  AND2_X1   g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT52), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n974), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT49), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n972), .B1(KEYINPUT117), .B2(new_n980), .ZN(new_n981));
  NAND2_X1  g556(.A1(G305), .A2(G1981), .ZN(new_n982));
  INV_X1    g557(.A(G1981), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n577), .A2(new_n983), .A3(new_n578), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  AND2_X1   g560(.A1(new_n980), .A2(KEYINPUT117), .ZN(new_n986));
  XNOR2_X1  g561(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NOR2_X1   g562(.A1(new_n981), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n977), .A2(new_n979), .A3(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n952), .A2(KEYINPUT50), .A3(new_n954), .ZN(new_n990));
  INV_X1    g565(.A(new_n471), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n470), .B1(new_n459), .B2(new_n461), .ZN(new_n992));
  OAI21_X1  g567(.A(G125), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(KEYINPUT68), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n472), .A2(new_n468), .A3(G125), .ZN(new_n995));
  AOI22_X1  g570(.A1(new_n994), .A2(new_n995), .B1(G113), .B2(G2104), .ZN(new_n996));
  OAI211_X1 g571(.A(G40), .B(new_n466), .C1(new_n996), .C2(new_n465), .ZN(new_n997));
  AOI21_X1  g572(.A(G1384), .B1(new_n827), .B2(new_n506), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT50), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n990), .A2(new_n1000), .ZN(new_n1001));
  OR2_X1    g576(.A1(new_n1001), .A2(G2090), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n949), .B1(new_n1002), .B2(new_n963), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1003), .A2(new_n967), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n970), .A2(new_n989), .A3(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n952), .A2(new_n932), .A3(new_n954), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n997), .B1(new_n998), .B2(KEYINPUT45), .ZN(new_n1008));
  AOI21_X1  g583(.A(G1966), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n971), .A2(new_n999), .ZN(new_n1011));
  INV_X1    g586(.A(new_n958), .ZN(new_n1012));
  NAND3_X1  g587(.A1(new_n1011), .A2(new_n1012), .A3(new_n728), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT124), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n955), .A2(new_n958), .A3(G2084), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  NOR3_X1   g591(.A1(new_n1015), .A2(new_n1009), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(G286), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1015), .A2(new_n1009), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G168), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1020), .A2(new_n1021), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n949), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1010), .A2(new_n1013), .A3(KEYINPUT124), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1016), .B1(new_n1015), .B2(new_n1009), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(new_n1025), .A3(G168), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1021), .B1(new_n1026), .B2(G8), .ZN(new_n1027));
  OAI21_X1  g602(.A(KEYINPUT62), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1026), .A2(G8), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(KEYINPUT51), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT62), .ZN(new_n1031));
  AOI21_X1  g606(.A(G168), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1032));
  AOI21_X1  g607(.A(KEYINPUT51), .B1(new_n1019), .B2(G168), .ZN(new_n1033));
  OAI21_X1  g608(.A(G8), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1030), .A2(new_n1031), .A3(new_n1034), .ZN(new_n1035));
  AND3_X1   g610(.A1(new_n960), .A2(new_n934), .A3(new_n961), .ZN(new_n1036));
  INV_X1    g611(.A(G2078), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT53), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1961), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1037), .A2(KEYINPUT53), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n1040), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND4_X1  g618(.A1(new_n1028), .A2(new_n1035), .A3(G171), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1001), .A2(new_n764), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT56), .B(G2072), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1036), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT121), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n567), .A2(KEYINPUT120), .A3(new_n568), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n1048), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1049), .A2(new_n1048), .A3(new_n1050), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1052), .A2(new_n601), .A3(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1053), .ZN(new_n1055));
  OAI21_X1  g630(.A(G299), .B1(new_n1055), .B2(new_n1051), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1045), .A2(new_n1047), .A3(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1046), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n962), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g636(.A(G1956), .B1(new_n990), .B2(new_n1000), .ZN(new_n1062));
  NOR2_X1   g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1057), .A2(KEYINPUT122), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT122), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1054), .A2(new_n1056), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1063), .A2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(G1348), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(new_n955), .B2(new_n958), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n971), .A2(new_n940), .A3(new_n934), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n596), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n1059), .B1(new_n1068), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT61), .ZN(new_n1074));
  AOI21_X1  g649(.A(new_n1058), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1075));
  NOR3_X1   g650(.A1(new_n1061), .A2(new_n1062), .A3(new_n1057), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n1071), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1080), .A2(new_n862), .A3(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1059), .B(KEYINPUT61), .C1(new_n1067), .C2(new_n1063), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1077), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1036), .A2(new_n942), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n971), .A2(new_n934), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n551), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT59), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1090), .A2(KEYINPUT123), .ZN(new_n1091));
  OR2_X1    g666(.A1(new_n1090), .A2(KEYINPUT123), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1089), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1070), .A2(KEYINPUT60), .A3(new_n596), .A4(new_n1071), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1093), .B(new_n1094), .C1(new_n1091), .C2(new_n1089), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1073), .B1(new_n1084), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1097));
  XNOR2_X1  g672(.A(G301), .B(KEYINPUT54), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1043), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n931), .A2(new_n932), .ZN(new_n1100));
  NOR2_X1   g675(.A1(new_n467), .A2(new_n1042), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n465), .B1(new_n996), .B2(KEYINPUT125), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n933), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1100), .A2(new_n960), .A3(new_n1101), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1098), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1040), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g683(.A(new_n1006), .B1(new_n1044), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g684(.A1(new_n1020), .A2(G8), .A3(G168), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1004), .A2(new_n1110), .A3(KEYINPUT63), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n989), .B1(new_n969), .B2(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1110), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(new_n989), .C1(new_n964), .C2(new_n967), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT63), .ZN(new_n1115));
  NOR2_X1   g690(.A1(G288), .A2(G1976), .ZN(new_n1116));
  XNOR2_X1  g691(.A(new_n1116), .B(KEYINPUT118), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1117), .B1(new_n981), .B2(new_n987), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1118), .A2(new_n984), .ZN(new_n1119));
  OR2_X1    g694(.A1(new_n1119), .A2(KEYINPUT119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(KEYINPUT119), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n972), .A3(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1112), .A2(new_n1115), .A3(new_n1122), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n948), .B1(new_n1109), .B2(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g699(.A(new_n936), .B(KEYINPUT48), .ZN(new_n1125));
  NOR2_X1   g700(.A1(new_n1125), .A2(new_n947), .ZN(new_n1126));
  INV_X1    g701(.A(new_n935), .ZN(new_n1127));
  INV_X1    g702(.A(new_n941), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1127), .B1(new_n698), .B2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1127), .A2(KEYINPUT46), .A3(new_n942), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT46), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(new_n935), .B2(G1996), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1129), .A2(new_n1130), .A3(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT47), .Z(new_n1134));
  OR2_X1    g709(.A1(new_n791), .A2(new_n793), .ZN(new_n1135));
  OAI22_X1  g710(.A1(new_n944), .A2(new_n1135), .B1(G2067), .B2(new_n742), .ZN(new_n1136));
  AOI211_X1 g711(.A(new_n1126), .B(new_n1134), .C1(new_n1127), .C2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1124), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT126), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1124), .A2(KEYINPUT126), .A3(new_n1137), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1140), .A2(new_n1141), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g717(.A(new_n858), .ZN(new_n1144));
  INV_X1    g718(.A(G227), .ZN(new_n1145));
  NAND3_X1  g719(.A1(new_n641), .A2(G319), .A3(new_n1145), .ZN(new_n1146));
  INV_X1    g720(.A(KEYINPUT127), .ZN(new_n1147));
  XNOR2_X1  g721(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  NOR2_X1   g722(.A1(new_n908), .A2(new_n913), .ZN(new_n1149));
  NOR4_X1   g723(.A1(new_n1144), .A2(new_n1148), .A3(G229), .A4(new_n1149), .ZN(G308));
  INV_X1    g724(.A(G308), .ZN(G225));
endmodule


