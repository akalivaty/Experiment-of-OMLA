//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 1 0 0 0 1 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 1 0 1 0 1 0 1 1 1 1 0 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  XNOR2_X1  g000(.A(G110), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G227), .ZN(new_n189));
  XNOR2_X1  g003(.A(new_n187), .B(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G143), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  AND2_X1   g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  NOR2_X1   g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n194), .B1(new_n195), .B2(new_n196), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n193), .B1(new_n197), .B2(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  OAI211_X1 g013(.A(new_n199), .B(new_n194), .C1(new_n195), .C2(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT64), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(new_n191), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT64), .A2(G146), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(G143), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  AOI22_X1  g019(.A1(new_n198), .A2(new_n200), .B1(new_n205), .B2(G128), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT1), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n194), .A2(G146), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n204), .A2(new_n207), .A3(G128), .A4(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT68), .B1(new_n206), .B2(new_n210), .ZN(new_n211));
  NOR3_X1   g025(.A1(new_n195), .A2(new_n196), .A3(new_n194), .ZN(new_n212));
  OAI21_X1  g026(.A(G128), .B1(new_n212), .B2(new_n207), .ZN(new_n213));
  AOI21_X1  g027(.A(G143), .B1(new_n202), .B2(new_n203), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n192), .B1(new_n214), .B2(new_n199), .ZN(new_n215));
  INV_X1    g029(.A(new_n200), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n213), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT68), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n217), .A2(new_n218), .A3(new_n209), .ZN(new_n219));
  XNOR2_X1  g033(.A(G104), .B(G107), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT76), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G104), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT3), .B1(new_n223), .B2(G107), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n225));
  INV_X1    g039(.A(G107), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n225), .A2(new_n226), .A3(G104), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n223), .A2(G107), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n224), .A2(new_n227), .A3(new_n221), .A4(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT76), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n223), .A2(G107), .ZN(new_n231));
  NOR2_X1   g045(.A1(new_n226), .A2(G104), .ZN(new_n232));
  OAI211_X1 g046(.A(new_n230), .B(G101), .C1(new_n231), .C2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n222), .A2(new_n229), .A3(new_n233), .ZN(new_n234));
  NAND4_X1  g048(.A1(new_n211), .A2(new_n219), .A3(KEYINPUT10), .A4(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT66), .ZN(new_n236));
  XOR2_X1   g050(.A(KEYINPUT0), .B(G128), .Z(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n238), .B1(new_n198), .B2(new_n200), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n204), .A2(new_n208), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  OAI21_X1  g056(.A(new_n236), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT75), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n245), .A2(new_n246), .A3(KEYINPUT4), .A4(new_n229), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(KEYINPUT4), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n244), .A2(G101), .A3(new_n248), .ZN(new_n249));
  AND2_X1   g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n237), .B1(new_n215), .B2(new_n216), .ZN(new_n251));
  INV_X1    g065(.A(new_n242), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n251), .A2(KEYINPUT66), .A3(new_n252), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n243), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT11), .ZN(new_n255));
  INV_X1    g069(.A(G134), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n255), .B1(new_n256), .B2(G137), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(G137), .ZN(new_n258));
  INV_X1    g072(.A(G137), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT11), .A3(G134), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n257), .A2(new_n258), .A3(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  INV_X1    g076(.A(G131), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n257), .A2(new_n260), .A3(new_n263), .A4(new_n258), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT67), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n262), .A2(KEYINPUT67), .A3(new_n264), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n192), .A2(new_n271), .A3(KEYINPUT1), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(G128), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n271), .B1(new_n192), .B2(KEYINPUT1), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n240), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(new_n209), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n234), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT10), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n235), .A2(new_n254), .A3(new_n270), .A4(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT78), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n222), .A2(new_n229), .A3(new_n233), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n217), .A2(new_n209), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n277), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n269), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT79), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT12), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n286), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  AOI22_X1  g103(.A1(new_n284), .A2(new_n277), .B1(new_n268), .B2(new_n267), .ZN(new_n290));
  OAI21_X1  g104(.A(KEYINPUT79), .B1(new_n290), .B2(KEYINPUT12), .ZN(new_n291));
  INV_X1    g105(.A(new_n265), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n288), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n289), .A2(new_n291), .B1(new_n285), .B2(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n190), .B1(new_n282), .B2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n190), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n235), .A2(new_n254), .A3(new_n279), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(new_n269), .ZN(new_n298));
  AND2_X1   g112(.A1(new_n280), .A2(KEYINPUT78), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n280), .A2(KEYINPUT78), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n296), .B(new_n298), .C1(new_n299), .C2(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(G902), .B1(new_n295), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G469), .ZN(new_n303));
  OAI21_X1  g117(.A(KEYINPUT80), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n254), .A2(new_n279), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n305), .A2(new_n281), .A3(new_n270), .A4(new_n235), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n280), .A2(KEYINPUT78), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n306), .A2(new_n307), .B1(new_n269), .B2(new_n297), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT82), .B1(new_n308), .B2(new_n296), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n310));
  INV_X1    g124(.A(new_n298), .ZN(new_n311));
  OAI211_X1 g125(.A(new_n310), .B(new_n190), .C1(new_n282), .C2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(new_n294), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n313), .B(new_n296), .C1(new_n300), .C2(new_n299), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(new_n312), .A3(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  XOR2_X1   g130(.A(KEYINPUT81), .B(G469), .Z(new_n317));
  NAND3_X1  g131(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n289), .A2(new_n291), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n285), .A2(new_n293), .ZN(new_n320));
  AOI22_X1  g134(.A1(new_n306), .A2(new_n307), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n301), .B1(new_n321), .B2(new_n296), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(new_n316), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT80), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n323), .A2(new_n324), .A3(G469), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n304), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n194), .A2(G128), .ZN(new_n327));
  INV_X1    g141(.A(G128), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G143), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT88), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  XNOR2_X1  g146(.A(G128), .B(G143), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT88), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n256), .B1(new_n332), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n333), .A2(KEYINPUT13), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n336), .B(G134), .C1(KEYINPUT13), .C2(new_n327), .ZN(new_n337));
  INV_X1    g151(.A(G122), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G116), .ZN(new_n339));
  INV_X1    g153(.A(G116), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(G122), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  XNOR2_X1  g156(.A(KEYINPUT87), .B(G107), .ZN(new_n343));
  OR2_X1    g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n342), .A2(new_n343), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n335), .A2(new_n337), .A3(new_n344), .A4(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n330), .A2(new_n331), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n333), .A2(KEYINPUT88), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(G134), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n335), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n226), .B1(new_n339), .B2(KEYINPUT14), .ZN(new_n351));
  XOR2_X1   g165(.A(new_n351), .B(new_n342), .Z(new_n352));
  AND3_X1   g166(.A1(new_n350), .A2(KEYINPUT89), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT89), .B1(new_n350), .B2(new_n352), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n346), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  XNOR2_X1  g169(.A(KEYINPUT72), .B(G217), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n356), .A2(new_n357), .A3(G953), .ZN(new_n358));
  INV_X1    g172(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n355), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n346), .B(new_n358), .C1(new_n353), .C2(new_n354), .ZN(new_n361));
  AOI21_X1  g175(.A(G902), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(G478), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n363), .A2(KEYINPUT15), .ZN(new_n364));
  XNOR2_X1  g178(.A(new_n362), .B(new_n364), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT16), .ZN(new_n366));
  INV_X1    g180(.A(G125), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(G140), .ZN(new_n368));
  XNOR2_X1  g182(.A(G125), .B(G140), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT73), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(KEYINPUT73), .A3(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n368), .B1(new_n373), .B2(new_n366), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G146), .ZN(new_n375));
  INV_X1    g189(.A(G237), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n376), .A2(new_n188), .A3(G214), .ZN(new_n377));
  XNOR2_X1  g191(.A(new_n377), .B(new_n194), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G131), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n377), .B(G143), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(new_n263), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT17), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n191), .B(new_n368), .C1(new_n373), .C2(new_n366), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(KEYINPUT17), .A3(G131), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n375), .A2(new_n383), .A3(new_n384), .A4(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(G113), .B(G122), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n387), .B(new_n223), .ZN(new_n388));
  NAND2_X1  g202(.A1(KEYINPUT18), .A2(G131), .ZN(new_n389));
  XNOR2_X1  g203(.A(new_n378), .B(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n195), .A2(new_n196), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(new_n369), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n392), .B1(new_n373), .B2(new_n191), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n386), .A2(new_n388), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n374), .A2(G146), .B1(new_n379), .B2(new_n381), .ZN(new_n396));
  AND2_X1   g210(.A1(new_n373), .A2(KEYINPUT19), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n369), .A2(KEYINPUT19), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n391), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  AOI22_X1  g213(.A1(new_n396), .A2(new_n399), .B1(new_n393), .B2(new_n390), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n395), .B1(new_n388), .B2(new_n400), .ZN(new_n401));
  NOR2_X1   g215(.A1(G475), .A2(G902), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(KEYINPUT20), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT20), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n401), .A2(new_n405), .A3(new_n402), .ZN(new_n406));
  INV_X1    g220(.A(new_n395), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n388), .B1(new_n386), .B2(new_n394), .ZN(new_n408));
  OAI21_X1  g222(.A(new_n316), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n404), .A2(new_n406), .B1(G475), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n188), .A2(G952), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n411), .B1(G234), .B2(G237), .ZN(new_n412));
  NAND2_X1  g226(.A1(G234), .A2(G237), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n413), .A2(G902), .A3(G953), .ZN(new_n414));
  XNOR2_X1  g228(.A(KEYINPUT21), .B(G898), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n365), .A2(new_n410), .A3(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT84), .ZN(new_n420));
  XNOR2_X1  g234(.A(G116), .B(G119), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(KEYINPUT2), .B(G113), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n423), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n421), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n247), .A2(new_n427), .A3(new_n249), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n421), .A2(KEYINPUT5), .ZN(new_n429));
  NOR3_X1   g243(.A1(new_n340), .A2(KEYINPUT5), .A3(G119), .ZN(new_n430));
  INV_X1    g244(.A(G113), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AOI22_X1  g246(.A1(new_n429), .A2(new_n432), .B1(new_n425), .B2(new_n421), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n234), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n428), .A2(new_n434), .ZN(new_n435));
  XNOR2_X1  g249(.A(G110), .B(G122), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n435), .A2(KEYINPUT83), .A3(new_n437), .ZN(new_n438));
  OAI211_X1 g252(.A(new_n438), .B(KEYINPUT6), .C1(new_n435), .C2(new_n437), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n436), .B1(new_n428), .B2(new_n434), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n440), .A2(KEYINPUT83), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n420), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n198), .A2(new_n200), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n210), .B1(new_n443), .B2(new_n213), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n367), .ZN(new_n445));
  OAI21_X1  g259(.A(G125), .B1(new_n239), .B2(new_n242), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n188), .A2(G224), .ZN(new_n448));
  XOR2_X1   g262(.A(new_n448), .B(KEYINPUT85), .Z(new_n449));
  XNOR2_X1  g263(.A(new_n447), .B(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT6), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n440), .A2(new_n451), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n435), .A2(new_n437), .ZN(new_n453));
  NOR2_X1   g267(.A1(new_n453), .A2(new_n451), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n440), .A2(KEYINPUT83), .ZN(new_n455));
  NAND4_X1  g269(.A1(new_n454), .A2(new_n455), .A3(KEYINPUT84), .A4(new_n438), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n442), .A2(new_n450), .A3(new_n452), .A4(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT7), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n449), .A2(new_n458), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n447), .B(new_n459), .ZN(new_n460));
  XOR2_X1   g274(.A(new_n436), .B(KEYINPUT8), .Z(new_n461));
  OR2_X1    g275(.A1(new_n234), .A2(new_n433), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n461), .B1(new_n462), .B2(new_n434), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n453), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g278(.A(G902), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n457), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(G210), .B1(G237), .B2(G902), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT86), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n466), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n457), .A2(new_n469), .A3(new_n465), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G214), .B1(G237), .B2(G902), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n419), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(G221), .B1(new_n357), .B2(G902), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n476), .B(KEYINPUT74), .Z(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n326), .A2(new_n475), .A3(new_n478), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT90), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n258), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n256), .A2(G137), .ZN(new_n483));
  OAI21_X1  g297(.A(G131), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(new_n264), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n211), .A2(new_n219), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n243), .A2(new_n253), .A3(new_n269), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT30), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT30), .ZN(new_n490));
  NOR2_X1   g304(.A1(new_n444), .A2(new_n485), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n292), .A2(new_n239), .A3(new_n242), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n489), .A2(new_n427), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(new_n427), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n487), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n376), .A2(new_n188), .A3(G210), .ZN(new_n498));
  XOR2_X1   g312(.A(new_n498), .B(KEYINPUT27), .Z(new_n499));
  XNOR2_X1  g313(.A(KEYINPUT26), .B(G101), .ZN(new_n500));
  XOR2_X1   g314(.A(new_n499), .B(new_n500), .Z(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n497), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT29), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  AND3_X1   g319(.A1(new_n487), .A2(new_n488), .A3(new_n495), .ZN(new_n506));
  OAI21_X1  g320(.A(KEYINPUT70), .B1(new_n506), .B2(KEYINPUT28), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT70), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT28), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n496), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n427), .B1(new_n491), .B2(new_n492), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n496), .B2(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n507), .B(new_n510), .C1(new_n512), .C2(KEYINPUT69), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(KEYINPUT69), .ZN(new_n514));
  INV_X1    g328(.A(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI21_X1  g330(.A(new_n505), .B1(new_n516), .B2(new_n501), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT71), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n495), .B1(new_n487), .B2(new_n488), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT28), .B1(new_n506), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n520), .A2(new_n507), .A3(new_n510), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n502), .A2(new_n504), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n518), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  AND3_X1   g338(.A1(new_n496), .A2(new_n508), .A3(new_n509), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n508), .B1(new_n496), .B2(new_n509), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n527), .A2(KEYINPUT71), .A3(new_n520), .A4(new_n522), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n524), .A2(new_n316), .A3(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G472), .B1(new_n517), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT32), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n494), .A2(new_n501), .A3(new_n496), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT31), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT31), .ZN(new_n534));
  NAND4_X1  g348(.A1(new_n494), .A2(new_n534), .A3(new_n501), .A4(new_n496), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n533), .A2(new_n535), .ZN(new_n536));
  OR2_X1    g350(.A1(new_n512), .A2(KEYINPUT69), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n537), .A2(new_n527), .A3(new_n514), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n536), .B1(new_n502), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(G472), .A2(G902), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n531), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n502), .B1(new_n513), .B2(new_n515), .ZN(new_n543));
  AND2_X1   g357(.A1(new_n533), .A2(new_n535), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n545), .A2(KEYINPUT32), .A3(new_n540), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n530), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n356), .B1(G234), .B2(new_n316), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n375), .A2(new_n384), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT23), .ZN(new_n551));
  INV_X1    g365(.A(G119), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n551), .B1(new_n552), .B2(G128), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n328), .A2(KEYINPUT23), .A3(G119), .ZN(new_n554));
  OAI211_X1 g368(.A(new_n553), .B(new_n554), .C1(G119), .C2(new_n328), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT24), .B(G110), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  XNOR2_X1  g371(.A(G119), .B(G128), .ZN(new_n558));
  AOI22_X1  g372(.A1(new_n555), .A2(G110), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  OAI22_X1  g374(.A1(new_n555), .A2(G110), .B1(new_n557), .B2(new_n558), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n375), .A2(new_n392), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  XNOR2_X1  g377(.A(KEYINPUT22), .B(G137), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n564), .B(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n560), .A2(new_n562), .A3(new_n566), .ZN(new_n569));
  AND2_X1   g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(KEYINPUT25), .A3(new_n316), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n568), .A2(new_n316), .A3(new_n569), .ZN(new_n572));
  INV_X1    g386(.A(KEYINPUT25), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n549), .B1(new_n571), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n548), .A2(G902), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR2_X1   g392(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  AND2_X1   g393(.A1(new_n547), .A2(new_n579), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n326), .A2(new_n475), .A3(KEYINPUT90), .A4(new_n478), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n481), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT91), .B(G101), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n582), .B(new_n583), .ZN(G3));
  INV_X1    g398(.A(KEYINPUT92), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(G472), .C1(new_n539), .C2(G902), .ZN(new_n586));
  INV_X1    g400(.A(G472), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n587), .B1(new_n545), .B2(new_n316), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT92), .B1(new_n545), .B2(new_n540), .ZN(new_n589));
  OAI211_X1 g403(.A(new_n586), .B(new_n579), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n324), .B1(new_n323), .B2(G469), .ZN(new_n592));
  AOI211_X1 g406(.A(KEYINPUT80), .B(new_n303), .C1(new_n322), .C2(new_n316), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n477), .B1(new_n594), .B2(new_n318), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n591), .A2(new_n595), .A3(KEYINPUT93), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT93), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n326), .A2(new_n478), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n590), .ZN(new_n599));
  AND2_X1   g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n474), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n601), .B1(new_n466), .B2(new_n467), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n457), .A2(new_n465), .A3(new_n468), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n360), .A2(new_n361), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n605), .A2(KEYINPUT33), .ZN(new_n606));
  INV_X1    g420(.A(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n360), .A2(new_n607), .A3(new_n361), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT94), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n363), .A2(G902), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n609), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n404), .A2(new_n406), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n409), .A2(G475), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  AOI211_X1 g429(.A(new_n363), .B(G902), .C1(new_n606), .C2(new_n608), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT94), .B1(new_n362), .B2(G478), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n612), .B(new_n615), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n604), .A2(new_n416), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n600), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(KEYINPUT95), .ZN(new_n621));
  XNOR2_X1  g435(.A(KEYINPUT34), .B(G104), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NOR2_X1   g437(.A1(new_n615), .A2(new_n365), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR3_X1   g439(.A1(new_n604), .A2(new_n625), .A3(new_n416), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n600), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(KEYINPUT35), .B(G107), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G9));
  NOR2_X1   g443(.A1(new_n567), .A2(KEYINPUT36), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT96), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n563), .B(new_n631), .ZN(new_n632));
  AND2_X1   g446(.A1(new_n632), .A2(new_n576), .ZN(new_n633));
  NOR2_X1   g447(.A1(new_n575), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n586), .B(new_n635), .C1(new_n588), .C2(new_n589), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n481), .A2(new_n581), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT37), .B(G110), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G12));
  AOI21_X1  g454(.A(KEYINPUT32), .B1(new_n545), .B2(new_n540), .ZN(new_n641));
  AOI211_X1 g455(.A(new_n531), .B(new_n541), .C1(new_n543), .C2(new_n544), .ZN(new_n642));
  NOR2_X1   g456(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n634), .B1(new_n643), .B2(new_n530), .ZN(new_n644));
  AND2_X1   g458(.A1(new_n602), .A2(new_n603), .ZN(new_n645));
  INV_X1    g459(.A(new_n412), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT97), .B(G900), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n414), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g463(.A1(new_n645), .A2(KEYINPUT98), .A3(new_n624), .A4(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n602), .A2(new_n624), .A3(new_n603), .A4(new_n649), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT98), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n650), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n644), .A2(new_n595), .A3(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G128), .ZN(G30));
  XOR2_X1   g470(.A(new_n649), .B(KEYINPUT39), .Z(new_n657));
  OR2_X1    g471(.A1(new_n598), .A2(new_n657), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(KEYINPUT40), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n471), .A2(new_n472), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT99), .B(KEYINPUT38), .Z(new_n662));
  OR2_X1    g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n497), .A2(new_n501), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n506), .A2(new_n519), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n316), .B1(new_n669), .B2(new_n501), .ZN(new_n670));
  OAI21_X1  g484(.A(G472), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n643), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n365), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n615), .ZN(new_n674));
  NOR3_X1   g488(.A1(new_n635), .A2(new_n674), .A3(new_n601), .ZN(new_n675));
  AND3_X1   g489(.A1(new_n666), .A2(new_n672), .A3(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n659), .A2(new_n660), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G143), .ZN(G45));
  NOR2_X1   g492(.A1(new_n604), .A2(new_n618), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n644), .A2(new_n595), .A3(new_n679), .A4(new_n649), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT100), .B(G146), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G48));
  NAND2_X1  g496(.A1(new_n315), .A2(new_n316), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n683), .A2(G469), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n476), .A3(new_n318), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT101), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT101), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n684), .A2(new_n687), .A3(new_n476), .A4(new_n318), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n580), .A2(new_n686), .A3(new_n619), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND4_X1  g505(.A1(new_n580), .A2(new_n686), .A3(new_n626), .A4(new_n688), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G116), .ZN(G18));
  AND3_X1   g507(.A1(new_n684), .A2(new_n476), .A3(new_n318), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n644), .A2(new_n419), .A3(new_n645), .A4(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G119), .ZN(G21));
  OAI21_X1  g510(.A(G472), .B1(new_n539), .B2(G902), .ZN(new_n697));
  INV_X1    g511(.A(KEYINPUT102), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n521), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n527), .A2(KEYINPUT102), .A3(new_n520), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n699), .A2(new_n700), .A3(new_n502), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n540), .B1(new_n701), .B2(new_n536), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n697), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n579), .A2(KEYINPUT103), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT103), .ZN(new_n705));
  NOR3_X1   g519(.A1(new_n575), .A2(new_n578), .A3(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  NOR2_X1   g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  NOR3_X1   g522(.A1(new_n604), .A2(new_n416), .A3(new_n674), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n686), .A2(new_n708), .A3(new_n688), .A4(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  NAND4_X1  g525(.A1(new_n684), .A2(new_n645), .A3(new_n476), .A4(new_n318), .ZN(new_n712));
  INV_X1    g526(.A(new_n649), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n618), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n714), .A2(new_n697), .A3(new_n702), .A4(new_n635), .ZN(new_n715));
  NOR2_X1   g529(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n367), .ZN(G27));
  NAND2_X1  g531(.A1(new_n323), .A2(G469), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n318), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n719), .A2(new_n476), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT104), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n661), .A2(new_n474), .ZN(new_n723));
  INV_X1    g537(.A(new_n476), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n724), .B1(new_n318), .B2(new_n718), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n723), .B1(new_n725), .B2(KEYINPUT104), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n722), .A2(new_n726), .A3(new_n714), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT105), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n542), .B2(new_n546), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n641), .A2(KEYINPUT105), .ZN(new_n731));
  OAI21_X1  g545(.A(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT105), .B1(new_n641), .B2(new_n642), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n542), .A2(new_n729), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(KEYINPUT106), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n732), .A2(new_n735), .A3(new_n530), .ZN(new_n736));
  OR2_X1    g550(.A1(new_n704), .A2(new_n706), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n727), .A2(new_n736), .A3(KEYINPUT42), .A4(new_n737), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n580), .A2(new_n722), .A3(new_n726), .A4(new_n714), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT107), .B(G131), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G33));
  AND2_X1   g558(.A1(new_n722), .A2(new_n726), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n625), .A2(new_n713), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n745), .A2(KEYINPUT108), .A3(new_n580), .A4(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n580), .A2(new_n722), .A3(new_n726), .A4(new_n746), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT108), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n747), .A2(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  INV_X1    g566(.A(KEYINPUT45), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n322), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n295), .A2(KEYINPUT45), .A3(new_n301), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(G469), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(G469), .A2(G902), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n758), .A2(new_n318), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT109), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT109), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n758), .A2(new_n761), .A3(new_n318), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n756), .A2(new_n757), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n760), .B(new_n762), .C1(KEYINPUT46), .C2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n476), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n657), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n585), .B1(new_n539), .B2(new_n541), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n697), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(new_n586), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n609), .A2(new_n611), .ZN(new_n770));
  INV_X1    g584(.A(new_n617), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n410), .A3(new_n612), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT43), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT43), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n772), .A2(new_n775), .A3(new_n410), .A4(new_n612), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n774), .A2(new_n635), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n769), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT44), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n723), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(KEYINPUT110), .C1(new_n780), .C2(new_n779), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT110), .ZN(new_n783));
  INV_X1    g597(.A(new_n723), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n777), .B1(new_n768), .B2(new_n586), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(new_n785), .B2(KEYINPUT44), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n779), .A2(new_n780), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n766), .A2(new_n782), .A3(new_n788), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(G137), .ZN(G39));
  INV_X1    g604(.A(new_n714), .ZN(new_n791));
  NOR4_X1   g605(.A1(new_n547), .A2(new_n791), .A3(new_n723), .A4(new_n579), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n476), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT47), .B1(new_n764), .B2(new_n476), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n792), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT111), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT47), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n765), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(new_n793), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n800), .A2(new_n801), .A3(new_n792), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n797), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G140), .ZN(G42));
  INV_X1    g618(.A(new_n716), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n604), .A2(new_n674), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n635), .A2(new_n713), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n672), .A2(new_n806), .A3(new_n725), .A4(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n680), .A2(new_n655), .A3(new_n805), .A4(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT115), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  AND4_X1   g625(.A1(new_n547), .A2(new_n478), .A3(new_n326), .A4(new_n635), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n716), .B1(new_n812), .B2(new_n654), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n813), .A2(KEYINPUT115), .A3(new_n680), .A4(new_n808), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(KEYINPUT52), .B1(new_n811), .B2(new_n814), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND4_X1   g631(.A1(new_n689), .A2(new_n692), .A3(new_n695), .A4(new_n710), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n703), .A2(new_n634), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n547), .A2(new_n635), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n820), .A2(new_n598), .A3(new_n713), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n723), .A2(new_n673), .A3(new_n615), .ZN(new_n822));
  AOI22_X1  g636(.A1(new_n727), .A2(new_n819), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n742), .A2(new_n818), .A3(new_n751), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n618), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n417), .B1(new_n825), .B2(new_n624), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n826), .A2(new_n601), .A3(new_n661), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n596), .A2(new_n599), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT114), .ZN(new_n829));
  OAI211_X1 g643(.A(new_n481), .B(new_n581), .C1(new_n580), .C2(new_n637), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  AOI21_X1  g645(.A(new_n829), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(new_n824), .A2(new_n833), .ZN(new_n834));
  AND3_X1   g648(.A1(new_n817), .A2(new_n834), .A3(KEYINPUT53), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n809), .A2(KEYINPUT52), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n816), .A2(new_n836), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT53), .B1(new_n834), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g652(.A(KEYINPUT54), .B1(new_n835), .B2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT53), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n811), .A2(new_n814), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT52), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n814), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n828), .A2(new_n830), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT114), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n828), .A2(new_n830), .A3(new_n829), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n689), .A2(new_n692), .A3(new_n695), .A4(new_n710), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n821), .A2(new_n822), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n722), .A2(new_n726), .A3(new_n714), .A4(new_n819), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND4_X1  g668(.A1(new_n849), .A2(new_n742), .A3(new_n751), .A4(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n840), .B1(new_n845), .B2(new_n855), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n834), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n736), .A2(new_n737), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n774), .A2(new_n412), .A3(new_n776), .ZN(new_n861));
  AND3_X1   g675(.A1(new_n694), .A2(new_n784), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT48), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n860), .A2(KEYINPUT48), .A3(new_n862), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n411), .B(KEYINPUT118), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n697), .A2(new_n702), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n868), .A3(new_n737), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n869), .B2(new_n712), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n694), .A2(new_n784), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n643), .A2(new_n579), .A3(new_n412), .A4(new_n671), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n870), .B1(new_n825), .B2(new_n873), .ZN(new_n874));
  AND3_X1   g688(.A1(new_n865), .A2(new_n866), .A3(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n861), .A2(new_n868), .A3(new_n737), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n474), .B1(new_n663), .B2(new_n664), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n876), .A2(KEYINPUT50), .A3(new_n694), .A4(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT50), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n665), .A2(new_n694), .A3(new_n601), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n869), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n862), .A2(new_n819), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n772), .A2(new_n612), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n410), .ZN(new_n885));
  INV_X1    g699(.A(new_n885), .ZN(new_n886));
  AOI21_X1  g700(.A(KEYINPUT116), .B1(new_n873), .B2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n888));
  NOR4_X1   g702(.A1(new_n871), .A2(new_n872), .A3(new_n888), .A4(new_n885), .ZN(new_n889));
  OAI211_X1 g703(.A(new_n882), .B(new_n883), .C1(new_n887), .C2(new_n889), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n684), .A2(new_n318), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n891), .B(KEYINPUT113), .ZN(new_n892));
  OAI211_X1 g706(.A(new_n799), .B(new_n793), .C1(new_n478), .C2(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n869), .A2(new_n723), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n890), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g709(.A(new_n875), .B1(new_n895), .B2(KEYINPUT51), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n893), .A2(new_n894), .ZN(new_n897));
  INV_X1    g711(.A(new_n890), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n897), .A2(KEYINPUT51), .A3(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT117), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n895), .A2(KEYINPUT117), .A3(KEYINPUT51), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n896), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n839), .A2(new_n859), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT119), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT119), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n839), .A2(new_n903), .A3(new_n906), .A4(new_n859), .ZN(new_n907));
  OR2_X1    g721(.A1(G952), .A2(G953), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n905), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n892), .B(KEYINPUT49), .ZN(new_n910));
  NOR4_X1   g724(.A1(new_n707), .A2(new_n477), .A3(new_n601), .A4(new_n773), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n911), .B(KEYINPUT112), .ZN(new_n912));
  OR4_X1    g726(.A1(new_n672), .A2(new_n910), .A3(new_n666), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n913), .ZN(G75));
  NAND2_X1  g728(.A1(new_n856), .A2(new_n857), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n915), .A2(G210), .A3(G902), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n442), .A2(new_n452), .A3(new_n456), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n450), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT55), .Z(new_n919));
  XOR2_X1   g733(.A(KEYINPUT120), .B(KEYINPUT56), .Z(new_n920));
  NAND3_X1  g734(.A1(new_n916), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n188), .A2(G952), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT121), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT56), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n919), .B1(new_n916), .B2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n924), .A2(new_n926), .ZN(G51));
  XOR2_X1   g741(.A(new_n757), .B(KEYINPUT57), .Z(new_n928));
  INV_X1    g742(.A(new_n859), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n858), .B1(new_n856), .B2(new_n857), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n928), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n931), .A2(new_n315), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n915), .A2(G902), .ZN(new_n933));
  OR2_X1    g747(.A1(new_n933), .A2(new_n756), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n922), .B1(new_n932), .B2(new_n934), .ZN(G54));
  NAND2_X1  g749(.A1(KEYINPUT58), .A2(G475), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n937), .A2(new_n401), .ZN(new_n938));
  INV_X1    g752(.A(new_n401), .ZN(new_n939));
  NOR3_X1   g753(.A1(new_n933), .A2(new_n939), .A3(new_n936), .ZN(new_n940));
  NOR3_X1   g754(.A1(new_n938), .A2(new_n922), .A3(new_n940), .ZN(G60));
  NAND2_X1  g755(.A1(G478), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT59), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n609), .B(new_n943), .C1(new_n929), .C2(new_n930), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n944), .A2(new_n923), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n839), .A2(new_n859), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n609), .B1(new_n946), .B2(new_n943), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(G63));
  XOR2_X1   g762(.A(new_n570), .B(KEYINPUT122), .Z(new_n949));
  AND2_X1   g763(.A1(new_n856), .A2(new_n857), .ZN(new_n950));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT60), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n949), .B1(new_n950), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n923), .B1(KEYINPUT123), .B2(KEYINPUT61), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n952), .B1(new_n856), .B2(new_n857), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n955), .B2(new_n632), .ZN(new_n956));
  NAND2_X1  g770(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n957));
  AND3_X1   g771(.A1(new_n953), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n957), .B1(new_n953), .B2(new_n956), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n958), .A2(new_n959), .ZN(G66));
  INV_X1    g774(.A(new_n415), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n188), .B1(new_n961), .B2(G224), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n833), .A2(new_n850), .ZN(new_n963));
  INV_X1    g777(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n962), .B1(new_n964), .B2(new_n188), .ZN(new_n965));
  INV_X1    g779(.A(G898), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n917), .B1(new_n966), .B2(G953), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n965), .B(new_n967), .ZN(G69));
  INV_X1    g782(.A(KEYINPUT126), .ZN(new_n969));
  INV_X1    g783(.A(new_n789), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n797), .B2(new_n802), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n766), .A2(new_n806), .A3(new_n860), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n813), .A2(new_n680), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n972), .A2(new_n742), .A3(new_n751), .A4(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(G953), .B1(new_n971), .B2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n188), .A2(G900), .ZN(new_n977));
  OAI21_X1  g791(.A(new_n969), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n801), .B1(new_n800), .B2(new_n792), .ZN(new_n979));
  INV_X1    g793(.A(new_n792), .ZN(new_n980));
  AOI211_X1 g794(.A(KEYINPUT111), .B(new_n980), .C1(new_n799), .C2(new_n793), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n789), .B1(new_n979), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n188), .B1(new_n982), .B2(new_n974), .ZN(new_n983));
  INV_X1    g797(.A(new_n977), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(KEYINPUT126), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n489), .A2(new_n493), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT124), .Z(new_n987));
  NOR2_X1   g801(.A1(new_n397), .A2(new_n398), .ZN(new_n988));
  XOR2_X1   g802(.A(new_n987), .B(new_n988), .Z(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n978), .A2(new_n985), .A3(new_n990), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n580), .B(new_n784), .C1(new_n825), .C2(new_n624), .ZN(new_n992));
  NOR2_X1   g806(.A1(new_n992), .A2(new_n658), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n677), .A2(new_n973), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n993), .B1(new_n994), .B2(KEYINPUT62), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(KEYINPUT62), .ZN(new_n996));
  INV_X1    g810(.A(KEYINPUT125), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n994), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n188), .B1(new_n1000), .B2(new_n982), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1001), .A2(new_n989), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n991), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1004), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n991), .A2(new_n1006), .A3(new_n1002), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(G72));
  OR3_X1    g822(.A1(new_n1000), .A2(new_n964), .A3(new_n982), .ZN(new_n1009));
  XNOR2_X1  g823(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1010));
  NOR2_X1   g824(.A1(new_n587), .A2(new_n316), .ZN(new_n1011));
  XNOR2_X1  g825(.A(new_n1010), .B(new_n1011), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n667), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n835), .A2(new_n838), .ZN(new_n1014));
  NAND2_X1  g828(.A1(new_n503), .A2(new_n532), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1015), .A2(new_n1012), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g831(.A1(new_n971), .A2(new_n975), .A3(new_n963), .ZN(new_n1018));
  AOI211_X1 g832(.A(new_n501), .B(new_n497), .C1(new_n1018), .C2(new_n1012), .ZN(new_n1019));
  NOR4_X1   g833(.A1(new_n1013), .A2(new_n1017), .A3(new_n1019), .A4(new_n922), .ZN(G57));
endmodule


