//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 1 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:56 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1036, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1094, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1241, new_n1242, new_n1243, new_n1244;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NOR2_X1   g0002(.A1(G58), .A2(G68), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g0005(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n206));
  NAND3_X1  g0006(.A1(new_n205), .A2(G50), .A3(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NAND2_X1  g0008(.A1(G1), .A2(G13), .ZN(new_n209));
  NOR3_X1   g0009(.A1(new_n207), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(new_n208), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n213), .A2(G13), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  AOI22_X1  g0016(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n217));
  XOR2_X1   g0017(.A(new_n217), .B(KEYINPUT65), .Z(new_n218));
  NAND2_X1  g0018(.A1(G68), .A2(G238), .ZN(new_n219));
  INV_X1    g0019(.A(G50), .ZN(new_n220));
  INV_X1    g0020(.A(G226), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n219), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g0022(.A(new_n222), .B1(G77), .B2(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G58), .ZN(new_n224));
  INV_X1    g0024(.A(G232), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n218), .B(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  AOI21_X1  g0026(.A(new_n226), .B1(G116), .B2(G270), .ZN(new_n227));
  INV_X1    g0027(.A(G107), .ZN(new_n228));
  INV_X1    g0028(.A(G264), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(new_n213), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT66), .ZN(new_n232));
  OR2_X1    g0032(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(KEYINPUT1), .ZN(new_n234));
  AOI211_X1 g0034(.A(new_n210), .B(new_n216), .C1(new_n233), .C2(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(KEYINPUT2), .B(G226), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(new_n229), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(G270), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G68), .B(G77), .Z(new_n244));
  XNOR2_X1  g0044(.A(G50), .B(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(G87), .B(G97), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  AOI21_X1  g0050(.A(new_n208), .B1(new_n203), .B2(new_n220), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n251), .B1(G150), .B2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(KEYINPUT67), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(new_n224), .B2(KEYINPUT8), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  OAI21_X1  g0056(.A(new_n255), .B1(new_n256), .B2(new_n254), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n257), .B(KEYINPUT68), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(G33), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n253), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n212), .A2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n209), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  AOI22_X1  g0064(.A1(new_n260), .A2(new_n262), .B1(new_n220), .B2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n262), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n211), .A2(G20), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n266), .A2(G50), .A3(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n269), .B(KEYINPUT9), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT3), .ZN(new_n271));
  INV_X1    g0071(.A(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(KEYINPUT3), .A2(G33), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G222), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G223), .A2(G1698), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n209), .B1(G33), .B2(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(new_n279), .B(new_n280), .C1(G77), .C2(new_n275), .ZN(new_n281));
  OAI211_X1 g0081(.A(new_n211), .B(G274), .C1(G41), .C2(G45), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(G1), .A3(G13), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI211_X1 g0086(.A(new_n281), .B(new_n282), .C1(new_n221), .C2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G190), .ZN(new_n288));
  OR2_X1    g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n270), .A2(KEYINPUT72), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n287), .A2(G200), .ZN(new_n291));
  INV_X1    g0091(.A(new_n291), .ZN(new_n292));
  OR3_X1    g0092(.A1(new_n290), .A2(KEYINPUT10), .A3(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(KEYINPUT10), .B1(new_n290), .B2(new_n292), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n287), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n269), .B(new_n297), .C1(G179), .C2(new_n287), .ZN(new_n298));
  XOR2_X1   g0098(.A(new_n298), .B(KEYINPUT69), .Z(new_n299));
  INV_X1    g0099(.A(KEYINPUT13), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT73), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n284), .A2(new_n301), .A3(new_n285), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G238), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n301), .B1(new_n284), .B2(new_n285), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n282), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT74), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(KEYINPUT74), .B(new_n282), .C1(new_n303), .C2(new_n304), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n221), .A2(new_n276), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n275), .B(new_n310), .C1(G232), .C2(new_n276), .ZN(new_n311));
  NAND2_X1  g0111(.A1(G33), .A2(G97), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n284), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n300), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  AOI211_X1 g0115(.A(KEYINPUT13), .B(new_n313), .C1(new_n307), .C2(new_n308), .ZN(new_n316));
  NOR3_X1   g0116(.A1(new_n315), .A2(new_n316), .A3(new_n288), .ZN(new_n317));
  INV_X1    g0117(.A(G68), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT70), .ZN(new_n319));
  XNOR2_X1  g0119(.A(new_n263), .B(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(new_n262), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(new_n267), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n318), .B1(new_n322), .B2(KEYINPUT12), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT12), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n263), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n320), .A2(KEYINPUT12), .A3(new_n318), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n318), .A2(G20), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  INV_X1    g0128(.A(new_n252), .ZN(new_n329));
  OAI221_X1 g0129(.A(new_n327), .B1(new_n259), .B2(new_n328), .C1(new_n329), .C2(new_n220), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n262), .ZN(new_n331));
  XNOR2_X1  g0131(.A(new_n331), .B(KEYINPUT11), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n325), .A2(new_n326), .A3(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n317), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g0134(.A(G200), .B1(new_n315), .B2(new_n316), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AND2_X1   g0136(.A1(new_n299), .A2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n273), .A2(new_n208), .A3(new_n274), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n273), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n274), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n318), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n224), .A2(new_n318), .ZN(new_n343));
  OAI21_X1  g0143(.A(G20), .B1(new_n343), .B2(new_n203), .ZN(new_n344));
  INV_X1    g0144(.A(G159), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n344), .B1(new_n345), .B2(new_n329), .ZN(new_n346));
  OAI21_X1  g0146(.A(KEYINPUT76), .B1(new_n342), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(KEYINPUT16), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT16), .ZN(new_n349));
  OAI211_X1 g0149(.A(KEYINPUT76), .B(new_n349), .C1(new_n342), .C2(new_n346), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n348), .A2(new_n262), .A3(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(KEYINPUT68), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n257), .B(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n266), .A2(new_n267), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n355), .B1(new_n264), .B2(new_n353), .ZN(new_n356));
  AND2_X1   g0156(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT3), .A2(G33), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT3), .A2(G33), .ZN(new_n359));
  OAI211_X1 g0159(.A(G223), .B(new_n276), .C1(new_n358), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT77), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT77), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n275), .A2(new_n362), .A3(G223), .A4(new_n276), .ZN(new_n363));
  NAND2_X1  g0163(.A1(G33), .A2(G87), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n275), .A2(G226), .A3(G1698), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n361), .A2(new_n363), .A3(new_n364), .A4(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(new_n280), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n282), .B1(new_n286), .B2(new_n225), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT78), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI211_X1 g0170(.A(KEYINPUT78), .B(new_n282), .C1(new_n286), .C2(new_n225), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n367), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n367), .A2(new_n372), .A3(G190), .ZN(new_n375));
  NAND4_X1  g0175(.A1(new_n357), .A2(KEYINPUT17), .A3(new_n374), .A4(new_n375), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n351), .A2(new_n356), .A3(new_n374), .A4(new_n375), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT17), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n351), .A2(new_n356), .ZN(new_n380));
  AOI21_X1  g0180(.A(G169), .B1(new_n367), .B2(new_n372), .ZN(new_n381));
  INV_X1    g0181(.A(G179), .ZN(new_n382));
  AND2_X1   g0182(.A1(new_n367), .A2(new_n372), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n380), .A2(new_n384), .A3(KEYINPUT18), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT18), .B1(new_n380), .B2(new_n384), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n376), .B(new_n379), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n321), .A2(G77), .A3(new_n267), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n320), .A2(new_n328), .ZN(new_n389));
  NAND2_X1  g0189(.A1(G20), .A2(G77), .ZN(new_n390));
  XNOR2_X1  g0190(.A(KEYINPUT15), .B(G87), .ZN(new_n391));
  OAI221_X1 g0191(.A(new_n390), .B1(new_n256), .B2(new_n329), .C1(new_n259), .C2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n262), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n388), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  OR2_X1    g0194(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(KEYINPUT71), .ZN(new_n396));
  NAND2_X1  g0196(.A1(G238), .A2(G1698), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n275), .B(new_n397), .C1(new_n225), .C2(G1698), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n398), .B(new_n280), .C1(G107), .C2(new_n275), .ZN(new_n399));
  INV_X1    g0199(.A(G244), .ZN(new_n400));
  OAI211_X1 g0200(.A(new_n399), .B(new_n282), .C1(new_n400), .C2(new_n286), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n401), .A2(G200), .ZN(new_n402));
  OR2_X1    g0202(.A1(new_n401), .A2(new_n288), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n395), .A2(new_n396), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  OR2_X1    g0205(.A1(new_n401), .A2(G179), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n401), .A2(new_n296), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n406), .A2(new_n394), .A3(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n387), .A2(new_n405), .A3(new_n409), .ZN(new_n410));
  AND2_X1   g0210(.A1(KEYINPUT75), .A2(G169), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n411), .B1(new_n315), .B2(new_n316), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT14), .ZN(new_n413));
  OR3_X1    g0213(.A1(new_n315), .A2(new_n316), .A3(new_n382), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT14), .ZN(new_n415));
  OAI211_X1 g0215(.A(new_n415), .B(new_n411), .C1(new_n315), .C2(new_n316), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n413), .A2(new_n414), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n333), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n295), .A2(new_n337), .A3(new_n410), .A4(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(G116), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G283), .ZN(new_n422));
  INV_X1    g0222(.A(G97), .ZN(new_n423));
  OAI211_X1 g0223(.A(new_n422), .B(new_n208), .C1(G33), .C2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n262), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT20), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n262), .A2(KEYINPUT20), .A3(new_n421), .A4(new_n424), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n427), .A2(KEYINPUT86), .A3(new_n428), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n272), .A2(G1), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n420), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n321), .A2(new_n431), .B1(new_n420), .B2(new_n320), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT86), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n425), .A2(new_n433), .A3(new_n426), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n429), .A2(new_n432), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n358), .A2(new_n359), .ZN(new_n436));
  INV_X1    g0236(.A(G303), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n284), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(G264), .A2(G1698), .ZN(new_n439));
  INV_X1    g0239(.A(G257), .ZN(new_n440));
  OAI21_X1  g0240(.A(new_n439), .B1(new_n440), .B2(G1698), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n438), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT5), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G41), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n280), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(G41), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT81), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n211), .A4(G45), .ZN(new_n448));
  INV_X1    g0248(.A(G41), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n211), .B(G45), .C1(new_n449), .C2(KEYINPUT5), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(KEYINPUT81), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n445), .A2(G274), .A3(new_n448), .A4(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(G270), .B(new_n284), .C1(new_n450), .C2(new_n444), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n442), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n435), .A2(G169), .A3(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT21), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n454), .A2(G200), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n458), .B1(new_n288), .B2(new_n454), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n459), .A2(new_n435), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n454), .A2(KEYINPUT21), .A3(G169), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n461), .B1(new_n382), .B2(new_n454), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT87), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n462), .A2(new_n463), .A3(new_n435), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n463), .B1(new_n462), .B2(new_n435), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n457), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT4), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n468), .B1(new_n275), .B2(G250), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n469), .A2(new_n276), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n468), .A2(G1698), .ZN(new_n471));
  OAI211_X1 g0271(.A(new_n471), .B(G244), .C1(new_n359), .C2(new_n358), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n400), .B1(new_n273), .B2(new_n274), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n472), .B(new_n422), .C1(new_n473), .C2(KEYINPUT4), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n280), .B1(new_n470), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n450), .A2(new_n444), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(new_n280), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G257), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n452), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G200), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n288), .B2(new_n479), .ZN(new_n481));
  NOR3_X1   g0281(.A1(new_n262), .A2(new_n264), .A3(new_n430), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n483), .A2(new_n423), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n264), .A2(new_n423), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n486), .B(KEYINPUT80), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n252), .A2(G77), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n228), .A2(KEYINPUT6), .A3(G97), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT6), .ZN(new_n492));
  XNOR2_X1  g0292(.A(G97), .B(G107), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n489), .B1(new_n494), .B2(new_n208), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n228), .B1(new_n340), .B2(new_n341), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n262), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT79), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT7), .B1(new_n436), .B2(new_n208), .ZN(new_n500));
  INV_X1    g0300(.A(new_n341), .ZN(new_n501));
  OAI21_X1  g0301(.A(G107), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  AND2_X1   g0302(.A1(G97), .A2(G107), .ZN(new_n503));
  NOR2_X1   g0303(.A1(G97), .A2(G107), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n492), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n490), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT79), .B1(new_n508), .B2(new_n262), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n485), .B(new_n488), .C1(new_n499), .C2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n481), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n497), .A2(new_n498), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n508), .A2(KEYINPUT79), .A3(new_n262), .ZN(new_n513));
  AOI211_X1 g0313(.A(new_n487), .B(new_n484), .C1(new_n512), .C2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n479), .A2(new_n296), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n515), .B1(G179), .B2(new_n479), .ZN(new_n516));
  OAI21_X1  g0316(.A(KEYINPUT82), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(new_n452), .ZN(new_n518));
  OAI21_X1  g0318(.A(G244), .B1(new_n358), .B2(new_n359), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n468), .B1(G33), .B2(G283), .ZN(new_n520));
  OAI211_X1 g0320(.A(new_n520), .B(new_n472), .C1(new_n276), .C2(new_n469), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n518), .B1(new_n521), .B2(new_n280), .ZN(new_n522));
  AOI21_X1  g0322(.A(G169), .B1(new_n522), .B2(new_n478), .ZN(new_n523));
  AND4_X1   g0323(.A1(new_n382), .A2(new_n475), .A3(new_n452), .A4(new_n478), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT82), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(new_n526), .A3(new_n510), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n511), .B1(new_n517), .B2(new_n527), .ZN(new_n528));
  OAI211_X1 g0328(.A(new_n208), .B(G87), .C1(new_n358), .C2(new_n359), .ZN(new_n529));
  XNOR2_X1  g0329(.A(new_n529), .B(KEYINPUT22), .ZN(new_n530));
  NOR2_X1   g0330(.A1(new_n208), .A2(G107), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n531), .B(KEYINPUT23), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n272), .A2(new_n420), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n208), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n530), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(KEYINPUT24), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT24), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n530), .A2(new_n537), .A3(new_n532), .A4(new_n534), .ZN(new_n538));
  AOI21_X1  g0338(.A(new_n266), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AOI21_X1  g0339(.A(KEYINPUT25), .B1(new_n264), .B2(new_n228), .ZN(new_n540));
  AND3_X1   g0340(.A1(new_n264), .A2(KEYINPUT25), .A3(new_n228), .ZN(new_n541));
  OAI22_X1  g0341(.A1(new_n483), .A2(new_n228), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n440), .A2(G1698), .ZN(new_n544));
  OAI221_X1 g0344(.A(new_n544), .B1(G250), .B2(G1698), .C1(new_n358), .C2(new_n359), .ZN(new_n545));
  INV_X1    g0345(.A(G294), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n545), .B1(new_n272), .B2(new_n546), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n547), .A2(new_n280), .B1(new_n477), .B2(G264), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n452), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(G200), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n548), .A2(G190), .A3(new_n452), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n543), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n547), .A2(new_n280), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n477), .A2(G264), .ZN(new_n554));
  AND4_X1   g0354(.A1(new_n382), .A2(new_n553), .A3(new_n554), .A4(new_n452), .ZN(new_n555));
  AOI21_X1  g0355(.A(G169), .B1(new_n548), .B2(new_n452), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI21_X1  g0357(.A(new_n557), .B1(new_n539), .B2(new_n542), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n552), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n400), .A2(G1698), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n275), .B(new_n560), .C1(G238), .C2(G1698), .ZN(new_n561));
  INV_X1    g0361(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n280), .B1(new_n562), .B2(new_n533), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n211), .A2(G45), .ZN(new_n564));
  INV_X1    g0364(.A(G250), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(new_n566), .B(new_n284), .C1(G274), .C2(new_n564), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n568), .B2(new_n288), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n208), .B(G68), .C1(new_n358), .C2(new_n359), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT19), .ZN(new_n572));
  INV_X1    g0372(.A(G87), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n573), .A2(new_n423), .A3(new_n228), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n312), .A2(new_n208), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n572), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n259), .A2(KEYINPUT19), .A3(new_n423), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n571), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT83), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g0380(.A(KEYINPUT83), .B(new_n571), .C1(new_n576), .C2(new_n577), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n580), .A2(new_n262), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n320), .A2(new_n391), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n582), .B(new_n583), .C1(new_n573), .C2(new_n483), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n570), .A2(new_n584), .ZN(new_n585));
  XOR2_X1   g0385(.A(new_n391), .B(KEYINPUT84), .Z(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(new_n482), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n582), .A2(new_n587), .A3(new_n583), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT85), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n582), .A2(KEYINPUT85), .A3(new_n587), .A4(new_n583), .ZN(new_n591));
  AOI22_X1  g0391(.A1(new_n590), .A2(new_n591), .B1(new_n296), .B2(new_n568), .ZN(new_n592));
  INV_X1    g0392(.A(new_n568), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(new_n382), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n585), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n467), .A2(new_n528), .A3(new_n559), .A4(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n419), .A2(new_n596), .ZN(G372));
  INV_X1    g0397(.A(new_n299), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n336), .A2(new_n409), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n418), .ZN(new_n600));
  XNOR2_X1  g0400(.A(new_n377), .B(KEYINPUT17), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n380), .A2(new_n384), .ZN(new_n603));
  INV_X1    g0403(.A(KEYINPUT18), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n380), .A2(new_n384), .A3(KEYINPUT18), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n602), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n598), .B1(new_n295), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n590), .A2(new_n591), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n568), .A2(new_n296), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n610), .A2(new_n611), .A3(new_n594), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n570), .A2(new_n584), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n517), .A2(new_n527), .A3(new_n612), .A4(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(KEYINPUT26), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n517), .A2(new_n527), .ZN(new_n616));
  INV_X1    g0416(.A(new_n511), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n616), .A2(new_n617), .A3(new_n595), .ZN(new_n618));
  INV_X1    g0418(.A(KEYINPUT88), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n558), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g0420(.A1(new_n455), .A2(new_n456), .B1(new_n435), .B2(new_n462), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n557), .B(KEYINPUT88), .C1(new_n539), .C2(new_n542), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n620), .A2(new_n621), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n552), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n615), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT89), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n612), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n514), .A2(new_n516), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n595), .A2(new_n628), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n627), .B1(KEYINPUT26), .B2(new_n629), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n625), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n609), .B1(new_n419), .B2(new_n631), .ZN(G369));
  XOR2_X1   g0432(.A(new_n466), .B(KEYINPUT92), .Z(new_n633));
  NAND3_X1  g0433(.A1(new_n211), .A2(new_n208), .A3(G13), .ZN(new_n634));
  XNOR2_X1  g0434(.A(new_n634), .B(KEYINPUT90), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT27), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  XNOR2_X1  g0437(.A(new_n637), .B(KEYINPUT91), .ZN(new_n638));
  OR2_X1    g0438(.A1(new_n635), .A2(new_n636), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n639), .A2(G213), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(G343), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n435), .ZN(new_n644));
  MUX2_X1   g0444(.A(new_n621), .B(new_n633), .S(new_n644), .Z(new_n645));
  INV_X1    g0445(.A(G330), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n643), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n559), .B1(new_n543), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n558), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n650), .A2(new_n643), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n457), .B1(new_n464), .B2(new_n465), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n654), .A2(new_n648), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(new_n559), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n620), .A2(new_n622), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n648), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n653), .A2(new_n660), .ZN(G399));
  INV_X1    g0461(.A(new_n214), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(G41), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n574), .A2(G116), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G1), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n666), .B1(new_n207), .B2(new_n664), .ZN(new_n667));
  XNOR2_X1  g0467(.A(new_n667), .B(KEYINPUT28), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n648), .B1(new_n625), .B2(new_n630), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(KEYINPUT93), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT29), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT93), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n672), .B(new_n648), .C1(new_n625), .C2(new_n630), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(KEYINPUT94), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n552), .B1(new_n654), .B2(new_n650), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT82), .ZN(new_n677));
  AOI21_X1  g0477(.A(new_n526), .B1(new_n525), .B2(new_n510), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n617), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI22_X1  g0479(.A1(new_n676), .A2(new_n679), .B1(KEYINPUT26), .B2(new_n616), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n595), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n629), .A2(KEYINPUT26), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n682), .A2(new_n627), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n643), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT29), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT94), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n670), .A2(new_n686), .A3(new_n671), .A4(new_n673), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n675), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(KEYINPUT31), .B1(new_n596), .B2(new_n643), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n548), .A2(new_n563), .A3(new_n567), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n454), .A2(new_n382), .ZN(new_n691));
  NAND4_X1  g0491(.A1(new_n690), .A2(new_n478), .A3(new_n522), .A4(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT30), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n568), .A2(new_n454), .ZN(new_n694));
  NAND4_X1  g0494(.A1(new_n694), .A2(new_n382), .A3(new_n549), .A4(new_n479), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n648), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n689), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n696), .A2(KEYINPUT31), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n646), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n688), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n668), .B1(new_n703), .B2(G1), .ZN(G364));
  INV_X1    g0504(.A(new_n647), .ZN(new_n705));
  INV_X1    g0505(.A(G13), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(G20), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n707), .A2(G45), .ZN(new_n708));
  OR2_X1    g0508(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(KEYINPUT95), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n709), .A2(G1), .A3(new_n710), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n663), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n645), .A2(new_n646), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n705), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(new_n209), .B1(G20), .B2(new_n296), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n208), .A2(new_n288), .ZN(new_n718));
  INV_X1    g0518(.A(G200), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G179), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n718), .A2(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(G179), .A2(G200), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G190), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(G20), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n722), .A2(G303), .B1(new_n725), .B2(G294), .ZN(new_n726));
  INV_X1    g0526(.A(G322), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n382), .A2(G200), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n718), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n726), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n208), .A2(G190), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n723), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g0533(.A(new_n275), .B1(new_n733), .B2(G329), .ZN(new_n734));
  NOR3_X1   g0534(.A1(new_n208), .A2(new_n382), .A3(new_n719), .ZN(new_n735));
  XNOR2_X1  g0535(.A(new_n735), .B(KEYINPUT97), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n736), .A2(new_n288), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(G326), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n734), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n736), .A2(G190), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT33), .B(G317), .ZN(new_n742));
  AOI211_X1 g0542(.A(new_n730), .B(new_n740), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G283), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n731), .A2(new_n720), .ZN(new_n745));
  INV_X1    g0545(.A(G311), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n731), .A2(new_n728), .ZN(new_n747));
  OAI221_X1 g0547(.A(new_n743), .B1(new_n744), .B2(new_n745), .C1(new_n746), .C2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n733), .A2(G159), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT32), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(KEYINPUT98), .ZN(new_n751));
  INV_X1    g0551(.A(new_n741), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n318), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n721), .A2(new_n573), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n725), .A2(G97), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n755), .B1(new_n224), .B2(new_n729), .C1(new_n228), .C2(new_n745), .ZN(new_n756));
  OAI21_X1  g0556(.A(new_n275), .B1(new_n747), .B2(new_n328), .ZN(new_n757));
  NOR4_X1   g0557(.A1(new_n753), .A2(new_n754), .A3(new_n756), .A4(new_n757), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n758), .B1(KEYINPUT98), .B2(new_n750), .C1(new_n220), .C2(new_n738), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n717), .B1(new_n748), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G13), .A2(G33), .ZN(new_n761));
  XOR2_X1   g0561(.A(new_n761), .B(KEYINPUT96), .Z(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G20), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n645), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n214), .A2(G355), .A3(new_n275), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n662), .A2(new_n275), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G45), .B2(new_n207), .ZN(new_n768));
  INV_X1    g0568(.A(G45), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n246), .A2(new_n769), .ZN(new_n770));
  OAI221_X1 g0570(.A(new_n766), .B1(G116), .B2(new_n214), .C1(new_n768), .C2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n764), .A2(new_n716), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n765), .A2(new_n773), .A3(new_n712), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n715), .B1(new_n760), .B2(new_n774), .ZN(G396));
  INV_X1    g0575(.A(KEYINPUT100), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n408), .A2(new_n643), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n643), .A2(new_n394), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n404), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n776), .B(new_n778), .C1(new_n780), .C2(new_n409), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n409), .B1(new_n779), .B2(new_n404), .ZN(new_n782));
  OAI21_X1  g0582(.A(KEYINPUT100), .B1(new_n782), .B2(new_n777), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n670), .A2(new_n673), .A3(new_n785), .ZN(new_n786));
  OAI211_X1 g0586(.A(new_n648), .B(new_n784), .C1(new_n625), .C2(new_n630), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  OR3_X1    g0588(.A1(new_n786), .A2(new_n701), .A3(new_n788), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n701), .B1(new_n786), .B2(new_n788), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n789), .A2(new_n713), .A3(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n729), .ZN(new_n792));
  AOI22_X1  g0592(.A1(new_n741), .A2(G150), .B1(G143), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n345), .B2(new_n747), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n794), .B1(G137), .B2(new_n737), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT99), .ZN(new_n796));
  XNOR2_X1  g0596(.A(new_n796), .B(KEYINPUT34), .ZN(new_n797));
  INV_X1    g0597(.A(G132), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n797), .B(new_n275), .C1(new_n798), .C2(new_n732), .ZN(new_n799));
  INV_X1    g0599(.A(new_n745), .ZN(new_n800));
  AOI22_X1  g0600(.A1(G50), .A2(new_n722), .B1(new_n800), .B2(G68), .ZN(new_n801));
  INV_X1    g0601(.A(new_n725), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n801), .B1(new_n224), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n721), .A2(new_n228), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n800), .A2(G87), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n546), .B2(new_n729), .ZN(new_n806));
  OAI221_X1 g0606(.A(new_n755), .B1(new_n746), .B2(new_n732), .C1(new_n738), .C2(new_n437), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G283), .C2(new_n741), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n808), .B(new_n436), .C1(new_n420), .C2(new_n747), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n799), .A2(new_n803), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g0610(.A(new_n713), .B1(new_n810), .B2(new_n716), .ZN(new_n811));
  NOR2_X1   g0611(.A1(new_n716), .A2(new_n761), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI221_X1 g0613(.A(new_n811), .B1(G77), .B2(new_n813), .C1(new_n763), .C2(new_n784), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n791), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(G384));
  INV_X1    g0616(.A(KEYINPUT104), .ZN(new_n817));
  INV_X1    g0617(.A(new_n641), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n380), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n387), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n603), .A2(new_n819), .A3(new_n377), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n822), .A2(KEYINPUT37), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT37), .ZN(new_n824));
  NAND4_X1  g0624(.A1(new_n603), .A2(new_n819), .A3(new_n824), .A4(new_n377), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n821), .A2(KEYINPUT38), .A3(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT103), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  AOI21_X1  g0629(.A(KEYINPUT38), .B1(new_n821), .B2(new_n826), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g0631(.A(new_n828), .B(KEYINPUT38), .C1(new_n821), .C2(new_n826), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n817), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(new_n832), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n823), .A2(new_n825), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n819), .B1(new_n601), .B2(new_n607), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n828), .A3(new_n827), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n834), .A2(new_n839), .A3(KEYINPUT104), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT107), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n699), .B(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n785), .B1(new_n698), .B2(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT101), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n418), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n417), .A2(KEYINPUT101), .A3(new_n333), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n334), .A2(new_n335), .B1(new_n333), .B2(new_n643), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT102), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND3_X1   g0649(.A1(new_n417), .A2(KEYINPUT101), .A3(new_n333), .ZN(new_n850));
  AOI21_X1  g0650(.A(KEYINPUT101), .B1(new_n417), .B2(new_n333), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n848), .B(KEYINPUT102), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  OAI22_X1  g0653(.A1(new_n849), .A2(new_n853), .B1(new_n418), .B2(new_n648), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n833), .A2(new_n840), .A3(new_n843), .A4(new_n854), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT40), .ZN(new_n856));
  INV_X1    g0656(.A(new_n618), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n857), .A2(new_n559), .A3(new_n467), .A4(new_n648), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n696), .B1(new_n858), .B2(KEYINPUT31), .ZN(new_n859));
  XNOR2_X1  g0659(.A(new_n699), .B(KEYINPUT107), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n784), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n418), .A2(new_n648), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n848), .B1(new_n850), .B2(new_n851), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT102), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n862), .B1(new_n865), .B2(new_n852), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n861), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n838), .A2(KEYINPUT105), .A3(new_n827), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT105), .ZN(new_n869));
  NAND4_X1  g0669(.A1(new_n821), .A2(new_n869), .A3(new_n826), .A4(KEYINPUT38), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n871), .A2(new_n856), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n855), .A2(new_n856), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n419), .B1(new_n698), .B2(new_n842), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n873), .B(new_n874), .Z(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(G330), .ZN(new_n876));
  INV_X1    g0676(.A(new_n847), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n877), .A2(new_n648), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT39), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT106), .B1(new_n871), .B2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT106), .ZN(new_n881));
  AOI211_X1 g0681(.A(new_n881), .B(KEYINPUT39), .C1(new_n868), .C2(new_n870), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n834), .A2(new_n839), .A3(KEYINPUT39), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n878), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n787), .A2(new_n778), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n833), .A2(new_n840), .A3(new_n854), .A4(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n605), .A2(new_n606), .A3(new_n641), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n885), .A2(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n419), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n675), .A2(new_n891), .A3(new_n685), .A4(new_n687), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n892), .A2(new_n609), .ZN(new_n893));
  XNOR2_X1  g0693(.A(new_n890), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n876), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n895), .B1(new_n211), .B2(new_n707), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n420), .B1(new_n506), .B2(KEYINPUT35), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n209), .A2(new_n208), .ZN(new_n898));
  OAI211_X1 g0698(.A(new_n897), .B(new_n898), .C1(KEYINPUT35), .C2(new_n506), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n899), .B(KEYINPUT36), .ZN(new_n900));
  OAI21_X1  g0700(.A(G77), .B1(new_n224), .B2(new_n318), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n207), .A2(new_n901), .B1(G50), .B2(new_n318), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n902), .A2(G1), .A3(new_n706), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n896), .A2(new_n900), .A3(new_n903), .ZN(G367));
  OAI21_X1  g0704(.A(new_n528), .B1(new_n514), .B2(new_n648), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n628), .A2(new_n643), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(new_n559), .A3(new_n655), .ZN(new_n908));
  XNOR2_X1  g0708(.A(new_n908), .B(KEYINPUT42), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n907), .A2(new_n650), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n643), .B1(new_n910), .B2(new_n616), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n643), .A2(new_n584), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n595), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n627), .B2(new_n913), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(new_n907), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n653), .A2(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n917), .A2(new_n919), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n912), .B(new_n916), .C1(new_n653), .C2(new_n918), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n915), .A2(KEYINPUT43), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n922), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(KEYINPUT108), .B1(new_n918), .B2(new_n659), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT108), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n660), .A2(new_n927), .A3(new_n907), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT45), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n918), .A2(new_n659), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT44), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n932), .B(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n926), .A2(new_n928), .A3(KEYINPUT45), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AND2_X1   g0736(.A1(new_n647), .A2(new_n652), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND4_X1  g0738(.A1(new_n653), .A2(new_n934), .A3(new_n931), .A4(new_n935), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NOR2_X1   g0740(.A1(new_n652), .A2(new_n655), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT109), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n656), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(new_n705), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n703), .B1(new_n940), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n663), .B(KEYINPUT41), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n711), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n764), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n915), .A2(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n767), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n772), .B1(new_n214), .B2(new_n391), .C1(new_n242), .C2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n721), .A2(new_n420), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT46), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n752), .A2(new_n546), .B1(new_n802), .B2(new_n228), .ZN(new_n954));
  INV_X1    g0754(.A(new_n747), .ZN(new_n955));
  AOI211_X1 g0755(.A(new_n953), .B(new_n954), .C1(G283), .C2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n733), .A2(G317), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n737), .A2(G311), .ZN(new_n958));
  OAI22_X1  g0758(.A1(new_n729), .A2(new_n437), .B1(new_n745), .B2(new_n423), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n959), .A2(new_n275), .ZN(new_n960));
  NAND4_X1  g0760(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT110), .B(G137), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n963), .A2(new_n732), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n722), .A2(G58), .B1(new_n725), .B2(G68), .ZN(new_n965));
  INV_X1    g0765(.A(G150), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n965), .B1(new_n220), .B2(new_n747), .C1(new_n966), .C2(new_n729), .ZN(new_n967));
  AOI211_X1 g0767(.A(new_n964), .B(new_n967), .C1(G143), .C2(new_n737), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n800), .A2(G77), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n741), .A2(G159), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n968), .A2(new_n275), .A3(new_n969), .A4(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n961), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT47), .Z(new_n973));
  OAI211_X1 g0773(.A(new_n712), .B(new_n951), .C1(new_n973), .C2(new_n717), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n925), .A2(new_n947), .B1(new_n949), .B2(new_n974), .ZN(G387));
  XNOR2_X1  g0775(.A(new_n943), .B(new_n647), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n976), .A2(new_n711), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n741), .A2(G311), .B1(G317), .B2(new_n792), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n437), .B2(new_n747), .C1(new_n727), .C2(new_n738), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n979), .B(KEYINPUT48), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n980), .B1(new_n744), .B2(new_n802), .C1(new_n546), .C2(new_n721), .ZN(new_n981));
  XOR2_X1   g0781(.A(KEYINPUT112), .B(KEYINPUT49), .Z(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n436), .B1(new_n732), .B2(new_n739), .C1(new_n420), .C2(new_n745), .ZN(new_n984));
  INV_X1    g0784(.A(new_n586), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n985), .A2(new_n802), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n721), .A2(new_n328), .B1(new_n745), .B2(new_n423), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n436), .B(new_n987), .C1(G150), .C2(new_n733), .ZN(new_n988));
  OR2_X1    g0788(.A1(new_n988), .A2(KEYINPUT111), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(KEYINPUT111), .ZN(new_n990));
  OAI211_X1 g0790(.A(new_n989), .B(new_n990), .C1(new_n345), .C2(new_n738), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n353), .B2(new_n741), .ZN(new_n992));
  OAI221_X1 g0792(.A(new_n992), .B1(new_n220), .B2(new_n729), .C1(new_n318), .C2(new_n747), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n983), .A2(new_n984), .B1(new_n986), .B2(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n713), .B1(new_n994), .B2(new_n716), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n256), .A2(G50), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT50), .Z(new_n997));
  NOR2_X1   g0797(.A1(new_n318), .A2(new_n328), .ZN(new_n998));
  INV_X1    g0798(.A(new_n665), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n997), .A2(G45), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n767), .B1(new_n239), .B2(new_n769), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n999), .A2(new_n214), .A3(new_n275), .ZN(new_n1002));
  AOI21_X1  g0802(.A(new_n1000), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n214), .A2(G107), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n772), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n995), .B(new_n1005), .C1(new_n652), .C2(new_n948), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n663), .B1(new_n703), .B2(new_n976), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n944), .A2(new_n702), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n977), .B(new_n1006), .C1(new_n1007), .C2(new_n1008), .ZN(G393));
  NAND3_X1  g0809(.A1(new_n1008), .A2(new_n938), .A3(new_n939), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n938), .A2(KEYINPUT113), .A3(new_n939), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(KEYINPUT113), .B2(new_n939), .ZN(new_n1012));
  OAI211_X1 g0812(.A(new_n1010), .B(new_n663), .C1(new_n1012), .C2(new_n1008), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1012), .A2(new_n711), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n802), .A2(new_n328), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n737), .A2(G150), .B1(G159), .B2(new_n792), .ZN(new_n1016));
  XOR2_X1   g0816(.A(new_n1016), .B(KEYINPUT51), .Z(new_n1017));
  NAND2_X1  g0817(.A1(new_n733), .A2(G143), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n1018), .B1(new_n318), .B2(new_n721), .C1(new_n256), .C2(new_n747), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n275), .A3(new_n805), .A4(new_n1020), .ZN(new_n1021));
  AOI211_X1 g0821(.A(new_n1015), .B(new_n1021), .C1(G50), .C2(new_n741), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT115), .Z(new_n1023));
  AOI22_X1  g0823(.A1(new_n737), .A2(G317), .B1(G311), .B2(new_n792), .ZN(new_n1024));
  XOR2_X1   g0824(.A(new_n1024), .B(KEYINPUT52), .Z(new_n1025));
  AOI22_X1  g0825(.A1(G107), .A2(new_n800), .B1(new_n733), .B2(G322), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1025), .B(new_n1026), .C1(new_n546), .C2(new_n747), .ZN(new_n1027));
  AOI211_X1 g0827(.A(new_n275), .B(new_n1027), .C1(G116), .C2(new_n725), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1028), .B1(new_n744), .B2(new_n721), .C1(new_n437), .C2(new_n752), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n717), .B1(new_n1023), .B2(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n772), .B1(new_n423), .B2(new_n214), .C1(new_n249), .C2(new_n950), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT114), .ZN(new_n1032));
  NOR3_X1   g0832(.A1(new_n1030), .A2(new_n713), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n948), .B2(new_n907), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1013), .A2(new_n1014), .A3(new_n1034), .ZN(G390));
  AND2_X1   g0835(.A1(new_n868), .A2(new_n870), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n881), .B1(new_n1036), .B2(KEYINPUT39), .ZN(new_n1037));
  AND2_X1   g0837(.A1(new_n787), .A2(new_n778), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n878), .B1(new_n1038), .B2(new_n866), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n871), .A2(KEYINPUT106), .A3(new_n879), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1037), .A2(new_n1039), .A3(new_n884), .A4(new_n1040), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n854), .A2(new_n700), .A3(new_n784), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n777), .B1(new_n684), .B2(new_n784), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1036), .B(new_n878), .C1(new_n1044), .C2(new_n866), .ZN(new_n1045));
  AND3_X1   g0845(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n861), .A2(new_n646), .A3(new_n866), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1047), .B1(new_n1041), .B2(new_n1045), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n711), .B1(new_n1046), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(KEYINPUT116), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT116), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1051), .B(new_n711), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1050), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n874), .A2(G330), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n892), .A2(new_n609), .A3(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n854), .B1(new_n700), .B2(new_n784), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n886), .B1(new_n1047), .B2(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n866), .B1(new_n861), .B2(new_n646), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(new_n1044), .A3(new_n1042), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1048), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1041), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1062), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  OAI211_X1 g0865(.A(new_n1056), .B(new_n1061), .C1(new_n1046), .C2(new_n1048), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1065), .A2(new_n663), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(G128), .ZN(new_n1068));
  NOR2_X1   g0868(.A1(new_n738), .A2(new_n1068), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n752), .A2(new_n963), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n722), .A2(G150), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(new_n1071), .B(KEYINPUT53), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n802), .A2(new_n345), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1069), .A2(new_n1070), .A3(new_n1072), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n733), .A2(G125), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n800), .A2(G50), .ZN(new_n1076));
  XOR2_X1   g0876(.A(KEYINPUT54), .B(G143), .Z(new_n1077));
  INV_X1    g0877(.A(new_n1077), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n275), .B1(new_n1078), .B2(new_n747), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1079), .B1(G132), .B2(new_n792), .ZN(new_n1080));
  NAND4_X1  g0880(.A1(new_n1074), .A2(new_n1075), .A3(new_n1076), .A4(new_n1080), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n754), .B(new_n1015), .C1(new_n741), .C2(G107), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n955), .A2(G97), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n737), .A2(G283), .ZN(new_n1084));
  OAI22_X1  g0884(.A1(new_n729), .A2(new_n420), .B1(new_n745), .B2(new_n318), .ZN(new_n1085));
  AOI211_X1 g0885(.A(new_n275), .B(new_n1085), .C1(G294), .C2(new_n733), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n717), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n713), .B(new_n1088), .C1(new_n258), .C2(new_n812), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1037), .A2(new_n884), .A3(new_n1040), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n763), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1053), .A2(new_n1067), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g0892(.A(new_n1092), .ZN(G378));
  INV_X1    g0893(.A(KEYINPUT120), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n878), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1090), .A2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n889), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1094), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n855), .A2(new_n856), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n867), .A2(new_n872), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n269), .A2(new_n818), .ZN(new_n1101));
  XOR2_X1   g0901(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1102));
  XOR2_X1   g0902(.A(new_n1101), .B(new_n1102), .Z(new_n1103));
  AND3_X1   g0903(.A1(new_n295), .A2(new_n298), .A3(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1103), .B1(new_n295), .B2(new_n298), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT119), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  AND4_X1   g0906(.A1(G330), .A2(new_n1099), .A3(new_n1100), .A4(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n295), .A2(new_n298), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1103), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT119), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n295), .A2(new_n298), .A3(new_n1103), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1110), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1106), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1114), .B1(new_n873), .B2(G330), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1098), .B1(new_n1107), .B2(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(KEYINPUT120), .B1(new_n885), .B2(new_n889), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1099), .A2(G330), .A3(new_n1100), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1114), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n873), .A2(G330), .A3(new_n1106), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n1117), .A2(new_n1120), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n711), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n436), .B1(new_n721), .B2(new_n328), .C1(new_n802), .C2(new_n318), .ZN(new_n1125));
  AOI21_X1  g0925(.A(G41), .B1(new_n800), .B2(G58), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n1126), .B1(new_n744), .B2(new_n732), .C1(new_n738), .C2(new_n420), .ZN(new_n1127));
  AOI211_X1 g0927(.A(new_n1125), .B(new_n1127), .C1(G107), .C2(new_n792), .ZN(new_n1128));
  OAI221_X1 g0928(.A(new_n1128), .B1(new_n423), .B2(new_n752), .C1(new_n985), .C2(new_n747), .ZN(new_n1129));
  XOR2_X1   g0929(.A(KEYINPUT117), .B(KEYINPUT58), .Z(new_n1130));
  XNOR2_X1  g0930(.A(new_n1129), .B(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n220), .B1(new_n358), .B2(G41), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n802), .A2(new_n966), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(G128), .A2(new_n792), .B1(new_n955), .B2(G137), .ZN(new_n1134));
  OAI221_X1 g0934(.A(new_n1134), .B1(new_n721), .B2(new_n1078), .C1(new_n752), .C2(new_n798), .ZN(new_n1135));
  AOI211_X1 g0935(.A(new_n1133), .B(new_n1135), .C1(G125), .C2(new_n737), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT59), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(G33), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1139));
  AOI21_X1  g0939(.A(G41), .B1(new_n733), .B2(G124), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n345), .C2(new_n745), .ZN(new_n1141));
  OAI211_X1 g0941(.A(new_n1131), .B(new_n1132), .C1(new_n1138), .C2(new_n1141), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1142), .B(KEYINPUT118), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n713), .B1(new_n1143), .B2(new_n716), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n762), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(G50), .C2(new_n813), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1124), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1120), .A2(new_n890), .A3(new_n1121), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT121), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1107), .A2(new_n1115), .B1(new_n885), .B2(new_n889), .ZN(new_n1152));
  NAND4_X1  g0952(.A1(new_n1120), .A2(new_n890), .A3(KEYINPUT121), .A4(new_n1121), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1046), .A2(new_n1048), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1056), .B1(new_n1155), .B2(new_n1062), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1154), .A2(KEYINPUT57), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n1116), .A2(new_n1122), .B1(new_n1066), .B2(new_n1056), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n663), .B1(new_n1159), .B2(KEYINPUT57), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1148), .B1(new_n1158), .B2(new_n1160), .ZN(G375));
  NOR2_X1   g0961(.A1(new_n813), .A2(G68), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n969), .B1(new_n423), .B2(new_n721), .C1(new_n744), .C2(new_n729), .ZN(new_n1163));
  AOI211_X1 g0963(.A(new_n1163), .B(new_n986), .C1(G107), .C2(new_n955), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n275), .B1(new_n737), .B2(G294), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n1164), .B(new_n1165), .C1(new_n437), .C2(new_n732), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G116), .B2(new_n741), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n955), .A2(G150), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n275), .B1(new_n802), .B2(new_n220), .C1(new_n752), .C2(new_n1078), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n737), .A2(G132), .B1(G58), .B2(new_n800), .ZN(new_n1170));
  OAI221_X1 g0970(.A(new_n1170), .B1(new_n1068), .B2(new_n732), .C1(new_n345), .C2(new_n721), .ZN(new_n1171));
  AOI211_X1 g0971(.A(new_n1169), .B(new_n1171), .C1(new_n792), .C2(new_n962), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1167), .B1(new_n1168), .B2(new_n1172), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT124), .ZN(new_n1174));
  AOI211_X1 g0974(.A(new_n713), .B(new_n1162), .C1(new_n1174), .C2(new_n716), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n866), .A2(new_n761), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(new_n1176), .B(KEYINPUT123), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n1061), .A2(new_n711), .B1(new_n1175), .B2(new_n1177), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n946), .B(KEYINPUT122), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1062), .A2(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1056), .A2(new_n1061), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1178), .B1(new_n1180), .B2(new_n1181), .ZN(G381));
  OR2_X1    g0982(.A1(G387), .A2(G390), .ZN(new_n1183));
  OR2_X1    g0983(.A1(G381), .A2(G384), .ZN(new_n1184));
  NOR4_X1   g0984(.A1(new_n1183), .A2(G396), .A3(G393), .A4(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1123), .A2(new_n1156), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT57), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n664), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1147), .B1(new_n1188), .B2(new_n1157), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1185), .A2(new_n1092), .A3(new_n1189), .ZN(G407));
  NOR2_X1   g0990(.A1(new_n1185), .A2(new_n642), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1189), .A2(new_n1092), .ZN(new_n1192));
  OAI21_X1  g0992(.A(G213), .B1(new_n1191), .B2(new_n1192), .ZN(G409));
  XNOR2_X1  g0993(.A(G393), .B(G396), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(G387), .A2(G390), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1183), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1194), .ZN(new_n1197));
  AND2_X1   g0997(.A1(G387), .A2(G390), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(G387), .A2(G390), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1197), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT61), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1196), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT126), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n642), .A2(G213), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1154), .A2(new_n711), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1159), .A2(new_n1179), .ZN(new_n1206));
  NAND4_X1  g1006(.A1(new_n1092), .A2(new_n1146), .A3(new_n1205), .A4(new_n1206), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1204), .B(new_n1207), .C1(new_n1189), .C2(new_n1092), .ZN(new_n1208));
  INV_X1    g1008(.A(KEYINPUT60), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1210));
  NAND4_X1  g1010(.A1(new_n1055), .A2(KEYINPUT60), .A3(new_n1058), .A4(new_n1060), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1210), .A2(new_n663), .A3(new_n1062), .A4(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1212), .A2(new_n1178), .ZN(new_n1213));
  OR2_X1    g1013(.A1(new_n815), .A2(KEYINPUT125), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n815), .A2(KEYINPUT125), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(KEYINPUT125), .A3(new_n815), .A4(new_n1178), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NOR2_X1   g1019(.A1(new_n1208), .A2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1220), .A2(KEYINPUT63), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n642), .A2(G213), .A3(G2897), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1218), .A2(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1216), .A2(new_n1222), .A3(new_n1217), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1208), .A2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1227), .A2(KEYINPUT63), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1203), .B(new_n1221), .C1(new_n1228), .C2(new_n1220), .ZN(new_n1229));
  AOI22_X1  g1029(.A1(G375), .A2(G378), .B1(G213), .B2(new_n642), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT62), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1207), .A4(new_n1218), .ZN(new_n1232));
  OAI21_X1  g1032(.A(KEYINPUT62), .B1(new_n1208), .B2(new_n1219), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1234));
  AOI21_X1  g1034(.A(KEYINPUT127), .B1(new_n1227), .B2(new_n1201), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT127), .ZN(new_n1236));
  AOI211_X1 g1036(.A(new_n1236), .B(KEYINPUT61), .C1(new_n1208), .C2(new_n1226), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(new_n1234), .A2(new_n1235), .A3(new_n1237), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n1196), .A2(new_n1200), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1229), .B1(new_n1238), .B2(new_n1239), .ZN(G405));
  XNOR2_X1  g1040(.A(new_n1239), .B(new_n1219), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(G375), .A2(G378), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(new_n1192), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1241), .B(new_n1244), .ZN(G402));
endmodule


