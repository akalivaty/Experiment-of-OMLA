

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U550 ( .A1(n763), .A2(n745), .ZN(n750) );
  OR2_X2 U551 ( .A1(n762), .A2(n748), .ZN(n745) );
  XNOR2_X1 U552 ( .A(n530), .B(KEYINPUT78), .ZN(G164) );
  NAND2_X2 U553 ( .A1(G8), .A2(n727), .ZN(n726) );
  NAND2_X1 U554 ( .A1(n727), .A2(G1348), .ZN(n681) );
  NOR2_X1 U555 ( .A1(n679), .A2(n678), .ZN(n700) );
  XNOR2_X1 U556 ( .A(KEYINPUT27), .B(KEYINPUT88), .ZN(n676) );
  INV_X1 U557 ( .A(KEYINPUT33), .ZN(n754) );
  NAND2_X1 U558 ( .A1(n525), .A2(n524), .ZN(n527) );
  XNOR2_X1 U559 ( .A(n523), .B(n522), .ZN(n616) );
  XNOR2_X1 U560 ( .A(n521), .B(KEYINPUT64), .ZN(n522) );
  INV_X1 U561 ( .A(KEYINPUT23), .ZN(n531) );
  AND2_X1 U562 ( .A1(n760), .A2(n759), .ZN(n517) );
  XNOR2_X1 U563 ( .A(KEYINPUT95), .B(KEYINPUT96), .ZN(n518) );
  XOR2_X1 U564 ( .A(n701), .B(KEYINPUT28), .Z(n519) );
  AND2_X1 U565 ( .A1(G126), .A2(n897), .ZN(n520) );
  INV_X1 U566 ( .A(KEYINPUT91), .ZN(n680) );
  INV_X1 U567 ( .A(KEYINPUT92), .ZN(n684) );
  XNOR2_X1 U568 ( .A(n685), .B(n684), .ZN(n693) );
  INV_X1 U569 ( .A(n727), .ZN(n704) );
  NOR2_X1 U570 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U571 ( .A(n714), .B(KEYINPUT93), .ZN(n715) );
  XNOR2_X1 U572 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X1 U573 ( .A1(n710), .A2(n709), .ZN(n723) );
  XNOR2_X1 U574 ( .A(n735), .B(n518), .ZN(n737) );
  INV_X1 U575 ( .A(n986), .ZN(n759) );
  INV_X1 U576 ( .A(KEYINPUT17), .ZN(n521) );
  NOR2_X1 U577 ( .A1(G164), .A2(G1384), .ZN(n778) );
  NOR2_X1 U578 ( .A1(G651), .A2(G543), .ZN(n645) );
  XNOR2_X1 U579 ( .A(n532), .B(n531), .ZN(n534) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n523) );
  NAND2_X1 U581 ( .A1(n616), .A2(G138), .ZN(n529) );
  AND2_X2 U582 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U583 ( .A1(G114), .A2(n898), .ZN(n525) );
  INV_X2 U584 ( .A(G2105), .ZN(n526) );
  AND2_X4 U585 ( .A1(n526), .A2(G2104), .ZN(n893) );
  NAND2_X1 U586 ( .A1(G102), .A2(n893), .ZN(n524) );
  NOR2_X4 U587 ( .A1(G2104), .A2(n526), .ZN(n897) );
  NOR2_X1 U588 ( .A1(n527), .A2(n520), .ZN(n528) );
  AND2_X1 U589 ( .A1(n529), .A2(n528), .ZN(n530) );
  NAND2_X1 U590 ( .A1(G101), .A2(n893), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n898), .A2(G113), .ZN(n533) );
  NAND2_X1 U592 ( .A1(n534), .A2(n533), .ZN(n538) );
  NAND2_X1 U593 ( .A1(G137), .A2(n616), .ZN(n536) );
  NAND2_X1 U594 ( .A1(G125), .A2(n897), .ZN(n535) );
  NAND2_X1 U595 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X2 U596 ( .A1(n538), .A2(n537), .ZN(G160) );
  INV_X1 U597 ( .A(G651), .ZN(n542) );
  NOR2_X1 U598 ( .A1(G543), .A2(n542), .ZN(n539) );
  XOR2_X1 U599 ( .A(KEYINPUT1), .B(n539), .Z(n637) );
  NAND2_X1 U600 ( .A1(G60), .A2(n637), .ZN(n541) );
  XOR2_X1 U601 ( .A(KEYINPUT0), .B(G543), .Z(n634) );
  NOR2_X2 U602 ( .A1(G651), .A2(n634), .ZN(n638) );
  NAND2_X1 U603 ( .A1(G47), .A2(n638), .ZN(n540) );
  NAND2_X1 U604 ( .A1(n541), .A2(n540), .ZN(n546) );
  NAND2_X1 U605 ( .A1(G85), .A2(n645), .ZN(n544) );
  NOR2_X1 U606 ( .A1(n634), .A2(n542), .ZN(n641) );
  NAND2_X1 U607 ( .A1(G72), .A2(n641), .ZN(n543) );
  NAND2_X1 U608 ( .A1(n544), .A2(n543), .ZN(n545) );
  OR2_X1 U609 ( .A1(n546), .A2(n545), .ZN(G290) );
  AND2_X1 U610 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U611 ( .A(G57), .ZN(G237) );
  INV_X1 U612 ( .A(G132), .ZN(G219) );
  INV_X1 U613 ( .A(G82), .ZN(G220) );
  NAND2_X1 U614 ( .A1(G88), .A2(n645), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G75), .A2(n641), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n552) );
  NAND2_X1 U617 ( .A1(G62), .A2(n637), .ZN(n550) );
  NAND2_X1 U618 ( .A1(G50), .A2(n638), .ZN(n549) );
  NAND2_X1 U619 ( .A1(n550), .A2(n549), .ZN(n551) );
  NOR2_X1 U620 ( .A1(n552), .A2(n551), .ZN(G166) );
  NAND2_X1 U621 ( .A1(G64), .A2(n637), .ZN(n554) );
  NAND2_X1 U622 ( .A1(G52), .A2(n638), .ZN(n553) );
  NAND2_X1 U623 ( .A1(n554), .A2(n553), .ZN(n561) );
  XNOR2_X1 U624 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n641), .A2(G77), .ZN(n557) );
  NAND2_X1 U626 ( .A1(n645), .A2(G90), .ZN(n555) );
  XOR2_X1 U627 ( .A(KEYINPUT65), .B(n555), .Z(n556) );
  NAND2_X1 U628 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U629 ( .A(n559), .B(n558), .Z(n560) );
  NOR2_X1 U630 ( .A1(n561), .A2(n560), .ZN(G171) );
  NAND2_X1 U631 ( .A1(n645), .A2(G89), .ZN(n562) );
  XNOR2_X1 U632 ( .A(n562), .B(KEYINPUT4), .ZN(n564) );
  NAND2_X1 U633 ( .A1(G76), .A2(n641), .ZN(n563) );
  NAND2_X1 U634 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U636 ( .A1(G63), .A2(n637), .ZN(n567) );
  NAND2_X1 U637 ( .A1(G51), .A2(n638), .ZN(n566) );
  NAND2_X1 U638 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U640 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U641 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U644 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n835) );
  NAND2_X1 U646 ( .A1(n835), .A2(G567), .ZN(n573) );
  XOR2_X1 U647 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  NAND2_X1 U648 ( .A1(n645), .A2(G81), .ZN(n574) );
  XNOR2_X1 U649 ( .A(n574), .B(KEYINPUT12), .ZN(n576) );
  NAND2_X1 U650 ( .A1(G68), .A2(n641), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(n577), .ZN(n583) );
  NAND2_X1 U653 ( .A1(G56), .A2(n637), .ZN(n578) );
  XOR2_X1 U654 ( .A(KEYINPUT14), .B(n578), .Z(n581) );
  NAND2_X1 U655 ( .A1(G43), .A2(n638), .ZN(n579) );
  XNOR2_X1 U656 ( .A(KEYINPUT69), .B(n579), .ZN(n580) );
  NOR2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U658 ( .A1(n583), .A2(n582), .ZN(n989) );
  INV_X1 U659 ( .A(G860), .ZN(n604) );
  OR2_X1 U660 ( .A1(n989), .A2(n604), .ZN(G153) );
  INV_X1 U661 ( .A(G171), .ZN(G301) );
  NAND2_X1 U662 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U663 ( .A1(G66), .A2(n637), .ZN(n585) );
  NAND2_X1 U664 ( .A1(G54), .A2(n638), .ZN(n584) );
  NAND2_X1 U665 ( .A1(n585), .A2(n584), .ZN(n589) );
  NAND2_X1 U666 ( .A1(G92), .A2(n645), .ZN(n587) );
  NAND2_X1 U667 ( .A1(G79), .A2(n641), .ZN(n586) );
  NAND2_X1 U668 ( .A1(n587), .A2(n586), .ZN(n588) );
  NOR2_X1 U669 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U670 ( .A(KEYINPUT15), .B(n590), .Z(n910) );
  INV_X1 U671 ( .A(n910), .ZN(n973) );
  INV_X1 U672 ( .A(G868), .ZN(n601) );
  NAND2_X1 U673 ( .A1(n973), .A2(n601), .ZN(n591) );
  NAND2_X1 U674 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U675 ( .A1(G78), .A2(n641), .ZN(n599) );
  NAND2_X1 U676 ( .A1(G65), .A2(n637), .ZN(n594) );
  NAND2_X1 U677 ( .A1(G91), .A2(n645), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n597) );
  NAND2_X1 U679 ( .A1(G53), .A2(n638), .ZN(n595) );
  XNOR2_X1 U680 ( .A(KEYINPUT67), .B(n595), .ZN(n596) );
  NOR2_X1 U681 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U682 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U683 ( .A(n600), .B(KEYINPUT68), .ZN(G299) );
  NOR2_X1 U684 ( .A1(G286), .A2(n601), .ZN(n603) );
  NOR2_X1 U685 ( .A1(G299), .A2(G868), .ZN(n602) );
  NOR2_X1 U686 ( .A1(n603), .A2(n602), .ZN(G297) );
  NAND2_X1 U687 ( .A1(n604), .A2(G559), .ZN(n605) );
  NAND2_X1 U688 ( .A1(n605), .A2(n910), .ZN(n606) );
  XNOR2_X1 U689 ( .A(n606), .B(KEYINPUT16), .ZN(n607) );
  XNOR2_X1 U690 ( .A(KEYINPUT70), .B(n607), .ZN(G148) );
  NOR2_X1 U691 ( .A1(G868), .A2(n989), .ZN(n610) );
  NAND2_X1 U692 ( .A1(G868), .A2(n910), .ZN(n608) );
  NOR2_X1 U693 ( .A1(G559), .A2(n608), .ZN(n609) );
  NOR2_X1 U694 ( .A1(n610), .A2(n609), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G99), .A2(n893), .ZN(n611) );
  XNOR2_X1 U696 ( .A(n611), .B(KEYINPUT72), .ZN(n615) );
  XOR2_X1 U697 ( .A(KEYINPUT71), .B(KEYINPUT18), .Z(n613) );
  NAND2_X1 U698 ( .A1(G123), .A2(n897), .ZN(n612) );
  XNOR2_X1 U699 ( .A(n613), .B(n612), .ZN(n614) );
  NAND2_X1 U700 ( .A1(n615), .A2(n614), .ZN(n620) );
  NAND2_X1 U701 ( .A1(G111), .A2(n898), .ZN(n618) );
  BUF_X1 U702 ( .A(n616), .Z(n894) );
  NAND2_X1 U703 ( .A1(G135), .A2(n894), .ZN(n617) );
  NAND2_X1 U704 ( .A1(n618), .A2(n617), .ZN(n619) );
  NOR2_X1 U705 ( .A1(n620), .A2(n619), .ZN(n929) );
  XNOR2_X1 U706 ( .A(n929), .B(G2096), .ZN(n622) );
  INV_X1 U707 ( .A(G2100), .ZN(n621) );
  NAND2_X1 U708 ( .A1(n622), .A2(n621), .ZN(G156) );
  NAND2_X1 U709 ( .A1(G559), .A2(n910), .ZN(n623) );
  XNOR2_X1 U710 ( .A(n623), .B(n989), .ZN(n656) );
  NOR2_X1 U711 ( .A1(n656), .A2(G860), .ZN(n630) );
  NAND2_X1 U712 ( .A1(G67), .A2(n637), .ZN(n625) );
  NAND2_X1 U713 ( .A1(G55), .A2(n638), .ZN(n624) );
  NAND2_X1 U714 ( .A1(n625), .A2(n624), .ZN(n629) );
  NAND2_X1 U715 ( .A1(G93), .A2(n645), .ZN(n627) );
  NAND2_X1 U716 ( .A1(G80), .A2(n641), .ZN(n626) );
  NAND2_X1 U717 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U718 ( .A1(n629), .A2(n628), .ZN(n652) );
  XNOR2_X1 U719 ( .A(n630), .B(n652), .ZN(G145) );
  NAND2_X1 U720 ( .A1(G49), .A2(n638), .ZN(n632) );
  NAND2_X1 U721 ( .A1(G74), .A2(G651), .ZN(n631) );
  NAND2_X1 U722 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U723 ( .A1(n637), .A2(n633), .ZN(n636) );
  NAND2_X1 U724 ( .A1(n634), .A2(G87), .ZN(n635) );
  NAND2_X1 U725 ( .A1(n636), .A2(n635), .ZN(G288) );
  NAND2_X1 U726 ( .A1(G61), .A2(n637), .ZN(n640) );
  NAND2_X1 U727 ( .A1(G48), .A2(n638), .ZN(n639) );
  NAND2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U729 ( .A1(n641), .A2(G73), .ZN(n642) );
  XOR2_X1 U730 ( .A(KEYINPUT2), .B(n642), .Z(n643) );
  NOR2_X1 U731 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U732 ( .A1(n645), .A2(G86), .ZN(n646) );
  NAND2_X1 U733 ( .A1(n647), .A2(n646), .ZN(G305) );
  NOR2_X1 U734 ( .A1(n652), .A2(G868), .ZN(n648) );
  XNOR2_X1 U735 ( .A(KEYINPUT75), .B(n648), .ZN(n660) );
  XNOR2_X1 U736 ( .A(G166), .B(G288), .ZN(n655) );
  XNOR2_X1 U737 ( .A(KEYINPUT19), .B(KEYINPUT73), .ZN(n650) );
  XNOR2_X1 U738 ( .A(G290), .B(G299), .ZN(n649) );
  XNOR2_X1 U739 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U740 ( .A(n652), .B(n651), .ZN(n653) );
  XNOR2_X1 U741 ( .A(n653), .B(G305), .ZN(n654) );
  XNOR2_X1 U742 ( .A(n655), .B(n654), .ZN(n911) );
  XNOR2_X1 U743 ( .A(n911), .B(n656), .ZN(n657) );
  NAND2_X1 U744 ( .A1(n657), .A2(G868), .ZN(n658) );
  XNOR2_X1 U745 ( .A(KEYINPUT74), .B(n658), .ZN(n659) );
  NAND2_X1 U746 ( .A1(n660), .A2(n659), .ZN(G295) );
  NAND2_X1 U747 ( .A1(G2078), .A2(G2084), .ZN(n661) );
  XOR2_X1 U748 ( .A(KEYINPUT20), .B(n661), .Z(n662) );
  NAND2_X1 U749 ( .A1(G2090), .A2(n662), .ZN(n663) );
  XNOR2_X1 U750 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U751 ( .A1(n664), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U752 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U753 ( .A1(G220), .A2(G219), .ZN(n665) );
  XOR2_X1 U754 ( .A(KEYINPUT22), .B(n665), .Z(n666) );
  NOR2_X1 U755 ( .A1(G218), .A2(n666), .ZN(n667) );
  XNOR2_X1 U756 ( .A(KEYINPUT76), .B(n667), .ZN(n668) );
  NAND2_X1 U757 ( .A1(n668), .A2(G96), .ZN(n839) );
  NAND2_X1 U758 ( .A1(n839), .A2(G2106), .ZN(n672) );
  NAND2_X1 U759 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U760 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U761 ( .A1(G108), .A2(n670), .ZN(n840) );
  NAND2_X1 U762 ( .A1(n840), .A2(G567), .ZN(n671) );
  NAND2_X1 U763 ( .A1(n672), .A2(n671), .ZN(n841) );
  NAND2_X1 U764 ( .A1(G483), .A2(G661), .ZN(n673) );
  NOR2_X1 U765 ( .A1(n841), .A2(n673), .ZN(n674) );
  XOR2_X1 U766 ( .A(KEYINPUT77), .B(n674), .Z(n838) );
  NAND2_X1 U767 ( .A1(n838), .A2(G36), .ZN(G176) );
  INV_X1 U768 ( .A(G166), .ZN(G303) );
  NAND2_X1 U769 ( .A1(G40), .A2(G160), .ZN(n675) );
  XNOR2_X2 U770 ( .A(n675), .B(KEYINPUT79), .ZN(n776) );
  NAND2_X2 U771 ( .A1(n778), .A2(n776), .ZN(n727) );
  NAND2_X1 U772 ( .A1(G2072), .A2(n704), .ZN(n677) );
  XNOR2_X1 U773 ( .A(n677), .B(n676), .ZN(n679) );
  INV_X1 U774 ( .A(G1956), .ZN(n976) );
  NOR2_X1 U775 ( .A1(n976), .A2(n704), .ZN(n678) );
  INV_X1 U776 ( .A(G299), .ZN(n699) );
  NAND2_X1 U777 ( .A1(n700), .A2(n699), .ZN(n698) );
  XNOR2_X1 U778 ( .A(n681), .B(n680), .ZN(n683) );
  NAND2_X1 U779 ( .A1(n704), .A2(G2067), .ZN(n682) );
  NAND2_X1 U780 ( .A1(n683), .A2(n682), .ZN(n685) );
  NAND2_X1 U781 ( .A1(n693), .A2(n910), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n727), .A2(G1341), .ZN(n686) );
  XNOR2_X1 U783 ( .A(n686), .B(KEYINPUT90), .ZN(n690) );
  XNOR2_X1 U784 ( .A(G1996), .B(KEYINPUT89), .ZN(n959) );
  NOR2_X1 U785 ( .A1(n959), .A2(n727), .ZN(n687) );
  XNOR2_X1 U786 ( .A(KEYINPUT26), .B(n687), .ZN(n688) );
  NOR2_X1 U787 ( .A1(n989), .A2(n688), .ZN(n689) );
  NAND2_X1 U788 ( .A1(n690), .A2(n689), .ZN(n691) );
  NAND2_X1 U789 ( .A1(n692), .A2(n691), .ZN(n696) );
  INV_X1 U790 ( .A(n693), .ZN(n694) );
  NAND2_X1 U791 ( .A1(n973), .A2(n694), .ZN(n695) );
  NAND2_X1 U792 ( .A1(n696), .A2(n695), .ZN(n697) );
  NAND2_X1 U793 ( .A1(n698), .A2(n697), .ZN(n702) );
  NAND2_X1 U794 ( .A1(n702), .A2(n519), .ZN(n703) );
  XNOR2_X1 U795 ( .A(n703), .B(KEYINPUT29), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n727), .A2(G1961), .ZN(n706) );
  XOR2_X1 U797 ( .A(G2078), .B(KEYINPUT25), .Z(n954) );
  NAND2_X1 U798 ( .A1(n704), .A2(n954), .ZN(n705) );
  NAND2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  XOR2_X1 U800 ( .A(n707), .B(KEYINPUT86), .Z(n718) );
  AND2_X1 U801 ( .A1(n718), .A2(G171), .ZN(n708) );
  XOR2_X1 U802 ( .A(KEYINPUT87), .B(n708), .Z(n709) );
  NOR2_X1 U803 ( .A1(G1966), .A2(n726), .ZN(n712) );
  INV_X1 U804 ( .A(KEYINPUT85), .ZN(n711) );
  XNOR2_X1 U805 ( .A(n712), .B(n711), .ZN(n738) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n727), .ZN(n741) );
  NOR2_X1 U807 ( .A1(n738), .A2(n741), .ZN(n713) );
  NAND2_X1 U808 ( .A1(G8), .A2(n713), .ZN(n716) );
  INV_X1 U809 ( .A(KEYINPUT30), .ZN(n714) );
  NOR2_X1 U810 ( .A1(G168), .A2(n717), .ZN(n720) );
  NOR2_X1 U811 ( .A1(G171), .A2(n718), .ZN(n719) );
  NOR2_X1 U812 ( .A1(n720), .A2(n719), .ZN(n721) );
  XNOR2_X1 U813 ( .A(n721), .B(KEYINPUT31), .ZN(n722) );
  NOR2_X2 U814 ( .A1(n723), .A2(n722), .ZN(n739) );
  INV_X1 U815 ( .A(n739), .ZN(n725) );
  AND2_X1 U816 ( .A1(G286), .A2(G8), .ZN(n724) );
  NAND2_X1 U817 ( .A1(n725), .A2(n724), .ZN(n734) );
  INV_X1 U818 ( .A(G8), .ZN(n732) );
  NOR2_X1 U819 ( .A1(G1971), .A2(n726), .ZN(n729) );
  NOR2_X1 U820 ( .A1(G2090), .A2(n727), .ZN(n728) );
  NOR2_X1 U821 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U822 ( .A1(n730), .A2(G303), .ZN(n731) );
  OR2_X1 U823 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U824 ( .A1(n734), .A2(n733), .ZN(n735) );
  INV_X1 U825 ( .A(KEYINPUT32), .ZN(n736) );
  XNOR2_X1 U826 ( .A(n737), .B(n736), .ZN(n763) );
  NOR2_X1 U827 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U828 ( .A(n740), .B(KEYINPUT94), .ZN(n744) );
  NAND2_X1 U829 ( .A1(G8), .A2(n741), .ZN(n742) );
  XNOR2_X1 U830 ( .A(KEYINPUT84), .B(n742), .ZN(n743) );
  AND2_X1 U831 ( .A1(n744), .A2(n743), .ZN(n762) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n978) );
  INV_X1 U833 ( .A(n978), .ZN(n748) );
  NOR2_X1 U834 ( .A1(G1976), .A2(G288), .ZN(n746) );
  XOR2_X1 U835 ( .A(KEYINPUT97), .B(n746), .Z(n756) );
  NOR2_X1 U836 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U837 ( .A1(n756), .A2(n747), .ZN(n979) );
  NOR2_X1 U838 ( .A1(n748), .A2(n979), .ZN(n749) );
  NOR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U840 ( .A(n751), .B(KEYINPUT98), .ZN(n752) );
  NOR2_X1 U841 ( .A1(n752), .A2(n726), .ZN(n753) );
  INV_X1 U842 ( .A(n753), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n755), .A2(n754), .ZN(n761) );
  INV_X1 U844 ( .A(n756), .ZN(n757) );
  NOR2_X1 U845 ( .A1(n726), .A2(n757), .ZN(n758) );
  NAND2_X1 U846 ( .A1(KEYINPUT33), .A2(n758), .ZN(n760) );
  XNOR2_X1 U847 ( .A(G1981), .B(G305), .ZN(n986) );
  NAND2_X1 U848 ( .A1(n761), .A2(n517), .ZN(n770) );
  NOR2_X1 U849 ( .A1(n762), .A2(n763), .ZN(n766) );
  NAND2_X1 U850 ( .A1(G8), .A2(G166), .ZN(n764) );
  NOR2_X1 U851 ( .A1(G2090), .A2(n764), .ZN(n765) );
  NOR2_X1 U852 ( .A1(n766), .A2(n765), .ZN(n767) );
  XNOR2_X1 U853 ( .A(n767), .B(KEYINPUT99), .ZN(n768) );
  NAND2_X1 U854 ( .A1(n768), .A2(n726), .ZN(n769) );
  NAND2_X1 U855 ( .A1(n770), .A2(n769), .ZN(n771) );
  XNOR2_X1 U856 ( .A(n771), .B(KEYINPUT100), .ZN(n775) );
  NOR2_X1 U857 ( .A1(G1981), .A2(G305), .ZN(n772) );
  XOR2_X1 U858 ( .A(n772), .B(KEYINPUT24), .Z(n773) );
  NOR2_X1 U859 ( .A1(n726), .A2(n773), .ZN(n774) );
  NOR2_X1 U860 ( .A1(n775), .A2(n774), .ZN(n808) );
  INV_X1 U861 ( .A(n776), .ZN(n777) );
  NOR2_X1 U862 ( .A1(n778), .A2(n777), .ZN(n821) );
  XNOR2_X1 U863 ( .A(KEYINPUT37), .B(G2067), .ZN(n811) );
  NAND2_X1 U864 ( .A1(G140), .A2(n894), .ZN(n779) );
  XNOR2_X1 U865 ( .A(n779), .B(KEYINPUT80), .ZN(n781) );
  NAND2_X1 U866 ( .A1(G104), .A2(n893), .ZN(n780) );
  NAND2_X1 U867 ( .A1(n781), .A2(n780), .ZN(n783) );
  XOR2_X1 U868 ( .A(KEYINPUT81), .B(KEYINPUT34), .Z(n782) );
  XNOR2_X1 U869 ( .A(n783), .B(n782), .ZN(n788) );
  NAND2_X1 U870 ( .A1(G128), .A2(n897), .ZN(n785) );
  NAND2_X1 U871 ( .A1(G116), .A2(n898), .ZN(n784) );
  NAND2_X1 U872 ( .A1(n785), .A2(n784), .ZN(n786) );
  XOR2_X1 U873 ( .A(KEYINPUT35), .B(n786), .Z(n787) );
  NOR2_X1 U874 ( .A1(n788), .A2(n787), .ZN(n789) );
  XNOR2_X1 U875 ( .A(KEYINPUT36), .B(n789), .ZN(n907) );
  NOR2_X1 U876 ( .A1(n811), .A2(n907), .ZN(n942) );
  NAND2_X1 U877 ( .A1(n821), .A2(n942), .ZN(n818) );
  NAND2_X1 U878 ( .A1(G129), .A2(n897), .ZN(n791) );
  NAND2_X1 U879 ( .A1(G117), .A2(n898), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n791), .A2(n790), .ZN(n795) );
  NAND2_X1 U881 ( .A1(G105), .A2(n893), .ZN(n792) );
  XNOR2_X1 U882 ( .A(n792), .B(KEYINPUT38), .ZN(n793) );
  XNOR2_X1 U883 ( .A(n793), .B(KEYINPUT83), .ZN(n794) );
  NOR2_X1 U884 ( .A1(n795), .A2(n794), .ZN(n797) );
  NAND2_X1 U885 ( .A1(G141), .A2(n894), .ZN(n796) );
  NAND2_X1 U886 ( .A1(n797), .A2(n796), .ZN(n880) );
  NAND2_X1 U887 ( .A1(G1996), .A2(n880), .ZN(n806) );
  NAND2_X1 U888 ( .A1(G95), .A2(n893), .ZN(n799) );
  NAND2_X1 U889 ( .A1(G119), .A2(n897), .ZN(n798) );
  NAND2_X1 U890 ( .A1(n799), .A2(n798), .ZN(n802) );
  NAND2_X1 U891 ( .A1(n898), .A2(G107), .ZN(n800) );
  XOR2_X1 U892 ( .A(KEYINPUT82), .B(n800), .Z(n801) );
  NOR2_X1 U893 ( .A1(n802), .A2(n801), .ZN(n804) );
  NAND2_X1 U894 ( .A1(G131), .A2(n894), .ZN(n803) );
  NAND2_X1 U895 ( .A1(n804), .A2(n803), .ZN(n876) );
  NAND2_X1 U896 ( .A1(G1991), .A2(n876), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n806), .A2(n805), .ZN(n930) );
  NAND2_X1 U898 ( .A1(n821), .A2(n930), .ZN(n814) );
  NAND2_X1 U899 ( .A1(n818), .A2(n814), .ZN(n807) );
  NOR2_X1 U900 ( .A1(n808), .A2(n807), .ZN(n810) );
  XNOR2_X1 U901 ( .A(G1986), .B(G290), .ZN(n975) );
  NAND2_X1 U902 ( .A1(n975), .A2(n821), .ZN(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n824) );
  NAND2_X1 U904 ( .A1(n811), .A2(n907), .ZN(n939) );
  NOR2_X1 U905 ( .A1(G1991), .A2(n876), .ZN(n931) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U907 ( .A1(n931), .A2(n812), .ZN(n813) );
  XNOR2_X1 U908 ( .A(n813), .B(KEYINPUT101), .ZN(n815) );
  NAND2_X1 U909 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U910 ( .A1(n880), .A2(G1996), .ZN(n934) );
  NAND2_X1 U911 ( .A1(n816), .A2(n934), .ZN(n817) );
  XOR2_X1 U912 ( .A(KEYINPUT39), .B(n817), .Z(n819) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n820) );
  NAND2_X1 U914 ( .A1(n939), .A2(n820), .ZN(n822) );
  NAND2_X1 U915 ( .A1(n822), .A2(n821), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n824), .A2(n823), .ZN(n825) );
  XNOR2_X1 U917 ( .A(n825), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U918 ( .A(G1348), .B(G2454), .ZN(n826) );
  XNOR2_X1 U919 ( .A(n826), .B(G2430), .ZN(n827) );
  XNOR2_X1 U920 ( .A(n827), .B(G1341), .ZN(n833) );
  XOR2_X1 U921 ( .A(G2443), .B(G2427), .Z(n829) );
  XNOR2_X1 U922 ( .A(G2438), .B(G2446), .ZN(n828) );
  XNOR2_X1 U923 ( .A(n829), .B(n828), .ZN(n831) );
  XOR2_X1 U924 ( .A(G2451), .B(G2435), .Z(n830) );
  XNOR2_X1 U925 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U926 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U927 ( .A1(n834), .A2(G14), .ZN(n918) );
  XOR2_X1 U928 ( .A(KEYINPUT102), .B(n918), .Z(G401) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U931 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U932 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U933 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U935 ( .A(G120), .ZN(G236) );
  INV_X1 U936 ( .A(G96), .ZN(G221) );
  INV_X1 U937 ( .A(G69), .ZN(G235) );
  NOR2_X1 U938 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U939 ( .A(G325), .ZN(G261) );
  INV_X1 U940 ( .A(n841), .ZN(G319) );
  XOR2_X1 U941 ( .A(G1966), .B(G1981), .Z(n843) );
  XNOR2_X1 U942 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U943 ( .A(n843), .B(n842), .ZN(n853) );
  XOR2_X1 U944 ( .A(KEYINPUT105), .B(KEYINPUT41), .Z(n845) );
  XNOR2_X1 U945 ( .A(G1956), .B(KEYINPUT106), .ZN(n844) );
  XNOR2_X1 U946 ( .A(n845), .B(n844), .ZN(n849) );
  XOR2_X1 U947 ( .A(G1976), .B(G1961), .Z(n847) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1971), .ZN(n846) );
  XNOR2_X1 U949 ( .A(n847), .B(n846), .ZN(n848) );
  XOR2_X1 U950 ( .A(n849), .B(n848), .Z(n851) );
  XNOR2_X1 U951 ( .A(KEYINPUT104), .B(G2474), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(G229) );
  XOR2_X1 U954 ( .A(KEYINPUT103), .B(G2072), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2090), .B(G2078), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n856), .B(G2100), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2084), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U960 ( .A(G2096), .B(KEYINPUT43), .Z(n860) );
  XNOR2_X1 U961 ( .A(G2678), .B(KEYINPUT42), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(n862), .B(n861), .Z(G227) );
  NAND2_X1 U964 ( .A1(G100), .A2(n893), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G112), .A2(n898), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n871) );
  NAND2_X1 U967 ( .A1(G136), .A2(n894), .ZN(n865) );
  XNOR2_X1 U968 ( .A(KEYINPUT107), .B(n865), .ZN(n868) );
  NAND2_X1 U969 ( .A1(n897), .A2(G124), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT44), .B(n866), .Z(n867) );
  NOR2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  XOR2_X1 U972 ( .A(KEYINPUT108), .B(n869), .Z(n870) );
  NOR2_X1 U973 ( .A1(n871), .A2(n870), .ZN(n872) );
  XOR2_X1 U974 ( .A(KEYINPUT109), .B(n872), .Z(G162) );
  XOR2_X1 U975 ( .A(KEYINPUT46), .B(KEYINPUT112), .Z(n874) );
  XNOR2_X1 U976 ( .A(KEYINPUT113), .B(KEYINPUT48), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U978 ( .A(KEYINPUT114), .B(n875), .ZN(n878) );
  XNOR2_X1 U979 ( .A(n876), .B(n929), .ZN(n877) );
  XNOR2_X1 U980 ( .A(n878), .B(n877), .ZN(n879) );
  XOR2_X1 U981 ( .A(n880), .B(n879), .Z(n882) );
  XNOR2_X1 U982 ( .A(G164), .B(G160), .ZN(n881) );
  XNOR2_X1 U983 ( .A(n882), .B(n881), .ZN(n892) );
  NAND2_X1 U984 ( .A1(G106), .A2(n893), .ZN(n884) );
  NAND2_X1 U985 ( .A1(G142), .A2(n894), .ZN(n883) );
  NAND2_X1 U986 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U987 ( .A(n885), .B(KEYINPUT45), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G130), .A2(n897), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n890) );
  NAND2_X1 U990 ( .A1(n898), .A2(G118), .ZN(n888) );
  XOR2_X1 U991 ( .A(KEYINPUT110), .B(n888), .Z(n889) );
  NOR2_X1 U992 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U993 ( .A(n892), .B(n891), .Z(n906) );
  NAND2_X1 U994 ( .A1(G103), .A2(n893), .ZN(n896) );
  NAND2_X1 U995 ( .A1(G139), .A2(n894), .ZN(n895) );
  NAND2_X1 U996 ( .A1(n896), .A2(n895), .ZN(n903) );
  NAND2_X1 U997 ( .A1(G127), .A2(n897), .ZN(n900) );
  NAND2_X1 U998 ( .A1(G115), .A2(n898), .ZN(n899) );
  NAND2_X1 U999 ( .A1(n900), .A2(n899), .ZN(n901) );
  XOR2_X1 U1000 ( .A(KEYINPUT47), .B(n901), .Z(n902) );
  NOR2_X1 U1001 ( .A1(n903), .A2(n902), .ZN(n904) );
  XOR2_X1 U1002 ( .A(KEYINPUT111), .B(n904), .Z(n923) );
  XNOR2_X1 U1003 ( .A(G162), .B(n923), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n908) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1006 ( .A1(G37), .A2(n909), .ZN(G395) );
  XOR2_X1 U1007 ( .A(n911), .B(n910), .Z(n913) );
  XNOR2_X1 U1008 ( .A(G286), .B(G171), .ZN(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(n914) );
  XNOR2_X1 U1010 ( .A(n914), .B(n989), .ZN(n915) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n915), .ZN(G397) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n916) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n916), .Z(n917) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n921) );
  NOR2_X1 U1015 ( .A1(G395), .A2(G397), .ZN(n919) );
  XNOR2_X1 U1016 ( .A(KEYINPUT115), .B(n919), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(n921), .A2(n920), .ZN(n922) );
  NAND2_X1 U1018 ( .A1(G319), .A2(n922), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(G2072), .B(n923), .ZN(n924) );
  XNOR2_X1 U1022 ( .A(n924), .B(KEYINPUT117), .ZN(n926) );
  XOR2_X1 U1023 ( .A(G2078), .B(G164), .Z(n925) );
  NOR2_X1 U1024 ( .A1(n926), .A2(n925), .ZN(n927) );
  XOR2_X1 U1025 ( .A(KEYINPUT50), .B(n927), .Z(n945) );
  XOR2_X1 U1026 ( .A(G2084), .B(G160), .Z(n928) );
  NOR2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n933) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n933), .A2(n932), .ZN(n938) );
  XNOR2_X1 U1030 ( .A(G162), .B(G2090), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  XOR2_X1 U1032 ( .A(KEYINPUT51), .B(n936), .Z(n937) );
  NOR2_X1 U1033 ( .A1(n938), .A2(n937), .ZN(n940) );
  NAND2_X1 U1034 ( .A1(n940), .A2(n939), .ZN(n941) );
  NOR2_X1 U1035 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1036 ( .A(KEYINPUT116), .B(n943), .Z(n944) );
  NOR2_X1 U1037 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1038 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  XOR2_X1 U1039 ( .A(KEYINPUT55), .B(KEYINPUT118), .Z(n949) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n949), .ZN(n948) );
  NAND2_X1 U1041 ( .A1(n948), .A2(G29), .ZN(n1030) );
  XOR2_X1 U1042 ( .A(n949), .B(KEYINPUT120), .Z(n969) );
  XNOR2_X1 U1043 ( .A(G2090), .B(G35), .ZN(n964) );
  XNOR2_X1 U1044 ( .A(KEYINPUT119), .B(G2067), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(n950), .B(G26), .ZN(n958) );
  XNOR2_X1 U1046 ( .A(G1991), .B(G25), .ZN(n952) );
  XNOR2_X1 U1047 ( .A(G33), .B(G2072), .ZN(n951) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(G28), .A2(n953), .ZN(n956) );
  XNOR2_X1 U1050 ( .A(G27), .B(n954), .ZN(n955) );
  NOR2_X1 U1051 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1052 ( .A1(n958), .A2(n957), .ZN(n961) );
  XOR2_X1 U1053 ( .A(G32), .B(n959), .Z(n960) );
  NOR2_X1 U1054 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1055 ( .A(KEYINPUT53), .B(n962), .ZN(n963) );
  NOR2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1057 ( .A(G2084), .B(G34), .Z(n965) );
  XNOR2_X1 U1058 ( .A(KEYINPUT54), .B(n965), .ZN(n966) );
  NAND2_X1 U1059 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1060 ( .A(n969), .B(n968), .ZN(n970) );
  NOR2_X1 U1061 ( .A1(G29), .A2(n970), .ZN(n971) );
  XNOR2_X1 U1062 ( .A(n971), .B(KEYINPUT121), .ZN(n972) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n972), .ZN(n1028) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n999) );
  XNOR2_X1 U1065 ( .A(G1348), .B(n973), .ZN(n974) );
  NOR2_X1 U1066 ( .A1(n975), .A2(n974), .ZN(n997) );
  NAND2_X1 U1067 ( .A1(G303), .A2(G1971), .ZN(n983) );
  XNOR2_X1 U1068 ( .A(G299), .B(KEYINPUT123), .ZN(n977) );
  XNOR2_X1 U1069 ( .A(n977), .B(n976), .ZN(n981) );
  NAND2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1071 ( .A1(n981), .A2(n980), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1073 ( .A(n984), .B(KEYINPUT124), .ZN(n995) );
  XOR2_X1 U1074 ( .A(G1966), .B(G168), .Z(n985) );
  NOR2_X1 U1075 ( .A1(n986), .A2(n985), .ZN(n987) );
  XOR2_X1 U1076 ( .A(KEYINPUT57), .B(n987), .Z(n988) );
  XNOR2_X1 U1077 ( .A(KEYINPUT122), .B(n988), .ZN(n993) );
  XNOR2_X1 U1078 ( .A(G301), .B(G1961), .ZN(n991) );
  XNOR2_X1 U1079 ( .A(n989), .B(G1341), .ZN(n990) );
  NOR2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NOR2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1084 ( .A1(n999), .A2(n998), .ZN(n1026) );
  INV_X1 U1085 ( .A(G16), .ZN(n1024) );
  XNOR2_X1 U1086 ( .A(G1961), .B(G5), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G21), .ZN(n1000) );
  NOR2_X1 U1088 ( .A1(n1001), .A2(n1000), .ZN(n1013) );
  XOR2_X1 U1089 ( .A(KEYINPUT126), .B(G4), .Z(n1003) );
  XNOR2_X1 U1090 ( .A(G1348), .B(KEYINPUT59), .ZN(n1002) );
  XNOR2_X1 U1091 ( .A(n1003), .B(n1002), .ZN(n1006) );
  XOR2_X1 U1092 ( .A(KEYINPUT125), .B(G1956), .Z(n1004) );
  XNOR2_X1 U1093 ( .A(G20), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1094 ( .A1(n1006), .A2(n1005), .ZN(n1010) );
  XNOR2_X1 U1095 ( .A(G1981), .B(G6), .ZN(n1008) );
  XNOR2_X1 U1096 ( .A(G1341), .B(G19), .ZN(n1007) );
  NOR2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NAND2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1099 ( .A(KEYINPUT60), .B(n1011), .Z(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1020) );
  XNOR2_X1 U1101 ( .A(G1971), .B(G22), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G23), .B(G1976), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1017) );
  XOR2_X1 U1104 ( .A(G1986), .B(G24), .Z(n1016) );
  NAND2_X1 U1105 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1106 ( .A(KEYINPUT58), .B(n1018), .ZN(n1019) );
  NOR2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XOR2_X1 U1108 ( .A(n1021), .B(KEYINPUT61), .Z(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT127), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1112 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1113 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1114 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1115 ( .A(G311), .ZN(G150) );
endmodule

