//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 1 0 0 1 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n239, new_n240, new_n241, new_n243, new_n244, new_n245,
    new_n246, new_n247, new_n248, new_n249, new_n250, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n257, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293;
  XNOR2_X1  g0000(.A(KEYINPUT64), .B(G50), .ZN(new_n201));
  NOR2_X1   g0001(.A1(G58), .A2(G68), .ZN(new_n202));
  INV_X1    g0002(.A(new_n202), .ZN(new_n203));
  NOR3_X1   g0003(.A1(new_n201), .A2(G77), .A3(new_n203), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XOR2_X1   g0008(.A(new_n208), .B(KEYINPUT0), .Z(new_n209));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G257), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G107), .A2(G264), .ZN(new_n213));
  INV_X1    g0013(.A(G50), .ZN(new_n214));
  INV_X1    g0014(.A(G226), .ZN(new_n215));
  INV_X1    g0015(.A(G116), .ZN(new_n216));
  INV_X1    g0016(.A(G270), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  AOI211_X1 g0018(.A(new_n212), .B(new_n218), .C1(G77), .C2(G244), .ZN(new_n219));
  INV_X1    g0019(.A(G58), .ZN(new_n220));
  INV_X1    g0020(.A(G232), .ZN(new_n221));
  INV_X1    g0021(.A(G238), .ZN(new_n222));
  AND2_X1   g0022(.A1(KEYINPUT68), .A2(G68), .ZN(new_n223));
  NOR2_X1   g0023(.A1(KEYINPUT68), .A2(G68), .ZN(new_n224));
  NOR2_X1   g0024(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g0025(.A(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n222), .C2(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(G87), .ZN(new_n228));
  INV_X1    g0028(.A(G250), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  OAI21_X1  g0030(.A(new_n206), .B1(new_n227), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(KEYINPUT1), .ZN(new_n232));
  NAND3_X1  g0032(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n233));
  INV_X1    g0033(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(KEYINPUT65), .B1(G1), .B2(G13), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g0036(.A(G20), .ZN(new_n237));
  NOR2_X1   g0037(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT66), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n203), .A2(G50), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n240), .B(KEYINPUT67), .Z(new_n241));
  AOI211_X1 g0041(.A(new_n209), .B(new_n232), .C1(new_n239), .C2(new_n241), .ZN(G361));
  XNOR2_X1  g0042(.A(G238), .B(G244), .ZN(new_n243));
  XNOR2_X1  g0043(.A(G226), .B(G232), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(G250), .B(G257), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(G264), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n249), .B(new_n217), .ZN(new_n250));
  XOR2_X1   g0050(.A(new_n247), .B(new_n250), .Z(G358));
  XNOR2_X1  g0051(.A(G68), .B(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(new_n214), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n253), .B(G58), .ZN(new_n254));
  XOR2_X1   g0054(.A(G107), .B(G116), .Z(new_n255));
  XNOR2_X1  g0055(.A(G87), .B(G97), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XNOR2_X1  g0057(.A(new_n254), .B(new_n257), .ZN(G351));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(KEYINPUT71), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT71), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G33), .A3(G41), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G1), .A2(G13), .ZN(new_n263));
  INV_X1    g0063(.A(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G1), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(G41), .B2(G45), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT70), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n266), .B(KEYINPUT70), .C1(G41), .C2(G45), .ZN(new_n270));
  NAND4_X1  g0070(.A1(new_n265), .A2(G274), .A3(new_n269), .A4(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n259), .B1(new_n234), .B2(new_n235), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G97), .ZN(new_n274));
  INV_X1    g0074(.A(G1698), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n215), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n221), .A2(G1698), .ZN(new_n277));
  AND2_X1   g0077(.A1(KEYINPUT3), .A2(G33), .ZN(new_n278));
  NOR2_X1   g0078(.A1(KEYINPUT3), .A2(G33), .ZN(new_n279));
  OAI211_X1 g0079(.A(new_n276), .B(new_n277), .C1(new_n278), .C2(new_n279), .ZN(new_n280));
  AOI21_X1  g0080(.A(new_n273), .B1(new_n274), .B2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n272), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT72), .ZN(new_n283));
  AND3_X1   g0083(.A1(new_n265), .A2(new_n283), .A3(new_n267), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n283), .B1(new_n265), .B2(new_n267), .ZN(new_n285));
  OAI21_X1  g0085(.A(G238), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n282), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n287), .B1(new_n282), .B2(new_n286), .ZN(new_n290));
  OAI21_X1  g0090(.A(G200), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n266), .A2(G13), .A3(G20), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(KEYINPUT12), .ZN(new_n294));
  INV_X1    g0094(.A(KEYINPUT65), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n263), .A2(new_n295), .ZN(new_n296));
  NAND3_X1  g0096(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n233), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(G1), .B2(new_n237), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT12), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n294), .B1(new_n301), .B2(G68), .ZN(new_n302));
  INV_X1    g0102(.A(G13), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n303), .A2(G1), .ZN(new_n304));
  NAND4_X1  g0104(.A1(new_n226), .A2(KEYINPUT12), .A3(G20), .A4(new_n304), .ZN(new_n305));
  NOR2_X1   g0105(.A1(G20), .A2(G33), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(G50), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n237), .A2(G33), .ZN(new_n309));
  OAI221_X1 g0109(.A(new_n307), .B1(new_n308), .B2(new_n309), .C1(new_n225), .C2(new_n237), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(new_n298), .ZN(new_n311));
  AND2_X1   g0111(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(KEYINPUT11), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n302), .B(new_n305), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n265), .A2(new_n267), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(KEYINPUT72), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n265), .A2(new_n283), .A3(new_n267), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n222), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n280), .A2(new_n274), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n271), .B1(new_n320), .B2(new_n273), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT13), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n322), .A2(new_n288), .A3(G190), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n291), .A2(new_n315), .A3(new_n323), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n322), .A2(new_n288), .A3(G179), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT78), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(KEYINPUT77), .B2(KEYINPUT14), .ZN(new_n328));
  OAI211_X1 g0128(.A(G169), .B(new_n328), .C1(new_n289), .C2(new_n290), .ZN(new_n329));
  INV_X1    g0129(.A(G169), .ZN(new_n330));
  AND2_X1   g0130(.A1(new_n327), .A2(KEYINPUT14), .ZN(new_n331));
  AOI211_X1 g0131(.A(new_n330), .B(new_n331), .C1(new_n322), .C2(new_n288), .ZN(new_n332));
  OAI211_X1 g0132(.A(new_n326), .B(new_n329), .C1(new_n332), .C2(new_n328), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n325), .B1(new_n333), .B2(new_n314), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n317), .A2(new_n318), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n272), .B1(new_n335), .B2(G226), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT73), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n278), .A2(new_n279), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(G223), .B2(G1698), .ZN(new_n339));
  INV_X1    g0139(.A(G222), .ZN(new_n340));
  OAI21_X1  g0140(.A(new_n339), .B1(new_n340), .B2(G1698), .ZN(new_n341));
  AOI22_X1  g0141(.A1(new_n296), .A2(new_n233), .B1(G33), .B2(G41), .ZN(new_n342));
  INV_X1    g0142(.A(KEYINPUT3), .ZN(new_n343));
  INV_X1    g0143(.A(G33), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(KEYINPUT3), .A2(G33), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n341), .B(new_n342), .C1(G77), .C2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n336), .A2(new_n337), .A3(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n337), .B1(new_n336), .B2(new_n348), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n350), .A2(new_n351), .A3(G169), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n336), .A2(new_n348), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(KEYINPUT73), .ZN(new_n354));
  AOI21_X1  g0154(.A(G179), .B1(new_n354), .B2(new_n349), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n306), .A2(G150), .ZN(new_n356));
  OAI21_X1  g0156(.A(G20), .B1(new_n201), .B2(new_n203), .ZN(new_n357));
  XNOR2_X1  g0157(.A(KEYINPUT8), .B(G58), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n358), .A2(KEYINPUT74), .ZN(new_n359));
  OR3_X1    g0159(.A1(new_n220), .A2(KEYINPUT74), .A3(KEYINPUT8), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n356), .B(new_n357), .C1(new_n361), .C2(new_n309), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n298), .ZN(new_n363));
  INV_X1    g0163(.A(new_n300), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(G50), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n293), .A2(new_n214), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n352), .A2(new_n355), .A3(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(G190), .B1(new_n350), .B2(new_n351), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n354), .A2(G200), .A3(new_n349), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n367), .A2(KEYINPUT9), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT9), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n363), .A2(new_n373), .A3(new_n365), .A4(new_n366), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT10), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT10), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n370), .A2(new_n371), .A3(new_n378), .A4(new_n375), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n369), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT75), .ZN(new_n381));
  INV_X1    g0181(.A(G244), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n317), .B2(new_n318), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n381), .B1(new_n383), .B2(new_n272), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n284), .A2(new_n285), .ZN(new_n385));
  OAI211_X1 g0185(.A(KEYINPUT75), .B(new_n271), .C1(new_n385), .C2(new_n382), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n338), .B1(G238), .B2(G1698), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n387), .B1(new_n221), .B2(G1698), .ZN(new_n388));
  OAI211_X1 g0188(.A(new_n388), .B(new_n342), .C1(G107), .C2(new_n347), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n384), .A2(new_n386), .A3(new_n389), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G20), .A2(G77), .ZN(new_n392));
  INV_X1    g0192(.A(new_n306), .ZN(new_n393));
  XNOR2_X1  g0193(.A(KEYINPUT15), .B(G87), .ZN(new_n394));
  OAI221_X1 g0194(.A(new_n392), .B1(new_n358), .B2(new_n393), .C1(new_n394), .C2(new_n309), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n364), .A2(G77), .B1(new_n298), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(G77), .B2(new_n292), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT76), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n397), .B1(new_n390), .B2(G200), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT76), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(G190), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n398), .B(new_n401), .C1(new_n402), .C2(new_n390), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n390), .A2(G179), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n390), .A2(new_n330), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n397), .A3(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(KEYINPUT18), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n361), .A2(new_n293), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n300), .B2(new_n361), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n393), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n202), .B1(new_n225), .B2(G58), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n237), .ZN(new_n414));
  INV_X1    g0214(.A(G68), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n345), .A2(new_n237), .A3(new_n346), .ZN(new_n416));
  INV_X1    g0216(.A(KEYINPUT7), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n345), .A2(KEYINPUT7), .A3(new_n237), .A4(new_n346), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n415), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n414), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n299), .B1(new_n421), .B2(KEYINPUT16), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT16), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n226), .B1(new_n418), .B2(new_n419), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n423), .B1(new_n414), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n409), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n215), .A2(G1698), .ZN(new_n427));
  OAI221_X1 g0227(.A(new_n427), .B1(G223), .B2(G1698), .C1(new_n278), .C2(new_n279), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n342), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n265), .A2(G232), .A3(new_n267), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n431), .A2(G179), .A3(new_n271), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n271), .A2(new_n432), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n273), .B1(new_n428), .B2(new_n429), .ZN(new_n435));
  OAI21_X1  g0235(.A(G169), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n433), .A2(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n407), .B1(new_n426), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(KEYINPUT7), .B1(new_n338), .B2(new_n237), .ZN(new_n440));
  INV_X1    g0240(.A(new_n419), .ZN(new_n441));
  OAI21_X1  g0241(.A(G68), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OR2_X1    g0242(.A1(KEYINPUT68), .A2(G68), .ZN(new_n443));
  NAND2_X1  g0243(.A1(KEYINPUT68), .A2(G68), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(G58), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n203), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n411), .B1(new_n446), .B2(G20), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n442), .A2(new_n447), .A3(KEYINPUT16), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n425), .A2(new_n298), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n409), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n451), .A2(KEYINPUT18), .A3(new_n437), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n439), .A2(new_n452), .ZN(new_n453));
  NAND4_X1  g0253(.A1(new_n431), .A2(G190), .A3(new_n271), .A4(new_n432), .ZN(new_n454));
  OAI21_X1  g0254(.A(G200), .B1(new_n434), .B2(new_n435), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n449), .A2(new_n450), .A3(new_n454), .A4(new_n455), .ZN(new_n456));
  XNOR2_X1  g0256(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT17), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(KEYINPUT79), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n459), .B1(new_n461), .B2(new_n456), .ZN(new_n462));
  AND3_X1   g0262(.A1(new_n406), .A2(new_n453), .A3(new_n462), .ZN(new_n463));
  AND4_X1   g0263(.A1(new_n334), .A2(new_n380), .A3(new_n403), .A4(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT4), .ZN(new_n465));
  NOR2_X1   g0265(.A1(new_n465), .A2(G1698), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n466), .B(G244), .C1(new_n279), .C2(new_n278), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G283), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n382), .B1(new_n345), .B2(new_n346), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n467), .B(new_n468), .C1(new_n469), .C2(KEYINPUT4), .ZN(new_n470));
  OAI21_X1  g0270(.A(G250), .B1(new_n278), .B2(new_n279), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n275), .B1(new_n471), .B2(KEYINPUT4), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n342), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G45), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n474), .A2(G1), .ZN(new_n475));
  XNOR2_X1  g0275(.A(KEYINPUT5), .B(G41), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n265), .A2(G274), .A3(new_n475), .A4(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(KEYINPUT5), .A2(G41), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n475), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n265), .A2(new_n481), .A3(G257), .ZN(new_n482));
  AND2_X1   g0282(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n473), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n330), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT81), .ZN(new_n486));
  AND3_X1   g0286(.A1(new_n477), .A2(new_n482), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n486), .B1(new_n477), .B2(new_n482), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n473), .A2(KEYINPUT80), .ZN(new_n490));
  INV_X1    g0290(.A(G179), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT80), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n492), .B(new_n342), .C1(new_n470), .C2(new_n472), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n489), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT82), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n292), .A2(G97), .ZN(new_n496));
  OAI21_X1  g0296(.A(G107), .B1(new_n440), .B2(new_n441), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT6), .ZN(new_n498));
  AND2_X1   g0298(.A1(G97), .A2(G107), .ZN(new_n499));
  NOR2_X1   g0299(.A1(G97), .A2(G107), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(G107), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n502), .A2(KEYINPUT6), .A3(G97), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n504), .A2(G20), .B1(G77), .B2(new_n306), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n496), .B1(new_n506), .B2(new_n298), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n266), .A2(G33), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n292), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n298), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G97), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n495), .B1(new_n507), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n299), .B1(new_n497), .B2(new_n505), .ZN(new_n513));
  INV_X1    g0313(.A(new_n511), .ZN(new_n514));
  NOR4_X1   g0314(.A1(new_n513), .A2(KEYINPUT82), .A3(new_n514), .A4(new_n496), .ZN(new_n515));
  OAI211_X1 g0315(.A(new_n485), .B(new_n494), .C1(new_n512), .C2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n489), .A2(new_n490), .A3(new_n493), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G200), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n506), .A2(new_n298), .ZN(new_n519));
  INV_X1    g0319(.A(new_n496), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(new_n511), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n521), .ZN(new_n522));
  INV_X1    g0322(.A(new_n484), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G190), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n518), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n222), .A2(new_n275), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n382), .A2(G1698), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n526), .B(new_n527), .C1(new_n278), .C2(new_n279), .ZN(new_n528));
  NAND2_X1  g0328(.A1(G33), .A2(G116), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n342), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  AND3_X1   g0332(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n229), .B1(new_n474), .B2(G1), .ZN(new_n534));
  INV_X1    g0334(.A(G274), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n266), .A2(new_n535), .A3(G45), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n532), .B1(new_n533), .B2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n265), .A2(KEYINPUT83), .A3(new_n534), .A4(new_n536), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n531), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n540), .A2(new_n330), .ZN(new_n541));
  XNOR2_X1  g0341(.A(new_n394), .B(KEYINPUT84), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n510), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n500), .A2(new_n228), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n274), .A2(new_n237), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n544), .A2(KEYINPUT19), .A3(new_n545), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n237), .B(G68), .C1(new_n278), .C2(new_n279), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n274), .A2(G20), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n546), .B(new_n547), .C1(KEYINPUT19), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n298), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n394), .A2(new_n293), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n543), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  OAI211_X1 g0352(.A(new_n541), .B(new_n552), .C1(G179), .C2(new_n540), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n510), .A2(G87), .ZN(new_n554));
  AND3_X1   g0354(.A1(new_n550), .A2(new_n551), .A3(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n540), .A2(G200), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n531), .A2(new_n538), .A3(G190), .A4(new_n539), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n553), .A2(new_n558), .ZN(new_n559));
  AND3_X1   g0359(.A1(new_n516), .A2(new_n525), .A3(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT21), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n292), .A2(G116), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n298), .A2(new_n509), .A3(new_n216), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n468), .B(new_n237), .C1(G33), .C2(new_n210), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n216), .A2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n298), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT20), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND4_X1  g0368(.A1(new_n298), .A2(KEYINPUT20), .A3(new_n564), .A4(new_n565), .ZN(new_n569));
  AOI211_X1 g0369(.A(new_n562), .B(new_n563), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(G303), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n345), .A2(new_n571), .A3(new_n346), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n275), .A2(G257), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G264), .A2(G1698), .ZN(new_n574));
  OAI211_X1 g0374(.A(new_n573), .B(new_n574), .C1(new_n278), .C2(new_n279), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n342), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n265), .A2(new_n481), .A3(G270), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n576), .A2(new_n477), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(G169), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n561), .B1(new_n570), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n568), .A2(new_n569), .ZN(new_n581));
  INV_X1    g0381(.A(new_n562), .ZN(new_n582));
  INV_X1    g0382(.A(new_n563), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n584), .A2(KEYINPUT21), .A3(G169), .A4(new_n578), .ZN(new_n585));
  AND3_X1   g0385(.A1(new_n576), .A2(new_n477), .A3(new_n577), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(G179), .A3(new_n586), .ZN(new_n587));
  AND3_X1   g0387(.A1(new_n580), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT87), .ZN(new_n589));
  OAI21_X1  g0389(.A(new_n589), .B1(new_n237), .B2(G107), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT23), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n237), .A2(G33), .A3(G116), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n502), .A2(G20), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n589), .A3(KEYINPUT23), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n592), .A2(new_n593), .A3(new_n595), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n237), .B(G87), .C1(new_n278), .C2(new_n279), .ZN(new_n597));
  XNOR2_X1  g0397(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n597), .A2(new_n598), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n596), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT24), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI211_X1 g0403(.A(new_n596), .B(KEYINPUT24), .C1(new_n599), .C2(new_n600), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n603), .A2(new_n298), .A3(new_n604), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n292), .A2(new_n508), .ZN(new_n606));
  NAND4_X1  g0406(.A1(new_n606), .A2(new_n236), .A3(G107), .A4(new_n297), .ZN(new_n607));
  INV_X1    g0407(.A(new_n304), .ZN(new_n608));
  OR3_X1    g0408(.A1(new_n608), .A2(KEYINPUT25), .A3(new_n594), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT25), .B1(new_n608), .B2(new_n594), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n607), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT88), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g0413(.A1(new_n607), .A2(new_n609), .A3(KEYINPUT88), .A4(new_n610), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n605), .A2(new_n615), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n265), .A2(new_n481), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n229), .A2(new_n275), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n211), .A2(G1698), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n618), .B(new_n619), .C1(new_n278), .C2(new_n279), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G33), .A2(G294), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  AOI22_X1  g0422(.A1(new_n617), .A2(G264), .B1(new_n622), .B2(new_n342), .ZN(new_n623));
  AOI21_X1  g0423(.A(G169), .B1(new_n623), .B2(new_n477), .ZN(new_n624));
  INV_X1    g0424(.A(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n622), .A2(new_n342), .ZN(new_n626));
  NAND3_X1  g0426(.A1(new_n265), .A2(new_n481), .A3(G264), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n626), .A2(new_n477), .A3(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n628), .A2(G179), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n616), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  INV_X1    g0431(.A(G200), .ZN(new_n632));
  OAI211_X1 g0432(.A(new_n570), .B(KEYINPUT85), .C1(new_n632), .C2(new_n586), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT85), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n586), .A2(new_n632), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n634), .B1(new_n635), .B2(new_n584), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n586), .A2(G190), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n633), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n628), .A2(new_n632), .ZN(new_n639));
  OAI211_X1 g0439(.A(new_n639), .B(KEYINPUT89), .C1(G190), .C2(new_n628), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT89), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n628), .A2(new_n641), .A3(new_n632), .ZN(new_n642));
  NAND4_X1  g0442(.A1(new_n640), .A2(new_n615), .A3(new_n605), .A4(new_n642), .ZN(new_n643));
  AND4_X1   g0443(.A1(new_n588), .A2(new_n631), .A3(new_n638), .A4(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n464), .A2(new_n560), .A3(new_n644), .ZN(G372));
  NAND2_X1  g0445(.A1(new_n553), .A2(new_n558), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n521), .B1(new_n517), .B2(G200), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n646), .B1(new_n647), .B2(new_n524), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n588), .A2(new_n631), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n648), .A2(new_n649), .A3(new_n516), .A4(new_n643), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n494), .A2(new_n553), .A3(new_n558), .A4(new_n485), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n651), .A2(KEYINPUT26), .A3(new_n522), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n512), .A2(new_n515), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT26), .B1(new_n651), .B2(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n553), .B(KEYINPUT90), .ZN(new_n656));
  INV_X1    g0456(.A(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n650), .A2(new_n653), .A3(new_n655), .A4(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n464), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n377), .A2(new_n379), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n333), .A2(new_n314), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n324), .A2(new_n404), .A3(new_n397), .A4(new_n405), .ZN(new_n662));
  INV_X1    g0462(.A(new_n461), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n426), .A2(new_n663), .A3(new_n454), .A4(new_n455), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n661), .A2(new_n662), .B1(new_n459), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n453), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n660), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n369), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n667), .A2(KEYINPUT91), .A3(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g0470(.A(KEYINPUT91), .B1(new_n667), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g0471(.A(new_n659), .B1(new_n670), .B2(new_n671), .ZN(G369));
  NAND2_X1  g0472(.A1(new_n588), .A2(new_n638), .ZN(new_n673));
  OR3_X1    g0473(.A1(new_n608), .A2(KEYINPUT27), .A3(G20), .ZN(new_n674));
  OAI21_X1  g0474(.A(KEYINPUT27), .B1(new_n608), .B2(G20), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(G213), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n584), .A2(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n580), .A2(new_n585), .A3(new_n587), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(new_n679), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT92), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n684), .A2(new_n685), .A3(G330), .ZN(new_n686));
  INV_X1    g0486(.A(G330), .ZN(new_n687));
  OAI21_X1  g0487(.A(KEYINPUT92), .B1(new_n683), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI211_X1 g0489(.A(new_n629), .B(new_n624), .C1(new_n605), .C2(new_n615), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n616), .A2(new_n678), .ZN(new_n691));
  AOI21_X1  g0491(.A(new_n690), .B1(new_n643), .B2(new_n691), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n631), .A2(new_n678), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n678), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n681), .A2(new_n696), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT93), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n693), .B1(new_n698), .B2(new_n694), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n695), .A2(new_n699), .ZN(G399));
  INV_X1    g0500(.A(new_n207), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n701), .A2(G41), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G1), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n500), .A2(new_n228), .A3(new_n216), .ZN(new_n705));
  OAI22_X1  g0505(.A1(new_n704), .A2(new_n705), .B1(new_n240), .B2(new_n703), .ZN(new_n706));
  XNOR2_X1  g0506(.A(new_n706), .B(KEYINPUT28), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT29), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n516), .A2(new_n525), .A3(new_n559), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n643), .B1(new_n690), .B2(new_n681), .ZN(new_n710));
  OAI211_X1 g0510(.A(new_n655), .B(new_n657), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  OAI211_X1 g0511(.A(new_n708), .B(new_n696), .C1(new_n711), .C2(new_n652), .ZN(new_n712));
  INV_X1    g0512(.A(new_n710), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n656), .B1(new_n560), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n654), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT26), .ZN(new_n716));
  AND2_X1   g0516(.A1(new_n494), .A2(new_n485), .ZN(new_n717));
  NAND4_X1  g0517(.A1(new_n715), .A2(new_n716), .A3(new_n717), .A4(new_n559), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT26), .B1(new_n651), .B2(new_n522), .ZN(new_n719));
  AND2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n678), .B1(new_n714), .B2(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n712), .B1(new_n721), .B2(new_n708), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n560), .A2(new_n644), .A3(new_n696), .ZN(new_n724));
  NOR3_X1   g0524(.A1(new_n540), .A2(new_n491), .A3(new_n578), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n523), .A2(new_n725), .A3(new_n623), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT30), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n523), .A2(new_n725), .A3(KEYINPUT30), .A4(new_n623), .ZN(new_n729));
  NAND4_X1  g0529(.A1(new_n517), .A2(new_n491), .A3(new_n540), .A4(new_n628), .ZN(new_n730));
  OAI211_X1 g0530(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n586), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(new_n678), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT31), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n678), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n724), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G330), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n723), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n707), .B1(new_n739), .B2(G1), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT94), .ZN(G364));
  INV_X1    g0541(.A(new_n689), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n303), .A2(G20), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n704), .B1(G45), .B2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n742), .B(new_n745), .C1(G330), .C2(new_n684), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n236), .B1(G20), .B2(new_n330), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n237), .A2(new_n402), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n632), .A2(G179), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n338), .B1(new_n751), .B2(new_n571), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT99), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n402), .A2(G20), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n491), .A2(new_n632), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G317), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(KEYINPUT33), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n758), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G322), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n491), .A2(G200), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n749), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n762), .B1(new_n763), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g0566(.A(new_n766), .B(KEYINPUT100), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G179), .A2(G200), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n755), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI211_X1 g0570(.A(new_n753), .B(new_n767), .C1(G329), .C2(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n749), .A2(new_n756), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT97), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  XNOR2_X1  g0574(.A(KEYINPUT98), .B(G326), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n754), .A2(G179), .A3(new_n632), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G283), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n755), .A2(new_n764), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n237), .B1(new_n768), .B2(G190), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(new_n780), .A2(G311), .B1(G294), .B2(new_n782), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n771), .A2(new_n776), .A3(new_n778), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n782), .A2(G97), .ZN(new_n785));
  OAI221_X1 g0585(.A(new_n785), .B1(new_n220), .B2(new_n765), .C1(new_n415), .C2(new_n757), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT32), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n787), .B1(new_n769), .B2(new_n410), .ZN(new_n788));
  NAND3_X1  g0588(.A1(new_n770), .A2(KEYINPUT32), .A3(G159), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n786), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n751), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n791), .A2(G87), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n780), .A2(G77), .ZN(new_n793));
  INV_X1    g0593(.A(new_n777), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n794), .A2(new_n502), .B1(new_n214), .B2(new_n772), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n338), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n790), .A2(new_n792), .A3(new_n793), .A4(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n748), .B1(new_n784), .B2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(G13), .A2(G33), .ZN(new_n799));
  XNOR2_X1  g0599(.A(new_n799), .B(KEYINPUT96), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n800), .A2(G20), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n745), .B(new_n798), .C1(new_n683), .C2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n241), .A2(new_n474), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n338), .A2(new_n207), .ZN(new_n804));
  XNOR2_X1  g0604(.A(new_n804), .B(KEYINPUT95), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n803), .B(new_n805), .C1(new_n254), .C2(new_n474), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n701), .A2(new_n338), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n807), .A2(G355), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n806), .B(new_n808), .C1(G116), .C2(new_n207), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n801), .A2(new_n747), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n802), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g0612(.A1(new_n746), .A2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  NOR2_X1   g0614(.A1(new_n399), .A2(new_n400), .ZN(new_n815));
  AOI211_X1 g0615(.A(KEYINPUT76), .B(new_n397), .C1(new_n390), .C2(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n390), .A2(new_n402), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n397), .A2(new_n678), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n406), .B1(new_n818), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n406), .A2(new_n678), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n800), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n747), .A2(new_n825), .ZN(new_n827));
  XOR2_X1   g0627(.A(new_n827), .B(KEYINPUT101), .Z(new_n828));
  INV_X1    g0628(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n308), .ZN(new_n830));
  OAI221_X1 g0630(.A(new_n785), .B1(new_n502), .B2(new_n751), .C1(new_n571), .C2(new_n772), .ZN(new_n831));
  INV_X1    g0631(.A(G311), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n794), .A2(new_n228), .B1(new_n769), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n338), .B1(new_n779), .B2(new_n216), .ZN(new_n834));
  NOR3_X1   g0634(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(G283), .ZN(new_n836));
  INV_X1    g0636(.A(G294), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n835), .B1(new_n836), .B2(new_n757), .C1(new_n837), .C2(new_n765), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n794), .A2(new_n415), .B1(new_n214), .B2(new_n751), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n338), .B(new_n839), .C1(G58), .C2(new_n782), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n769), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT102), .ZN(new_n843));
  INV_X1    g0643(.A(new_n765), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n780), .A2(G159), .B1(new_n844), .B2(G143), .ZN(new_n845));
  INV_X1    g0645(.A(G137), .ZN(new_n846));
  INV_X1    g0646(.A(G150), .ZN(new_n847));
  OAI221_X1 g0647(.A(new_n845), .B1(new_n846), .B2(new_n772), .C1(new_n847), .C2(new_n757), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT34), .Z(new_n849));
  OAI21_X1  g0649(.A(new_n838), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(new_n747), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n826), .A2(new_n744), .A3(new_n830), .A4(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n696), .B1(new_n711), .B2(new_n652), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n824), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n818), .A2(new_n820), .ZN(new_n855));
  NAND4_X1  g0655(.A1(new_n658), .A2(new_n855), .A3(new_n406), .A4(new_n696), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g0657(.A(new_n857), .B(new_n737), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n852), .B1(new_n858), .B2(new_n744), .ZN(G384));
  XNOR2_X1  g0659(.A(KEYINPUT107), .B(KEYINPUT40), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT38), .ZN(new_n861));
  OAI21_X1  g0661(.A(new_n423), .B1(new_n414), .B2(new_n420), .ZN(new_n862));
  NAND3_X1  g0662(.A1(new_n862), .A2(new_n298), .A3(new_n448), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(new_n450), .ZN(new_n864));
  INV_X1    g0664(.A(new_n676), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(new_n453), .B2(new_n462), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n425), .A2(new_n298), .A3(new_n448), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n868), .A2(new_n409), .B1(new_n437), .B2(new_n865), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n869), .A2(new_n870), .A3(new_n456), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n433), .A2(new_n436), .A3(new_n676), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n864), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n870), .B1(new_n873), .B2(new_n456), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n861), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT105), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n873), .A2(new_n456), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(KEYINPUT37), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n869), .A2(new_n870), .A3(new_n456), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g0681(.A1(new_n439), .A2(new_n452), .B1(new_n664), .B2(new_n459), .ZN(new_n882));
  OAI211_X1 g0682(.A(KEYINPUT38), .B(new_n881), .C1(new_n882), .C2(new_n866), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(new_n877), .A3(new_n883), .ZN(new_n884));
  OAI211_X1 g0684(.A(KEYINPUT105), .B(new_n861), .C1(new_n867), .C2(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n314), .A2(new_n678), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n661), .A2(new_n324), .A3(new_n887), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n314), .B(new_n678), .C1(new_n325), .C2(new_n333), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND4_X1  g0690(.A1(new_n736), .A2(new_n890), .A3(new_n823), .A4(new_n821), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n860), .B1(new_n886), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT40), .ZN(new_n893));
  AOI22_X1  g0693(.A1(new_n438), .A2(new_n676), .B1(new_n449), .B2(new_n450), .ZN(new_n894));
  OAI21_X1  g0694(.A(KEYINPUT37), .B1(new_n894), .B2(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n869), .A2(new_n456), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g0697(.A1(new_n869), .A2(KEYINPUT106), .A3(KEYINPUT37), .A4(new_n456), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n451), .A2(new_n865), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n453), .B2(new_n462), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n861), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n893), .B1(new_n902), .B2(new_n883), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n403), .A2(new_n819), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n822), .B1(new_n904), .B2(new_n406), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n903), .A2(new_n736), .A3(new_n905), .A4(new_n890), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n892), .A2(G330), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n464), .A2(G330), .A3(new_n736), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT108), .Z(new_n910));
  NAND2_X1  g0710(.A1(new_n464), .A2(new_n736), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n892), .A2(new_n906), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n406), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n914), .B1(new_n403), .B2(new_n819), .ZN(new_n915));
  OAI21_X1  g0715(.A(new_n823), .B1(new_n853), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n916), .A2(new_n890), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(KEYINPUT104), .ZN(new_n918));
  INV_X1    g0718(.A(new_n886), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n916), .A2(new_n920), .A3(new_n890), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n918), .A2(new_n919), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n884), .A2(KEYINPUT39), .A3(new_n885), .ZN(new_n923));
  INV_X1    g0723(.A(KEYINPUT39), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n902), .A2(new_n924), .A3(new_n883), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n661), .A2(new_n678), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n666), .A2(new_n676), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n922), .A2(new_n928), .A3(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n671), .ZN(new_n931));
  AOI22_X1  g0731(.A1(new_n931), .A2(new_n669), .B1(new_n722), .B2(new_n464), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n930), .B(new_n932), .ZN(new_n933));
  XNOR2_X1  g0733(.A(new_n913), .B(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n934), .B1(new_n266), .B2(new_n743), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n504), .B(KEYINPUT103), .Z(new_n936));
  AOI21_X1  g0736(.A(new_n216), .B1(new_n936), .B2(KEYINPUT35), .ZN(new_n937));
  OAI211_X1 g0737(.A(new_n937), .B(new_n239), .C1(KEYINPUT35), .C2(new_n936), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT36), .ZN(new_n939));
  NAND4_X1  g0739(.A1(new_n445), .A2(G50), .A3(G77), .A4(new_n203), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n415), .B2(new_n201), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n941), .A2(G1), .A3(new_n303), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n935), .A2(new_n939), .A3(new_n942), .ZN(G367));
  NAND2_X1  g0743(.A1(new_n698), .A2(new_n694), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n516), .B(new_n525), .C1(new_n522), .C2(new_n696), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n717), .A2(new_n521), .A3(new_n678), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  OR3_X1    g0748(.A1(new_n944), .A2(new_n948), .A3(KEYINPUT42), .ZN(new_n949));
  OAI21_X1  g0749(.A(KEYINPUT42), .B1(new_n944), .B2(new_n948), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n947), .A2(new_n690), .B1(new_n717), .B2(new_n715), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n949), .B(new_n950), .C1(new_n951), .C2(new_n678), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n696), .A2(new_n555), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n656), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n646), .B2(new_n953), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n689), .A2(new_n694), .A3(new_n947), .ZN(new_n958));
  INV_X1    g0758(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n952), .A2(new_n958), .A3(new_n956), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT109), .ZN(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n962), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n702), .B(KEYINPUT41), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(KEYINPUT110), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n699), .B2(new_n947), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n699), .A2(new_n969), .A3(new_n947), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n971), .A2(KEYINPUT45), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT45), .ZN(new_n974));
  INV_X1    g0774(.A(new_n972), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n970), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  INV_X1    g0777(.A(new_n699), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n977), .B1(new_n978), .B2(new_n948), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n699), .A2(KEYINPUT44), .A3(new_n947), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n976), .A3(new_n981), .ZN(new_n982));
  INV_X1    g0782(.A(new_n695), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND4_X1  g0784(.A1(new_n973), .A2(new_n976), .A3(new_n981), .A4(new_n695), .ZN(new_n985));
  INV_X1    g0785(.A(new_n694), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(new_n698), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n742), .A2(new_n987), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n742), .A2(new_n987), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND4_X1  g0790(.A1(new_n984), .A2(new_n739), .A3(new_n985), .A4(new_n990), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n968), .B1(new_n991), .B2(new_n739), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n266), .B1(new_n743), .B2(G45), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n966), .B1(new_n992), .B2(new_n994), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n773), .A2(new_n832), .B1(new_n571), .B2(new_n765), .ZN(new_n996));
  XOR2_X1   g0796(.A(new_n996), .B(KEYINPUT111), .Z(new_n997));
  OAI22_X1  g0797(.A1(new_n794), .A2(new_n210), .B1(new_n781), .B2(new_n502), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n347), .B(new_n998), .C1(G317), .C2(new_n770), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n997), .B(new_n999), .C1(new_n836), .C2(new_n779), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(G294), .B2(new_n758), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n791), .A2(G116), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT46), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n774), .A2(G143), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n757), .A2(new_n410), .B1(new_n781), .B2(new_n415), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n769), .A2(new_n846), .B1(new_n751), .B2(new_n220), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1006), .B(KEYINPUT112), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n844), .A2(G150), .B1(new_n777), .B2(G77), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1007), .A2(new_n347), .A3(new_n1008), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1005), .B(new_n1009), .C1(new_n201), .C2(new_n780), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1001), .A2(new_n1003), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT47), .Z(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n747), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n801), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n955), .A2(new_n1014), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n805), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n810), .B1(new_n207), .B2(new_n394), .C1(new_n250), .C2(new_n1016), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1013), .A2(new_n744), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  AND3_X1   g0818(.A1(new_n995), .A2(KEYINPUT113), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(KEYINPUT113), .B1(new_n995), .B2(new_n1018), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1020), .A2(new_n1022), .ZN(G387));
  NAND2_X1  g0823(.A1(new_n990), .A2(new_n739), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n738), .A2(new_n988), .A3(new_n989), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1024), .A2(new_n702), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1016), .B1(new_n247), .B2(G45), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n1027), .B1(new_n705), .B2(new_n807), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n358), .A2(G50), .ZN(new_n1029));
  XOR2_X1   g0829(.A(new_n1029), .B(KEYINPUT50), .Z(new_n1030));
  NOR2_X1   g0830(.A1(new_n415), .A2(new_n308), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1030), .A2(G45), .A3(new_n1031), .A4(new_n705), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1028), .A2(new_n1032), .B1(G107), .B2(new_n207), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n745), .B1(new_n1033), .B2(new_n810), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1034), .B1(new_n694), .B2(new_n1014), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n765), .A2(new_n214), .ZN(new_n1036));
  INV_X1    g0836(.A(new_n542), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(new_n781), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n1036), .B(new_n1038), .C1(G150), .C2(new_n770), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n791), .A2(G77), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n410), .B2(new_n772), .C1(new_n361), .C2(new_n757), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n338), .B(new_n1041), .C1(G68), .C2(new_n780), .ZN(new_n1042));
  OAI211_X1 g0842(.A(new_n1039), .B(new_n1042), .C1(new_n210), .C2(new_n794), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(new_n758), .A2(G311), .B1(new_n844), .B2(G317), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n571), .B2(new_n779), .C1(new_n773), .C2(new_n763), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT48), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n1046), .B1(new_n836), .B2(new_n781), .C1(new_n837), .C2(new_n751), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OR2_X1    g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n770), .A2(new_n775), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n777), .A2(G116), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n1049), .A2(new_n338), .A3(new_n1050), .A4(new_n1051), .ZN(new_n1052));
  AND2_X1   g0852(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1043), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1035), .B1(new_n1054), .B2(new_n747), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1055), .B1(new_n990), .B2(new_n994), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1026), .A2(new_n1056), .ZN(G393));
  NAND2_X1  g0857(.A1(new_n984), .A2(new_n985), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1058), .A2(new_n1024), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1059), .A2(new_n702), .A3(new_n991), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n984), .A2(new_n994), .A3(new_n985), .ZN(new_n1061));
  OAI221_X1 g0861(.A(new_n810), .B1(new_n210), .B2(new_n207), .C1(new_n1016), .C2(new_n257), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n769), .A2(new_n763), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n772), .A2(new_n759), .B1(new_n765), .B2(new_n832), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT114), .B(KEYINPUT52), .Z(new_n1065));
  XNOR2_X1  g0865(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n794), .A2(new_n502), .B1(new_n836), .B2(new_n751), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1067), .B1(G294), .B2(new_n780), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n782), .A2(G116), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n347), .B1(new_n758), .B2(G303), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .A4(new_n1070), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n772), .A2(new_n847), .B1(new_n765), .B2(new_n410), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT51), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n770), .A2(G143), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n338), .B1(new_n777), .B2(G87), .ZN(new_n1075));
  OAI22_X1  g0875(.A1(new_n226), .A2(new_n751), .B1(new_n779), .B2(new_n358), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n201), .B2(new_n758), .ZN(new_n1077));
  NAND4_X1  g0877(.A1(new_n1073), .A2(new_n1074), .A3(new_n1075), .A4(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n781), .A2(new_n308), .ZN(new_n1079));
  OAI22_X1  g0879(.A1(new_n1063), .A2(new_n1071), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n745), .B1(new_n1080), .B2(new_n747), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1062), .B(new_n1081), .C1(new_n947), .C2(new_n1014), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1060), .A2(new_n1061), .A3(new_n1082), .ZN(G390));
  INV_X1    g0883(.A(new_n890), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1084), .B1(new_n737), .B2(new_n824), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n905), .A2(G330), .A3(new_n736), .A4(new_n890), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n822), .B1(new_n721), .B2(new_n821), .ZN(new_n1087));
  AND3_X1   g0887(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1085), .A2(new_n1086), .B1(new_n823), .B2(new_n856), .ZN(new_n1089));
  OAI211_X1 g0889(.A(new_n932), .B(new_n908), .C1(new_n1088), .C2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n927), .B1(new_n902), .B2(new_n883), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n1087), .B2(new_n1084), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n927), .B1(new_n916), .B2(new_n890), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1092), .B(new_n1086), .C1(new_n1093), .C2(new_n926), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1084), .B1(new_n856), .B2(new_n823), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n923), .B(new_n925), .C1(new_n1096), .C2(new_n927), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1086), .B1(new_n1097), .B2(new_n1092), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1090), .B1(new_n1095), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n712), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n650), .A2(new_n657), .A3(new_n719), .A4(new_n718), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n708), .B1(new_n1101), .B2(new_n696), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n464), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1103), .B(new_n908), .C1(new_n670), .C2(new_n671), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1085), .A2(new_n1086), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n916), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1085), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1104), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1092), .B1(new_n1093), .B2(new_n926), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n1086), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1108), .A2(new_n1111), .A3(new_n1094), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1099), .A2(new_n1112), .A3(new_n702), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT115), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1099), .A2(new_n1112), .A3(KEYINPUT115), .A4(new_n702), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1115), .A2(new_n1116), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n926), .A2(new_n800), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n791), .A2(G150), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT53), .ZN(new_n1120));
  OAI22_X1  g0920(.A1(new_n765), .A2(new_n841), .B1(new_n781), .B2(new_n410), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n777), .A2(new_n201), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1123), .B1(new_n846), .B2(new_n757), .ZN(new_n1124));
  XOR2_X1   g0924(.A(KEYINPUT54), .B(G143), .Z(new_n1125));
  AOI211_X1 g0925(.A(new_n338), .B(new_n1124), .C1(new_n780), .C2(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g0927(.A(G125), .ZN(new_n1128));
  INV_X1    g0928(.A(G128), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1127), .B1(new_n1128), .B2(new_n769), .C1(new_n1129), .C2(new_n772), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n792), .A2(new_n338), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT116), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n1079), .B1(G68), .B2(new_n777), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n757), .A2(new_n502), .B1(new_n779), .B2(new_n210), .ZN(new_n1134));
  INV_X1    g0934(.A(new_n772), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1134), .B1(G283), .B2(new_n1135), .ZN(new_n1136));
  AND3_X1   g0936(.A1(new_n1132), .A2(new_n1133), .A3(new_n1136), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n216), .B2(new_n765), .C1(new_n837), .C2(new_n769), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n748), .B1(new_n1130), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n828), .B1(new_n360), .B2(new_n359), .ZN(new_n1140));
  NOR4_X1   g0940(.A1(new_n1118), .A2(new_n745), .A3(new_n1139), .A4(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1095), .A2(new_n1098), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n1142), .B2(new_n994), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1117), .A2(new_n1143), .ZN(G378));
  AOI211_X1 g0944(.A(G41), .B(new_n347), .C1(new_n777), .C2(G58), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1145), .B(new_n1040), .C1(new_n836), .C2(new_n769), .ZN(new_n1146));
  XOR2_X1   g0946(.A(new_n1146), .B(KEYINPUT117), .Z(new_n1147));
  NOR2_X1   g0947(.A1(new_n772), .A2(new_n216), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n757), .A2(new_n210), .B1(new_n781), .B2(new_n415), .ZN(new_n1149));
  NOR3_X1   g0949(.A1(new_n1147), .A2(new_n1148), .A3(new_n1149), .ZN(new_n1150));
  OAI221_X1 g0950(.A(new_n1150), .B1(new_n502), .B2(new_n765), .C1(new_n1037), .C2(new_n779), .ZN(new_n1151));
  XNOR2_X1  g0951(.A(new_n1151), .B(KEYINPUT58), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n214), .B1(new_n278), .B2(G41), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n781), .A2(new_n847), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n779), .A2(new_n846), .B1(new_n765), .B2(new_n1129), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1154), .B(new_n1155), .C1(new_n791), .C2(new_n1125), .ZN(new_n1156));
  OAI221_X1 g0956(.A(new_n1156), .B1(new_n1128), .B2(new_n772), .C1(new_n841), .C2(new_n757), .ZN(new_n1157));
  XOR2_X1   g0957(.A(new_n1157), .B(KEYINPUT59), .Z(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n770), .C2(G124), .ZN(new_n1159));
  OAI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(new_n410), .C2(new_n794), .ZN(new_n1160));
  AND3_X1   g0960(.A1(new_n1152), .A2(new_n1153), .A3(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n744), .B1(new_n201), .B2(new_n828), .C1(new_n1161), .C2(new_n748), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n660), .A2(new_n668), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  XNOR2_X1  g0964(.A(new_n1164), .B(KEYINPUT118), .ZN(new_n1165));
  AND2_X1   g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(new_n368), .B2(new_n676), .ZN(new_n1168));
  OR2_X1    g0968(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n368), .A2(new_n676), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1162), .B1(new_n825), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT119), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1174), .B(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n922), .A2(new_n928), .A3(new_n929), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1168), .A2(new_n1172), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n907), .A2(new_n1179), .ZN(new_n1180));
  NAND4_X1  g0980(.A1(new_n1173), .A2(new_n892), .A3(G330), .A4(new_n906), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n930), .A2(new_n1181), .A3(new_n1180), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1104), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1112), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1177), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1176), .B1(new_n1188), .B2(new_n702), .ZN(new_n1189));
  AND2_X1   g0989(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1190));
  OAI21_X1  g0990(.A(KEYINPUT121), .B1(new_n1190), .B2(new_n930), .ZN(new_n1191));
  INV_X1    g0991(.A(KEYINPUT121), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1178), .A2(new_n1182), .A3(new_n1192), .ZN(new_n1193));
  OAI21_X1  g0993(.A(KEYINPUT120), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT120), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n930), .A2(new_n1195), .A3(new_n1181), .A4(new_n1180), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1191), .A2(new_n1193), .A3(new_n1194), .A4(new_n1196), .ZN(new_n1197));
  AOI211_X1 g0997(.A(KEYINPUT57), .B(new_n703), .C1(new_n1112), .C2(new_n1186), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1197), .B1(new_n994), .B2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1189), .A2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(KEYINPUT122), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g1002(.A1(new_n1189), .A2(new_n1199), .A3(KEYINPUT122), .ZN(new_n1203));
  AND2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(G375));
  NOR2_X1   g1005(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1206), .A2(new_n993), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n794), .A2(new_n308), .B1(new_n502), .B2(new_n779), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n338), .B1(new_n769), .B2(new_n571), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n751), .A2(new_n210), .ZN(new_n1210));
  OR3_X1    g1010(.A1(new_n1038), .A2(new_n1209), .A3(new_n1210), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1208), .B(new_n1211), .C1(G283), .C2(new_n844), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n1212), .B1(new_n216), .B2(new_n757), .C1(new_n837), .C2(new_n772), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1135), .A2(G132), .B1(G58), .B2(new_n777), .ZN(new_n1214));
  OAI221_X1 g1014(.A(new_n1214), .B1(new_n847), .B2(new_n779), .C1(new_n410), .C2(new_n751), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1215), .B1(G50), .B2(new_n782), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n844), .A2(G137), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n758), .A2(new_n1125), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n338), .B1(new_n770), .B2(G128), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1216), .A2(new_n1217), .A3(new_n1218), .A4(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n748), .B1(new_n1213), .B2(new_n1220), .ZN(new_n1221));
  AOI211_X1 g1021(.A(new_n745), .B(new_n1221), .C1(new_n415), .C2(new_n829), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT124), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n890), .A2(new_n800), .ZN(new_n1224));
  XNOR2_X1  g1024(.A(new_n1224), .B(KEYINPUT123), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1207), .B1(new_n1223), .B2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1206), .A2(new_n1104), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1227), .A2(new_n967), .A3(new_n1090), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(G381));
  NAND2_X1  g1029(.A1(new_n1113), .A2(new_n1143), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1204), .A2(new_n1231), .ZN(new_n1232));
  OR3_X1    g1032(.A1(new_n1232), .A2(G384), .A3(G381), .ZN(new_n1233));
  NOR3_X1   g1033(.A1(new_n1019), .A2(new_n1021), .A3(G390), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1234), .A2(new_n813), .A3(new_n1056), .A4(new_n1026), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1233), .A2(new_n1235), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n677), .A2(G213), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT125), .Z(new_n1238));
  OAI221_X1 g1038(.A(G213), .B1(new_n1232), .B2(new_n1238), .C1(new_n1233), .C2(new_n1235), .ZN(G409));
  INV_X1    g1039(.A(KEYINPUT61), .ZN(new_n1240));
  INV_X1    g1040(.A(KEYINPUT60), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n702), .B(new_n1090), .C1(new_n1227), .C2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(KEYINPUT60), .B1(new_n1206), .B2(new_n1104), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1226), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  XNOR2_X1  g1044(.A(new_n1244), .B(G384), .ZN(new_n1245));
  AND3_X1   g1045(.A1(G378), .A2(new_n1189), .A3(new_n1199), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1197), .A2(new_n967), .A3(new_n1187), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1174), .B1(new_n1185), .B2(new_n994), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1230), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1249));
  OAI211_X1 g1049(.A(new_n1237), .B(new_n1245), .C1(new_n1246), .C2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT63), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G393), .A2(G396), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1026), .A2(new_n813), .A3(new_n1056), .ZN(new_n1254));
  AND2_X1   g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n995), .A2(new_n1018), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(G390), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1256), .B1(new_n1234), .B2(new_n1259), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1257), .A2(G390), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1261), .A2(new_n1255), .A3(new_n1258), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1260), .A2(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1264), .A2(new_n1231), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(G378), .A2(new_n1189), .A3(new_n1199), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1267), .A2(KEYINPUT63), .A3(new_n1238), .A4(new_n1245), .ZN(new_n1268));
  AND4_X1   g1068(.A1(new_n1240), .A2(new_n1252), .A3(new_n1263), .A4(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n1245), .A2(new_n1238), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1237), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1271), .A2(G2897), .ZN(new_n1272));
  AOI22_X1  g1072(.A1(new_n1270), .A2(G2897), .B1(new_n1245), .B2(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(KEYINPUT126), .B1(new_n1267), .B2(new_n1237), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT126), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1275), .B(new_n1271), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1273), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(KEYINPUT127), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT127), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1279), .B(new_n1273), .C1(new_n1274), .C2(new_n1276), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1269), .A2(new_n1278), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1267), .A2(new_n1238), .ZN(new_n1282));
  AOI21_X1  g1082(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1273), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1245), .ZN(new_n1284));
  OAI21_X1  g1084(.A(KEYINPUT62), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1283), .B(new_n1285), .C1(KEYINPUT62), .C2(new_n1250), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1263), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1281), .A2(new_n1288), .ZN(G405));
  OAI211_X1 g1089(.A(new_n1284), .B(new_n1266), .C1(new_n1204), .C2(new_n1230), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1230), .B1(new_n1202), .B2(new_n1203), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1245), .B1(new_n1291), .B2(new_n1246), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  XNOR2_X1  g1093(.A(new_n1293), .B(new_n1287), .ZN(G402));
endmodule


