//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:35 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n570, new_n571, new_n572, new_n573, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1213, new_n1214, new_n1215;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT65), .B(G44), .Z(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  INV_X1    g023(.A(new_n447), .ZN(new_n449));
  NAND2_X1  g024(.A1(new_n449), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n449), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XOR2_X1   g033(.A(new_n458), .B(KEYINPUT67), .Z(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  OAI21_X1  g039(.A(G125), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  OAI211_X1 g042(.A(G137), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n468));
  AND3_X1   g043(.A1(new_n462), .A2(G101), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g047(.A(new_n472), .B(KEYINPUT68), .ZN(G160));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G2105), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  AOI21_X1  g056(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G136), .ZN(new_n483));
  MUX2_X1   g058(.A(G100), .B(G112), .S(G2105), .Z(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2104), .ZN(new_n485));
  NAND3_X1  g060(.A1(new_n481), .A2(new_n483), .A3(new_n485), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(G162));
  OAI211_X1 g062(.A(G138), .B(new_n462), .C1(new_n463), .C2(new_n464), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT4), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n478), .A2(KEYINPUT4), .A3(G138), .A4(new_n462), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n463), .C2(new_n464), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G102), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(G2105), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n497), .A2(G2104), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT69), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n497), .A2(KEYINPUT69), .A3(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n494), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n492), .A2(new_n502), .A3(KEYINPUT70), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT70), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n462), .A2(G102), .ZN(new_n505));
  AOI211_X1 g080(.A(new_n499), .B(new_n475), .C1(new_n505), .C2(new_n495), .ZN(new_n506));
  AOI21_X1  g081(.A(KEYINPUT69), .B1(new_n497), .B2(G2104), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n493), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n490), .A2(new_n491), .ZN(new_n509));
  OAI21_X1  g084(.A(new_n504), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n503), .A2(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(new_n511), .ZN(G164));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  AND2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  NOR2_X1   g089(.A1(KEYINPUT6), .A2(G651), .ZN(new_n515));
  OR2_X1    g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT5), .B(G543), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n516), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  OAI22_X1  g095(.A1(new_n513), .A2(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  AOI22_X1  g096(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n522));
  INV_X1    g097(.A(G651), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n521), .A2(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND3_X1  g101(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n527));
  XNOR2_X1  g102(.A(new_n527), .B(KEYINPUT7), .ZN(new_n528));
  INV_X1    g103(.A(G51), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n516), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n530));
  XOR2_X1   g105(.A(KEYINPUT5), .B(G543), .Z(new_n531));
  OAI221_X1 g106(.A(new_n528), .B1(new_n517), .B2(new_n529), .C1(new_n530), .C2(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n533), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n534), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(G52), .ZN(new_n537));
  INV_X1    g112(.A(G90), .ZN(new_n538));
  OAI22_X1  g113(.A1(new_n537), .A2(new_n517), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n540));
  NOR2_X1   g115(.A1(new_n540), .A2(new_n523), .ZN(new_n541));
  OR3_X1    g116(.A1(new_n539), .A2(KEYINPUT72), .A3(new_n541), .ZN(new_n542));
  OAI21_X1  g117(.A(KEYINPUT72), .B1(new_n539), .B2(new_n541), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n542), .A2(new_n543), .ZN(G171));
  AOI22_X1  g119(.A1(new_n518), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n545));
  OR2_X1    g120(.A1(new_n545), .A2(new_n523), .ZN(new_n546));
  AND2_X1   g121(.A1(new_n516), .A2(G543), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G43), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n514), .A2(new_n515), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n531), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G81), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n546), .A2(new_n548), .A3(new_n551), .ZN(new_n552));
  INV_X1    g127(.A(G860), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT73), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT75), .ZN(new_n559));
  XOR2_X1   g134(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n560));
  XNOR2_X1  g135(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n556), .A2(new_n561), .ZN(G188));
  NAND2_X1  g137(.A1(new_n547), .A2(G53), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT9), .ZN(new_n564));
  NAND2_X1  g139(.A1(G78), .A2(G543), .ZN(new_n565));
  INV_X1    g140(.A(G65), .ZN(new_n566));
  OAI21_X1  g141(.A(new_n565), .B1(new_n531), .B2(new_n566), .ZN(new_n567));
  AOI22_X1  g142(.A1(new_n567), .A2(G651), .B1(new_n550), .B2(G91), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n564), .A2(new_n568), .ZN(G299));
  INV_X1    g144(.A(KEYINPUT76), .ZN(new_n570));
  AOI21_X1  g145(.A(new_n570), .B1(new_n542), .B2(new_n543), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n542), .A2(new_n570), .A3(new_n543), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(new_n573), .ZN(G301));
  AND2_X1   g149(.A1(new_n534), .A2(new_n535), .ZN(G286));
  NAND3_X1  g150(.A1(new_n516), .A2(G49), .A3(G543), .ZN(new_n576));
  XOR2_X1   g151(.A(new_n576), .B(KEYINPUT77), .Z(new_n577));
  OR2_X1    g152(.A1(new_n518), .A2(G74), .ZN(new_n578));
  AOI22_X1  g153(.A1(G651), .A2(new_n578), .B1(new_n550), .B2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n577), .A2(new_n579), .ZN(G288));
  AOI22_X1  g155(.A1(new_n518), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n523), .ZN(new_n582));
  OR2_X1    g157(.A1(new_n582), .A2(KEYINPUT78), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n547), .A2(G48), .B1(new_n550), .B2(G86), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n582), .A2(KEYINPUT78), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  NOR2_X1   g162(.A1(new_n587), .A2(new_n523), .ZN(new_n588));
  XNOR2_X1  g163(.A(new_n588), .B(KEYINPUT79), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n547), .A2(G47), .B1(new_n550), .B2(G85), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G290));
  NAND2_X1  g166(.A1(new_n550), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n531), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(G54), .A2(new_n547), .B1(new_n596), .B2(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G301), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n601), .B2(new_n599), .ZN(G321));
  XOR2_X1   g177(.A(G321), .B(KEYINPUT80), .Z(G284));
  NAND2_X1  g178(.A1(G299), .A2(new_n599), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n599), .ZN(G280));
  XOR2_X1   g180(.A(G280), .B(KEYINPUT81), .Z(G297));
  INV_X1    g181(.A(new_n598), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NOR2_X1   g184(.A1(new_n552), .A2(G868), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n598), .A2(G559), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(new_n611), .B2(G868), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g188(.A(new_n482), .ZN(new_n614));
  OAI21_X1  g189(.A(KEYINPUT12), .B1(new_n614), .B2(new_n475), .ZN(new_n615));
  INV_X1    g190(.A(KEYINPUT12), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n482), .A2(new_n616), .A3(G2104), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT13), .ZN(new_n619));
  INV_X1    g194(.A(G2100), .ZN(new_n620));
  OR2_X1    g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n619), .A2(new_n620), .ZN(new_n622));
  MUX2_X1   g197(.A(G99), .B(G111), .S(G2105), .Z(new_n623));
  AOI22_X1  g198(.A1(new_n480), .A2(G123), .B1(G2104), .B2(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G135), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(new_n614), .ZN(new_n626));
  INV_X1    g201(.A(G2096), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n621), .A2(new_n622), .A3(new_n628), .ZN(G156));
  INV_X1    g204(.A(G14), .ZN(new_n630));
  XOR2_X1   g205(.A(G2443), .B(G2446), .Z(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2438), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2430), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AND3_X1   g210(.A1(new_n635), .A2(KEYINPUT82), .A3(KEYINPUT14), .ZN(new_n636));
  AOI21_X1  g211(.A(KEYINPUT82), .B1(new_n635), .B2(KEYINPUT14), .ZN(new_n637));
  OAI22_X1  g212(.A1(new_n636), .A2(new_n637), .B1(new_n633), .B2(new_n634), .ZN(new_n638));
  XOR2_X1   g213(.A(G2451), .B(G2454), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n638), .A2(new_n640), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n631), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g219(.A(new_n643), .ZN(new_n645));
  INV_X1    g220(.A(new_n631), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n644), .A2(new_n647), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  AOI21_X1  g226(.A(new_n630), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  AND3_X1   g227(.A1(new_n648), .A2(KEYINPUT83), .A3(new_n650), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT83), .B1(new_n648), .B2(new_n650), .ZN(new_n654));
  OAI21_X1  g229(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(G401));
  XOR2_X1   g231(.A(G2084), .B(G2090), .Z(new_n657));
  XNOR2_X1  g232(.A(G2067), .B(G2678), .ZN(new_n658));
  XNOR2_X1  g233(.A(G2072), .B(G2078), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(new_n660), .B(KEYINPUT18), .Z(new_n661));
  INV_X1    g236(.A(new_n658), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT84), .ZN(new_n663));
  AND2_X1   g238(.A1(new_n659), .A2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n659), .A2(new_n663), .ZN(new_n665));
  OAI21_X1  g240(.A(new_n662), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  INV_X1    g241(.A(new_n657), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n659), .B(KEYINPUT17), .Z(new_n668));
  OAI211_X1 g243(.A(new_n666), .B(new_n667), .C1(new_n668), .C2(new_n662), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n668), .A2(new_n662), .A3(new_n657), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n661), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(new_n627), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(G227));
  XNOR2_X1  g248(.A(G1956), .B(G2474), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n674), .B(KEYINPUT85), .ZN(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G1971), .B(G1976), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT19), .ZN(new_n679));
  NOR2_X1   g254(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT20), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n675), .A2(new_n679), .A3(new_n676), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(new_n675), .B2(new_n676), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(KEYINPUT86), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n684), .A2(new_n685), .ZN(new_n687));
  NAND3_X1  g262(.A1(new_n682), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  XOR2_X1   g263(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n689));
  INV_X1    g264(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  NOR2_X1   g267(.A1(new_n688), .A2(new_n690), .ZN(new_n693));
  XOR2_X1   g268(.A(G1991), .B(G1996), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g270(.A1(new_n692), .A2(new_n693), .A3(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT87), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n695), .B1(new_n692), .B2(new_n693), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n697), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(new_n699), .ZN(new_n702));
  INV_X1    g277(.A(new_n693), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n694), .B1(new_n703), .B2(new_n691), .ZN(new_n704));
  OAI21_X1  g279(.A(new_n702), .B1(new_n704), .B2(new_n696), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n701), .A2(new_n705), .ZN(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(G229));
  NOR2_X1   g282(.A1(G6), .A2(G16), .ZN(new_n708));
  AND3_X1   g283(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n708), .B1(new_n709), .B2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT32), .B(G1981), .Z(new_n711));
  XOR2_X1   g286(.A(new_n710), .B(new_n711), .Z(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G23), .ZN(new_n714));
  AND2_X1   g289(.A1(new_n577), .A2(new_n579), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n714), .B1(new_n715), .B2(new_n713), .ZN(new_n716));
  XNOR2_X1  g291(.A(KEYINPUT33), .B(G1976), .ZN(new_n717));
  XOR2_X1   g292(.A(new_n716), .B(new_n717), .Z(new_n718));
  NAND2_X1  g293(.A1(new_n713), .A2(G22), .ZN(new_n719));
  XOR2_X1   g294(.A(new_n719), .B(KEYINPUT88), .Z(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G303), .B2(G16), .ZN(new_n721));
  INV_X1    g296(.A(G1971), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NOR3_X1   g298(.A1(new_n712), .A2(new_n718), .A3(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n726));
  OR2_X1    g301(.A1(new_n725), .A2(KEYINPUT34), .ZN(new_n727));
  OR2_X1    g302(.A1(G16), .A2(G24), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G290), .B2(new_n713), .ZN(new_n729));
  INV_X1    g304(.A(G1986), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n482), .A2(G131), .ZN(new_n733));
  AND2_X1   g308(.A1(G107), .A2(G2105), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(G95), .B2(new_n462), .ZN(new_n735));
  INV_X1    g310(.A(G119), .ZN(new_n736));
  OAI221_X1 g311(.A(new_n733), .B1(new_n475), .B2(new_n735), .C1(new_n736), .C2(new_n479), .ZN(new_n737));
  MUX2_X1   g312(.A(G25), .B(new_n737), .S(G29), .Z(new_n738));
  XOR2_X1   g313(.A(KEYINPUT35), .B(G1991), .Z(new_n739));
  INV_X1    g314(.A(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n738), .B(new_n740), .ZN(new_n741));
  NOR3_X1   g316(.A1(new_n732), .A2(new_n741), .A3(KEYINPUT89), .ZN(new_n742));
  AND4_X1   g317(.A1(new_n726), .A2(new_n727), .A3(new_n731), .A4(new_n742), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n743), .A2(KEYINPUT36), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n607), .A2(G16), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G4), .B2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G1348), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n480), .A2(G129), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n475), .A2(G2105), .ZN(new_n750));
  AOI22_X1  g325(.A1(new_n482), .A2(G141), .B1(G105), .B2(new_n750), .ZN(new_n751));
  AND2_X1   g326(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n753));
  XNOR2_X1  g328(.A(new_n753), .B(KEYINPUT93), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT26), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n752), .A2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(G29), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n758), .B2(G32), .ZN(new_n760));
  XNOR2_X1  g335(.A(KEYINPUT27), .B(G1996), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n748), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n758), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT90), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT28), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n480), .A2(G128), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n482), .A2(G140), .ZN(new_n767));
  MUX2_X1   g342(.A(G104), .B(G116), .S(G2105), .Z(new_n768));
  NAND2_X1  g343(.A1(new_n768), .A2(G2104), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n766), .A2(new_n767), .A3(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n765), .B1(new_n771), .B2(new_n758), .ZN(new_n772));
  XNOR2_X1  g347(.A(new_n772), .B(G2067), .ZN(new_n773));
  NOR2_X1   g348(.A1(G16), .A2(G19), .ZN(new_n774));
  INV_X1    g349(.A(new_n552), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n774), .B1(new_n775), .B2(G16), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G1341), .ZN(new_n777));
  NOR3_X1   g352(.A1(new_n762), .A2(new_n773), .A3(new_n777), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT31), .B(G11), .Z(new_n779));
  XNOR2_X1  g354(.A(KEYINPUT30), .B(G28), .ZN(new_n780));
  AOI21_X1  g355(.A(new_n779), .B1(new_n758), .B2(new_n780), .ZN(new_n781));
  OAI221_X1 g356(.A(new_n781), .B1(new_n758), .B2(new_n626), .C1(new_n746), .C2(new_n747), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n713), .A2(G20), .ZN(new_n783));
  XOR2_X1   g358(.A(new_n783), .B(KEYINPUT23), .Z(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(G299), .B2(G16), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(G1956), .Z(new_n786));
  NOR2_X1   g361(.A1(new_n782), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G29), .A2(G35), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G162), .B2(G29), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT29), .ZN(new_n790));
  INV_X1    g365(.A(G2090), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NOR2_X1   g367(.A1(G5), .A2(G16), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n793), .B1(G171), .B2(G16), .ZN(new_n794));
  INV_X1    g369(.A(G1961), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n778), .A2(new_n787), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n758), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n758), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(G34), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(KEYINPUT24), .ZN(new_n803));
  NOR2_X1   g378(.A1(new_n802), .A2(KEYINPUT24), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n758), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(G160), .B2(new_n758), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(KEYINPUT92), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n801), .B1(G2084), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n713), .A2(G21), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(G168), .B2(new_n713), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT95), .ZN(new_n811));
  INV_X1    g386(.A(G1966), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NOR3_X1   g388(.A1(new_n797), .A2(new_n808), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n743), .A2(KEYINPUT36), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n750), .A2(G103), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT91), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT25), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n482), .A2(G139), .ZN(new_n819));
  AOI22_X1  g394(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n820));
  OAI211_X1 g395(.A(new_n818), .B(new_n819), .C1(new_n462), .C2(new_n820), .ZN(new_n821));
  MUX2_X1   g396(.A(G33), .B(new_n821), .S(G29), .Z(new_n822));
  XOR2_X1   g397(.A(new_n822), .B(G2072), .Z(new_n823));
  NAND2_X1  g398(.A1(new_n807), .A2(G2084), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n760), .A2(new_n761), .ZN(new_n825));
  NAND3_X1  g400(.A1(new_n823), .A2(new_n824), .A3(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT94), .Z(new_n827));
  AND4_X1   g402(.A1(new_n744), .A2(new_n814), .A3(new_n815), .A4(new_n827), .ZN(G311));
  NAND4_X1  g403(.A1(new_n744), .A2(new_n815), .A3(new_n827), .A4(new_n814), .ZN(G150));
  NAND2_X1  g404(.A1(new_n607), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT38), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n775), .A2(KEYINPUT96), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n552), .A2(new_n833), .ZN(new_n834));
  INV_X1    g409(.A(G55), .ZN(new_n835));
  INV_X1    g410(.A(G93), .ZN(new_n836));
  OAI22_X1  g411(.A1(new_n835), .A2(new_n517), .B1(new_n519), .B2(new_n836), .ZN(new_n837));
  AOI22_X1  g412(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n838));
  NOR2_X1   g413(.A1(new_n838), .A2(new_n523), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n837), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n832), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(new_n840), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n842), .A2(new_n833), .A3(new_n552), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n831), .B(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(KEYINPUT39), .ZN(new_n846));
  AOI21_X1  g421(.A(G860), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(new_n846), .B2(new_n845), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n848), .B(KEYINPUT97), .Z(new_n849));
  NOR2_X1   g424(.A1(new_n840), .A2(new_n553), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT37), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(G145));
  XNOR2_X1  g427(.A(new_n618), .B(new_n737), .ZN(new_n853));
  MUX2_X1   g428(.A(G106), .B(G118), .S(G2105), .Z(new_n854));
  AOI22_X1  g429(.A1(new_n480), .A2(G130), .B1(G2104), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(G142), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n855), .B1(new_n856), .B2(new_n614), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n853), .B(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n508), .A2(new_n509), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(new_n770), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n858), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n821), .B(new_n757), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(new_n486), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(new_n626), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n858), .A2(new_n860), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n858), .A2(new_n860), .ZN(new_n867));
  INV_X1    g442(.A(new_n862), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n863), .A2(new_n865), .A3(new_n869), .ZN(new_n870));
  INV_X1    g445(.A(G37), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n865), .ZN(new_n873));
  AND3_X1   g448(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n868), .B1(new_n866), .B2(new_n867), .ZN(new_n875));
  OAI21_X1  g450(.A(new_n873), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  OAI211_X1 g453(.A(KEYINPUT98), .B(new_n873), .C1(new_n874), .C2(new_n875), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT40), .Z(G395));
  XNOR2_X1  g456(.A(G303), .B(KEYINPUT100), .ZN(new_n882));
  OR2_X1    g457(.A1(new_n882), .A2(G305), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(G305), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n715), .B(G290), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g462(.A(new_n886), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n888), .A2(new_n883), .A3(new_n884), .ZN(new_n889));
  AND2_X1   g464(.A1(new_n887), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n593), .A2(new_n564), .A3(new_n568), .A4(new_n597), .ZN(new_n892));
  INV_X1    g467(.A(new_n892), .ZN(new_n893));
  AOI22_X1  g468(.A1(new_n593), .A2(new_n597), .B1(new_n564), .B2(new_n568), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT41), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n598), .A2(G299), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n896), .A2(new_n897), .A3(new_n892), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n895), .A2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n844), .B(new_n611), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g477(.A1(new_n893), .A2(new_n894), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(KEYINPUT99), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(KEYINPUT99), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n902), .B1(new_n906), .B2(new_n901), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n891), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n887), .A2(new_n889), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n909), .B(KEYINPUT42), .ZN(new_n910));
  INV_X1    g485(.A(new_n907), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n599), .B1(new_n908), .B2(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n842), .A2(G868), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(G295));
  NOR2_X1   g490(.A1(G295), .A2(KEYINPUT101), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT101), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n913), .A2(new_n917), .A3(new_n914), .ZN(new_n918));
  NOR2_X1   g493(.A1(new_n916), .A2(new_n918), .ZN(G331));
  NAND3_X1  g494(.A1(new_n895), .A2(KEYINPUT103), .A3(new_n898), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT103), .ZN(new_n921));
  OAI211_X1 g496(.A(new_n921), .B(KEYINPUT41), .C1(new_n893), .C2(new_n894), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n920), .A2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(G286), .B1(new_n572), .B2(new_n573), .ZN(new_n924));
  AND2_X1   g499(.A1(new_n841), .A2(new_n843), .ZN(new_n925));
  AOI21_X1  g500(.A(G168), .B1(new_n542), .B2(new_n543), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(G301), .A2(G168), .ZN(new_n928));
  INV_X1    g503(.A(new_n926), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n844), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n923), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n844), .ZN(new_n932));
  OAI21_X1  g507(.A(new_n925), .B1(new_n924), .B2(new_n926), .ZN(new_n933));
  NAND4_X1  g508(.A1(new_n932), .A2(new_n904), .A3(new_n933), .A4(new_n905), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n931), .A2(new_n890), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n899), .B1(new_n930), .B2(new_n927), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n932), .A2(new_n933), .A3(new_n903), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n936), .A2(new_n909), .A3(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n935), .A2(new_n938), .A3(new_n871), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT43), .ZN(new_n940));
  AND2_X1   g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n938), .ZN(new_n942));
  INV_X1    g517(.A(new_n937), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n900), .B1(new_n933), .B2(new_n932), .ZN(new_n944));
  OAI21_X1  g519(.A(new_n890), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(KEYINPUT102), .A3(new_n871), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT102), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n909), .B1(new_n936), .B2(new_n937), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n947), .B1(new_n948), .B2(G37), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n942), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g525(.A(new_n941), .B1(new_n950), .B2(KEYINPUT43), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n951), .A2(KEYINPUT44), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT44), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n950), .A2(new_n940), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n939), .A2(KEYINPUT43), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n953), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n952), .A2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G8), .ZN(new_n958));
  INV_X1    g533(.A(G125), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n476), .B2(new_n477), .ZN(new_n960));
  INV_X1    g535(.A(new_n466), .ZN(new_n961));
  OAI21_X1  g536(.A(G2105), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n469), .B1(new_n482), .B2(G137), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT105), .B(G40), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT106), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n962), .A2(new_n963), .A3(new_n967), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  AOI21_X1  g544(.A(G1384), .B1(new_n492), .B2(new_n502), .ZN(new_n970));
  AOI21_X1  g545(.A(new_n958), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(G1981), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n709), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n584), .A2(new_n582), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n975), .A2(G1981), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT49), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n972), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g554(.A(new_n979), .B1(new_n978), .B2(new_n977), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n715), .A2(G1976), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n982), .A2(new_n971), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT52), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n981), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT110), .B(G1976), .ZN(new_n986));
  NAND2_X1  g561(.A1(G288), .A2(new_n986), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n983), .A2(new_n984), .A3(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n983), .A2(new_n981), .A3(new_n984), .A4(new_n987), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n980), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n967), .B1(new_n472), .B2(new_n964), .ZN(new_n993));
  INV_X1    g568(.A(new_n968), .ZN(new_n994));
  INV_X1    g569(.A(G1384), .ZN(new_n995));
  OAI21_X1  g570(.A(new_n995), .B1(new_n508), .B2(new_n509), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT45), .ZN(new_n997));
  OAI22_X1  g572(.A1(new_n993), .A2(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n511), .A2(new_n995), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT104), .B(KEYINPUT45), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n998), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT108), .B1(new_n1001), .B2(G1971), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n993), .A2(new_n994), .ZN(new_n1003));
  AOI21_X1  g578(.A(KEYINPUT70), .B1(new_n492), .B2(new_n502), .ZN(new_n1004));
  NOR3_X1   g579(.A1(new_n508), .A2(new_n509), .A3(new_n504), .ZN(new_n1005));
  OAI211_X1 g580(.A(KEYINPUT50), .B(new_n995), .C1(new_n1004), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n996), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g583(.A(new_n1003), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(new_n791), .ZN(new_n1010));
  AOI22_X1  g585(.A1(new_n970), .A2(KEYINPUT45), .B1(new_n966), .B2(new_n968), .ZN(new_n1011));
  INV_X1    g586(.A(new_n1000), .ZN(new_n1012));
  AOI21_X1  g587(.A(G1384), .B1(new_n503), .B2(new_n510), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1011), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT108), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(new_n1015), .A3(new_n722), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1002), .A2(new_n1010), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(G303), .A2(G8), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n1019), .B(KEYINPUT55), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1020), .B(KEYINPUT109), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1018), .A2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n992), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(G288), .A2(G1976), .ZN(new_n1024));
  XOR2_X1   g599(.A(new_n1024), .B(KEYINPUT113), .Z(new_n1025));
  AOI22_X1  g600(.A1(new_n980), .A2(new_n1025), .B1(new_n973), .B2(new_n709), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n971), .B(KEYINPUT112), .ZN(new_n1027));
  OAI21_X1  g602(.A(new_n1023), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1020), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1018), .A2(KEYINPUT117), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT117), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1017), .A2(new_n1031), .A3(G8), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(KEYINPUT118), .B1(new_n1033), .B2(new_n991), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1032), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1031), .B1(new_n1017), .B2(G8), .ZN(new_n1036));
  OAI21_X1  g611(.A(new_n1020), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT118), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1037), .A2(new_n1038), .A3(new_n992), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT63), .ZN(new_n1040));
  INV_X1    g615(.A(G2084), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1009), .A2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g617(.A(new_n969), .B1(KEYINPUT45), .B2(new_n970), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n511), .A2(new_n995), .A3(new_n1012), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT116), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n1013), .A2(KEYINPUT116), .A3(new_n1012), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n1043), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1042), .B1(new_n1048), .B2(G1966), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  NOR4_X1   g625(.A1(new_n1022), .A2(new_n1040), .A3(G286), .A4(new_n1050), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1034), .A2(new_n1039), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n970), .A2(KEYINPUT50), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(new_n1013), .B2(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n1055));
  AND3_X1   g630(.A1(new_n1054), .A2(new_n1055), .A3(new_n969), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1055), .B1(new_n1054), .B2(new_n969), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n791), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1014), .A2(new_n722), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(KEYINPUT115), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(G8), .ZN(new_n1061));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1020), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g638(.A1(new_n1022), .A2(new_n991), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1050), .A2(G286), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1063), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1040), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1028), .B1(new_n1052), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT125), .ZN(new_n1069));
  AND2_X1   g644(.A1(new_n1006), .A2(new_n1008), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n795), .B1(new_n1070), .B2(new_n1003), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1011), .B(new_n800), .C1(new_n1012), .C2(new_n1013), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT124), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n1074));
  AND3_X1   g649(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1073), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1071), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1048), .A2(KEYINPUT123), .A3(new_n800), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1043), .ZN(new_n1079));
  AND4_X1   g654(.A1(KEYINPUT116), .A2(new_n511), .A3(new_n995), .A4(new_n1012), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT116), .B1(new_n1013), .B2(new_n1012), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n800), .B(new_n1079), .C1(new_n1080), .C2(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT123), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1074), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1077), .B1(new_n1078), .B2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1069), .B1(new_n1085), .B2(G301), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1078), .ZN(new_n1087));
  NOR2_X1   g662(.A1(new_n1009), .A2(G1961), .ZN(new_n1088));
  INV_X1    g663(.A(new_n1076), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1088), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1087), .A2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1092), .A2(KEYINPUT125), .A3(new_n601), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1088), .A2(KEYINPUT126), .ZN(new_n1094));
  NOR2_X1   g669(.A1(new_n970), .A2(new_n1012), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n472), .A2(KEYINPUT53), .A3(G40), .A4(new_n800), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g672(.A(new_n1097), .B1(new_n997), .B2(new_n996), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT126), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1099), .B1(new_n1009), .B2(G1961), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1094), .A2(new_n1098), .A3(new_n1100), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1102));
  OR3_X1    g677(.A1(new_n1101), .A2(new_n1102), .A3(new_n601), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1086), .A2(new_n1093), .A3(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT51), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G286), .A2(G8), .ZN(new_n1108));
  AOI211_X1 g683(.A(G2084), .B(new_n1003), .C1(new_n1006), .C2(new_n1008), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1079), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1109), .B1(new_n1110), .B2(new_n812), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1107), .B(new_n1108), .C1(new_n1111), .C2(new_n958), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT122), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1050), .A2(KEYINPUT122), .A3(new_n1107), .A4(new_n1108), .ZN(new_n1115));
  OAI211_X1 g690(.A(KEYINPUT51), .B(G8), .C1(new_n1049), .C2(G286), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1114), .A2(new_n1115), .A3(new_n1116), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1049), .A2(G8), .A3(G286), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g694(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1120));
  NAND2_X1  g695(.A1(G299), .A2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT119), .ZN(new_n1122));
  NOR2_X1   g697(.A1(new_n1122), .A2(KEYINPUT57), .ZN(new_n1123));
  INV_X1    g698(.A(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1121), .B1(G299), .B2(new_n1124), .ZN(new_n1125));
  XOR2_X1   g700(.A(KEYINPUT56), .B(G2072), .Z(new_n1126));
  NOR2_X1   g701(.A1(new_n1014), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g702(.A(G1956), .B1(new_n1054), .B2(new_n969), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1125), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1131));
  INV_X1    g706(.A(new_n1125), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n969), .A2(new_n970), .ZN(new_n1134));
  OAI22_X1  g709(.A1(new_n1009), .A2(G1348), .B1(G2067), .B2(new_n1134), .ZN(new_n1135));
  AND2_X1   g710(.A1(new_n1135), .A2(new_n607), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1130), .B1(new_n1133), .B2(new_n1136), .ZN(new_n1137));
  OR2_X1    g712(.A1(new_n598), .A2(KEYINPUT60), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1135), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT58), .B(G1341), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1134), .A2(new_n1141), .ZN(new_n1142));
  OAI21_X1  g717(.A(new_n1142), .B1(new_n1014), .B2(G1996), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1143), .A2(new_n1144), .A3(KEYINPUT59), .A4(new_n775), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT59), .ZN(new_n1146));
  INV_X1    g721(.A(G1996), .ZN(new_n1147));
  AOI22_X1  g722(.A1(new_n1001), .A2(new_n1147), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1148));
  NAND2_X1  g723(.A1(new_n775), .A2(new_n1144), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1146), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AND3_X1   g725(.A1(new_n1139), .A2(new_n1145), .A3(new_n1150), .ZN(new_n1151));
  OAI221_X1 g726(.A(new_n598), .B1(G2067), .B2(new_n1134), .C1(new_n1009), .C2(G1348), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT60), .B1(new_n1136), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT61), .ZN(new_n1155));
  AOI21_X1  g730(.A(KEYINPUT121), .B1(new_n1133), .B2(new_n1129), .ZN(new_n1156));
  OAI211_X1 g731(.A(new_n1151), .B(new_n1154), .C1(new_n1155), .C2(new_n1156), .ZN(new_n1157));
  AND2_X1   g732(.A1(new_n1156), .A2(new_n1155), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1137), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1087), .A2(new_n1091), .A3(G301), .ZN(new_n1160));
  OAI21_X1  g735(.A(G171), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1161));
  NAND3_X1  g736(.A1(new_n1160), .A2(new_n1161), .A3(KEYINPUT54), .ZN(new_n1162));
  AND3_X1   g737(.A1(new_n1063), .A2(new_n1162), .A3(new_n1064), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1106), .A2(new_n1119), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1086), .A2(new_n1093), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1166));
  AND3_X1   g741(.A1(new_n1117), .A2(KEYINPUT62), .A3(new_n1118), .ZN(new_n1167));
  AOI21_X1  g742(.A(KEYINPUT62), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1165), .B(new_n1166), .C1(new_n1167), .C2(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1068), .A2(new_n1164), .A3(new_n1169), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1095), .A2(new_n969), .ZN(new_n1171));
  XOR2_X1   g746(.A(new_n770), .B(G2067), .Z(new_n1172));
  NAND2_X1  g747(.A1(new_n757), .A2(new_n1147), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n756), .A2(G1996), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1175), .ZN(new_n1176));
  XNOR2_X1  g751(.A(new_n737), .B(new_n739), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1176), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(G290), .A2(G1986), .ZN(new_n1179));
  INV_X1    g754(.A(new_n1179), .ZN(new_n1180));
  NOR2_X1   g755(.A1(G290), .A2(G1986), .ZN(new_n1181));
  OR3_X1    g756(.A1(new_n1180), .A2(KEYINPUT107), .A3(new_n1181), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1171), .B1(new_n1180), .B2(KEYINPUT107), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1178), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1170), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1171), .A2(G1996), .ZN(new_n1186));
  XNOR2_X1  g761(.A(new_n1186), .B(KEYINPUT46), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1171), .B1(new_n1172), .B2(new_n757), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1187), .A2(new_n1188), .ZN(new_n1189));
  XOR2_X1   g764(.A(new_n1189), .B(KEYINPUT47), .Z(new_n1190));
  OR2_X1    g765(.A1(new_n737), .A2(new_n740), .ZN(new_n1191));
  OAI22_X1  g766(.A1(new_n1175), .A2(new_n1191), .B1(G2067), .B2(new_n770), .ZN(new_n1192));
  INV_X1    g767(.A(new_n1171), .ZN(new_n1193));
  NAND2_X1  g768(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1181), .ZN(new_n1195));
  INV_X1    g770(.A(new_n1195), .ZN(new_n1196));
  AOI21_X1  g771(.A(new_n1178), .B1(KEYINPUT48), .B2(new_n1196), .ZN(new_n1197));
  OAI21_X1  g772(.A(new_n1197), .B1(KEYINPUT48), .B2(new_n1196), .ZN(new_n1198));
  AND3_X1   g773(.A1(new_n1190), .A2(new_n1194), .A3(new_n1198), .ZN(new_n1199));
  NAND2_X1  g774(.A1(new_n1185), .A2(new_n1199), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g775(.A(KEYINPUT127), .ZN(new_n1202));
  NOR2_X1   g776(.A1(G227), .A2(new_n460), .ZN(new_n1203));
  NAND3_X1  g777(.A1(new_n706), .A2(new_n655), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g778(.A1(new_n880), .A2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g779(.A(new_n1202), .B1(new_n951), .B2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g780(.A(KEYINPUT102), .B1(new_n945), .B2(new_n871), .ZN(new_n1207));
  NOR3_X1   g781(.A1(new_n948), .A2(new_n947), .A3(G37), .ZN(new_n1208));
  OAI211_X1 g782(.A(KEYINPUT43), .B(new_n938), .C1(new_n1207), .C2(new_n1208), .ZN(new_n1209));
  INV_X1    g783(.A(new_n941), .ZN(new_n1210));
  AND4_X1   g784(.A1(new_n1202), .A2(new_n1209), .A3(new_n1210), .A4(new_n1205), .ZN(new_n1211));
  NOR2_X1   g785(.A1(new_n1206), .A2(new_n1211), .ZN(G308));
  NAND3_X1  g786(.A1(new_n1209), .A2(new_n1210), .A3(new_n1205), .ZN(new_n1213));
  NAND2_X1  g787(.A1(new_n1213), .A2(KEYINPUT127), .ZN(new_n1214));
  NAND3_X1  g788(.A1(new_n951), .A2(new_n1202), .A3(new_n1205), .ZN(new_n1215));
  NAND2_X1  g789(.A1(new_n1214), .A2(new_n1215), .ZN(G225));
endmodule


