//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 0 0 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n810, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n985, new_n986,
    new_n987, new_n989, new_n990, new_n991, new_n992, new_n994, new_n995;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G64gat), .B(G92gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n202), .B(new_n203), .Z(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(G197gat), .B(G204gat), .Z(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G211gat), .B(G218gat), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT74), .B(G211gat), .ZN(new_n209));
  AND2_X1   g008(.A1(new_n209), .A2(G218gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n207), .B(new_n208), .C1(new_n210), .C2(KEYINPUT22), .ZN(new_n211));
  INV_X1    g010(.A(new_n208), .ZN(new_n212));
  AOI21_X1  g011(.A(KEYINPUT22), .B1(new_n209), .B2(G218gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(new_n206), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G226gat), .ZN(new_n216));
  INV_X1    g015(.A(G233gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(KEYINPUT27), .B(G183gat), .ZN(new_n220));
  INV_X1    g019(.A(G190gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n222), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n223));
  INV_X1    g022(.A(G169gat), .ZN(new_n224));
  INV_X1    g023(.A(G176gat), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT70), .ZN(new_n226));
  AOI22_X1  g025(.A1(new_n226), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n227), .B1(KEYINPUT26), .B2(new_n226), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT69), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT27), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n229), .B(G183gat), .C1(new_n230), .C2(KEYINPUT68), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT68), .ZN(new_n232));
  INV_X1    g031(.A(G183gat), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n232), .B(KEYINPUT27), .C1(new_n233), .C2(KEYINPUT69), .ZN(new_n234));
  NOR2_X1   g033(.A1(KEYINPUT28), .A2(G190gat), .ZN(new_n235));
  OAI21_X1  g034(.A(KEYINPUT68), .B1(new_n230), .B2(G183gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n223), .A2(new_n228), .A3(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT23), .ZN(new_n240));
  AOI22_X1  g039(.A1(new_n240), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n241), .B1(KEYINPUT65), .B2(new_n240), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n224), .A2(new_n225), .ZN(new_n243));
  XOR2_X1   g042(.A(KEYINPUT64), .B(G176gat), .Z(new_n244));
  NOR2_X1   g043(.A1(new_n240), .A2(G169gat), .ZN(new_n245));
  AOI22_X1  g044(.A1(new_n242), .A2(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n221), .ZN(new_n249));
  NAND3_X1  g048(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n249), .A3(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT25), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT65), .ZN(new_n253));
  OAI22_X1  g052(.A1(new_n224), .A2(new_n225), .B1(new_n253), .B2(KEYINPUT23), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n240), .A2(KEYINPUT65), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n243), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT25), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n257), .B1(new_n245), .B2(new_n225), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n256), .A2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n249), .A2(new_n250), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n263));
  AOI21_X1  g062(.A(new_n260), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT67), .B1(new_n252), .B2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(new_n263), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n247), .A2(KEYINPUT66), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI211_X1 g068(.A(new_n256), .B(new_n258), .C1(new_n269), .C2(new_n260), .ZN(new_n270));
  OR2_X1    g069(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n271));
  NAND2_X1  g070(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n245), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n251), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(new_n257), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT67), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n270), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  AOI211_X1 g076(.A(new_n219), .B(new_n239), .C1(new_n266), .C2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n218), .A2(KEYINPUT29), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n270), .A2(new_n275), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(new_n238), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n215), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT75), .ZN(new_n284));
  INV_X1    g083(.A(new_n215), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n281), .A2(new_n218), .A3(new_n238), .ZN(new_n286));
  AOI21_X1  g085(.A(new_n239), .B1(new_n266), .B2(new_n277), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n285), .B(new_n286), .C1(new_n287), .C2(new_n280), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n283), .A2(new_n284), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n284), .B1(new_n283), .B2(new_n288), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n205), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n283), .A2(new_n288), .A3(new_n204), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n293), .A2(new_n294), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n292), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  XOR2_X1   g096(.A(KEYINPUT84), .B(KEYINPUT0), .Z(new_n298));
  XNOR2_X1  g097(.A(new_n298), .B(KEYINPUT85), .ZN(new_n299));
  XNOR2_X1  g098(.A(G1gat), .B(G29gat), .ZN(new_n300));
  XNOR2_X1  g099(.A(new_n299), .B(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G57gat), .B(G85gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n301), .B(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT78), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n305), .B1(new_n306), .B2(G148gat), .ZN(new_n307));
  INV_X1    g106(.A(G148gat), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n306), .A2(G148gat), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n307), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(G155gat), .A2(G162gat), .ZN(new_n312));
  INV_X1    g111(.A(G155gat), .ZN(new_n313));
  INV_X1    g112(.A(G162gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n312), .B1(new_n315), .B2(KEYINPUT2), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n311), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n308), .A2(G141gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(new_n310), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n312), .A2(KEYINPUT2), .ZN(new_n320));
  AND2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n313), .A2(new_n314), .A3(KEYINPUT77), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT76), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n312), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT77), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(G155gat), .B2(G162gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(KEYINPUT76), .A2(G155gat), .A3(G162gat), .ZN(new_n327));
  NAND4_X1  g126(.A1(new_n322), .A2(new_n324), .A3(new_n326), .A4(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n317), .B1(new_n321), .B2(new_n328), .ZN(new_n329));
  XOR2_X1   g128(.A(G127gat), .B(G134gat), .Z(new_n330));
  XNOR2_X1  g129(.A(G113gat), .B(G120gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n330), .B1(KEYINPUT1), .B2(new_n331), .ZN(new_n332));
  XOR2_X1   g131(.A(G113gat), .B(G120gat), .Z(new_n333));
  INV_X1    g132(.A(KEYINPUT1), .ZN(new_n334));
  XNOR2_X1  g133(.A(G127gat), .B(G134gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n332), .A2(new_n336), .A3(KEYINPUT79), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g137(.A(KEYINPUT79), .B1(new_n332), .B2(new_n336), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n329), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n332), .A2(new_n336), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  AND4_X1   g141(.A1(new_n326), .A2(new_n322), .A3(new_n324), .A4(new_n327), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n319), .A2(new_n320), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n343), .A2(new_n344), .B1(new_n311), .B2(new_n316), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n342), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n340), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(G225gat), .A2(G233gat), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  AOI21_X1  g148(.A(KEYINPUT83), .B1(new_n347), .B2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT83), .ZN(new_n351));
  AOI211_X1 g150(.A(new_n351), .B(new_n348), .C1(new_n340), .C2(new_n346), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT5), .B1(new_n350), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(KEYINPUT80), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT80), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT3), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n345), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n341), .A2(new_n359), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n360), .A2(new_n337), .B1(new_n329), .B2(KEYINPUT3), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n349), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT4), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n342), .A2(new_n345), .A3(new_n363), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT4), .B1(new_n329), .B2(new_n341), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT81), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n364), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n346), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(new_n367), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g170(.A1(new_n367), .A2(new_n368), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n372), .A2(KEYINPUT82), .A3(new_n362), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n353), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT5), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n364), .A2(new_n365), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n362), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(KEYINPUT6), .B(new_n304), .C1(new_n374), .C2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n304), .B1(new_n374), .B2(new_n378), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n347), .A2(new_n349), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n351), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n347), .A2(KEYINPUT83), .A3(new_n349), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n375), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n373), .ZN(new_n385));
  AOI21_X1  g184(.A(KEYINPUT82), .B1(new_n372), .B2(new_n362), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n387), .A2(new_n303), .A3(new_n377), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT6), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n380), .A2(new_n388), .A3(new_n389), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n297), .B1(new_n379), .B2(new_n390), .ZN(new_n391));
  AND2_X1   g190(.A1(new_n391), .A2(KEYINPUT35), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT86), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT29), .B1(new_n354), .B2(new_n357), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n393), .B1(new_n394), .B2(new_n215), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT29), .B1(new_n211), .B2(new_n214), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n329), .B1(new_n396), .B2(KEYINPUT3), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n394), .B2(new_n215), .ZN(new_n398));
  NAND2_X1  g197(.A1(G228gat), .A2(G233gat), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n399), .ZN(new_n401));
  OAI221_X1 g200(.A(new_n397), .B1(new_n393), .B2(new_n401), .C1(new_n394), .C2(new_n215), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(G22gat), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT87), .ZN(new_n405));
  INV_X1    g204(.A(G22gat), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n400), .A2(new_n406), .A3(new_n402), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n404), .A2(new_n405), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g207(.A(G78gat), .B(G106gat), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT31), .B(G50gat), .ZN(new_n410));
  XOR2_X1   g209(.A(new_n409), .B(new_n410), .Z(new_n411));
  NAND3_X1  g210(.A1(new_n403), .A2(KEYINPUT87), .A3(G22gat), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n408), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n404), .A2(KEYINPUT88), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT88), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n403), .A2(new_n415), .A3(G22gat), .ZN(new_n416));
  INV_X1    g215(.A(new_n411), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n414), .A2(new_n416), .A3(new_n417), .A4(new_n407), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n270), .A2(new_n275), .A3(new_n276), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n276), .B1(new_n270), .B2(new_n275), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n238), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n341), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n287), .A2(new_n342), .ZN(new_n425));
  NAND2_X1  g224(.A1(G227gat), .A2(G233gat), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT73), .B(KEYINPUT34), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(new_n428), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n424), .A2(new_n425), .A3(new_n426), .A4(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XOR2_X1   g231(.A(G71gat), .B(G99gat), .Z(new_n433));
  XNOR2_X1  g232(.A(G15gat), .B(G43gat), .ZN(new_n434));
  XNOR2_X1  g233(.A(new_n433), .B(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n426), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n287), .A2(new_n342), .ZN(new_n438));
  AOI211_X1 g237(.A(new_n341), .B(new_n239), .C1(new_n266), .C2(new_n277), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n436), .B1(new_n440), .B2(KEYINPUT32), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT33), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OR2_X1    g242(.A1(new_n435), .A2(KEYINPUT71), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n435), .A2(KEYINPUT71), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT33), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n440), .A2(KEYINPUT32), .A3(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT72), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT32), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n424), .A2(new_n425), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n437), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n452), .A2(KEYINPUT72), .A3(new_n446), .ZN(new_n453));
  AOI221_X4 g252(.A(new_n432), .B1(new_n441), .B2(new_n443), .C1(new_n449), .C2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(new_n432), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n449), .A2(new_n453), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n441), .A2(new_n443), .ZN(new_n457));
  AOI21_X1  g256(.A(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  OAI211_X1 g257(.A(new_n419), .B(new_n420), .C1(new_n454), .C2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT72), .B1(new_n452), .B2(new_n446), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n426), .B1(new_n424), .B2(new_n425), .ZN(new_n462));
  INV_X1    g261(.A(new_n446), .ZN(new_n463));
  NOR4_X1   g262(.A1(new_n462), .A2(new_n448), .A3(new_n450), .A4(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n457), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n432), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n456), .A2(new_n457), .A3(new_n455), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n420), .B1(new_n468), .B2(new_n419), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n392), .B1(new_n460), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n390), .A2(new_n379), .ZN(new_n471));
  INV_X1    g270(.A(new_n297), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n419), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AOI22_X1  g274(.A1(new_n358), .A2(new_n361), .B1(new_n365), .B2(new_n364), .ZN(new_n476));
  OR3_X1    g275(.A1(new_n476), .A2(KEYINPUT39), .A3(new_n348), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n340), .A2(new_n348), .A3(new_n346), .ZN(new_n478));
  OAI211_X1 g277(.A(KEYINPUT39), .B(new_n478), .C1(new_n476), .C2(new_n348), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n303), .A3(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT40), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n303), .A4(new_n479), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AOI21_X1  g283(.A(new_n303), .B1(new_n387), .B2(new_n377), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n486), .A2(new_n297), .B1(new_n418), .B2(new_n413), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n283), .A2(new_n488), .A3(new_n288), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n215), .B(new_n286), .C1(new_n287), .C2(new_n280), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n282), .B1(new_n287), .B2(new_n218), .ZN(new_n491));
  OAI211_X1 g290(.A(new_n490), .B(KEYINPUT37), .C1(new_n491), .C2(new_n215), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n489), .A2(new_n492), .A3(new_n205), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT38), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n288), .B1(new_n491), .B2(new_n285), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT75), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n488), .B1(new_n497), .B2(new_n289), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n489), .A2(KEYINPUT38), .A3(new_n205), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n495), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n500), .A2(new_n390), .A3(new_n379), .A4(new_n293), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n487), .A2(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n466), .A2(KEYINPUT36), .A3(new_n467), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT36), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n468), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n475), .A2(new_n502), .A3(new_n503), .A4(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n466), .A2(new_n467), .B1(new_n418), .B2(new_n413), .ZN(new_n507));
  AOI21_X1  g306(.A(KEYINPUT35), .B1(new_n507), .B2(new_n391), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n470), .A2(new_n506), .A3(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G197gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT11), .B(G169gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT12), .ZN(new_n515));
  INV_X1    g314(.A(G50gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n516), .A2(G43gat), .ZN(new_n517));
  INV_X1    g316(.A(G43gat), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(G50gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT15), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT91), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n523), .A2(G29gat), .ZN(new_n524));
  INV_X1    g323(.A(G29gat), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n526));
  OAI21_X1  g325(.A(G36gat), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n525), .A2(new_n528), .A3(KEYINPUT90), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(new_n531), .A3(KEYINPUT14), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT14), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n530), .B(new_n533), .C1(G29gat), .C2(G36gat), .ZN(new_n534));
  NAND4_X1  g333(.A1(new_n522), .A2(new_n527), .A3(new_n532), .A4(new_n534), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n519), .A3(KEYINPUT15), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(KEYINPUT15), .B1(new_n517), .B2(new_n519), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n525), .A2(KEYINPUT91), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n523), .A2(G29gat), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n528), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(new_n536), .A3(new_n532), .A4(new_n534), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n538), .A2(new_n544), .A3(KEYINPUT17), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT93), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g346(.A1(new_n538), .A2(new_n544), .A3(KEYINPUT93), .A4(KEYINPUT17), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(G8gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT16), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n551), .B1(new_n552), .B2(G1gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT92), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n550), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n553), .B1(G1gat), .B2(new_n551), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  OAI221_X1 g356(.A(new_n553), .B1(new_n554), .B2(new_n550), .C1(G1gat), .C2(new_n551), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n538), .A2(new_n544), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT17), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n549), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT94), .ZN(new_n564));
  NAND2_X1  g363(.A1(G229gat), .A2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n565), .B(KEYINPUT95), .ZN(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n559), .A2(new_n560), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT94), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n549), .A2(new_n569), .A3(new_n562), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n567), .A3(new_n568), .A4(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT18), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n515), .B1(new_n573), .B2(KEYINPUT96), .ZN(new_n574));
  AND2_X1   g373(.A1(new_n570), .A2(new_n568), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n575), .A2(KEYINPUT18), .A3(new_n567), .A4(new_n564), .ZN(new_n576));
  XOR2_X1   g375(.A(new_n559), .B(new_n560), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n566), .B(KEYINPUT13), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n573), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n571), .A2(new_n572), .B1(new_n578), .B2(new_n579), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT96), .ZN(new_n584));
  AOI21_X1  g383(.A(new_n584), .B1(new_n571), .B2(new_n572), .ZN(new_n585));
  OAI211_X1 g384(.A(new_n583), .B(new_n576), .C1(new_n585), .C2(new_n515), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(G71gat), .B(G78gat), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(new_n589), .B(KEYINPUT97), .ZN(new_n590));
  XOR2_X1   g389(.A(G57gat), .B(G64gat), .Z(new_n591));
  AOI21_X1  g390(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT97), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(KEYINPUT98), .A2(G57gat), .A3(G64gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(KEYINPUT98), .A2(G57gat), .ZN(new_n596));
  INV_X1    g395(.A(G64gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n588), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n592), .A2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT21), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(G231gat), .A2(G233gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G127gat), .B(G155gat), .ZN(new_n607));
  XOR2_X1   g406(.A(new_n607), .B(KEYINPUT99), .Z(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n606), .B(new_n609), .ZN(new_n610));
  OAI211_X1 g409(.A(new_n558), .B(new_n557), .C1(new_n602), .C2(new_n603), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n611), .B(KEYINPUT100), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n606), .B(new_n608), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G183gat), .B(G211gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n617), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n613), .A2(new_n616), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT102), .ZN(new_n625));
  XOR2_X1   g424(.A(G99gat), .B(G106gat), .Z(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G85gat), .A2(G92gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT7), .ZN(new_n629));
  NOR2_X1   g428(.A1(G85gat), .A2(G92gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(G99gat), .A2(G106gat), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(KEYINPUT8), .B2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n627), .A2(new_n629), .A3(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n627), .B1(new_n629), .B2(new_n632), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n625), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n629), .A2(new_n632), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n626), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n638), .A2(KEYINPUT102), .A3(new_n633), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g439(.A1(G232gat), .A2(G233gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(new_n640), .A2(new_n560), .B1(KEYINPUT41), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g441(.A1(new_n560), .A2(new_n561), .B1(new_n636), .B2(new_n639), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n549), .A2(new_n643), .A3(KEYINPUT103), .ZN(new_n644));
  AOI21_X1  g443(.A(KEYINPUT103), .B1(new_n549), .B2(new_n643), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G190gat), .B(G218gat), .Z(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n641), .A2(KEYINPUT41), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT101), .ZN(new_n650));
  XNOR2_X1  g449(.A(G134gat), .B(G162gat), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n650), .B(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(new_n647), .ZN(new_n653));
  OAI211_X1 g452(.A(new_n642), .B(new_n653), .C1(new_n644), .C2(new_n645), .ZN(new_n654));
  NAND3_X1  g453(.A1(new_n648), .A2(new_n652), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n652), .B1(new_n648), .B2(new_n654), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(G176gat), .B(G204gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n659), .B(new_n660), .Z(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n590), .A2(new_n591), .ZN(new_n663));
  INV_X1    g462(.A(new_n588), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  OR2_X1    g464(.A1(new_n594), .A2(new_n599), .ZN(new_n666));
  NAND4_X1  g465(.A1(new_n665), .A2(new_n666), .A3(new_n633), .A4(new_n638), .ZN(new_n667));
  OAI22_X1  g466(.A1(new_n634), .A2(new_n635), .B1(new_n592), .B2(new_n600), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(G230gat), .A2(G233gat), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n669), .A2(KEYINPUT105), .A3(new_n671), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT10), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n667), .A2(new_n668), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n636), .A2(KEYINPUT10), .A3(new_n601), .A4(new_n639), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n671), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n662), .B1(new_n676), .B2(new_n680), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n674), .A2(new_n661), .A3(new_n675), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n678), .A2(new_n679), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n671), .B1(new_n683), .B2(KEYINPUT104), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT104), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n678), .A2(new_n679), .A3(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n688), .B1(new_n682), .B2(new_n687), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n681), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n624), .A2(new_n658), .A3(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n510), .A2(new_n587), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT107), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT107), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n510), .A2(new_n697), .A3(new_n587), .A4(new_n694), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n471), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g501(.A(KEYINPUT16), .B(G8gat), .Z(new_n703));
  NAND3_X1  g502(.A1(new_n699), .A2(new_n297), .A3(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(KEYINPUT42), .ZN(new_n705));
  NOR3_X1   g504(.A1(new_n704), .A2(KEYINPUT108), .A3(new_n705), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n550), .B1(new_n699), .B2(new_n297), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n704), .B1(new_n707), .B2(new_n705), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n709));
  INV_X1    g508(.A(new_n703), .ZN(new_n710));
  AOI211_X1 g509(.A(new_n472), .B(new_n710), .C1(new_n696), .C2(new_n698), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(KEYINPUT42), .ZN(new_n712));
  AOI21_X1  g511(.A(new_n706), .B1(new_n708), .B2(new_n712), .ZN(G1325gat));
  INV_X1    g512(.A(new_n699), .ZN(new_n714));
  INV_X1    g513(.A(new_n468), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n714), .A2(G15gat), .A3(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(new_n503), .ZN(new_n717));
  AOI21_X1  g516(.A(KEYINPUT36), .B1(new_n466), .B2(new_n467), .ZN(new_n718));
  NOR2_X1   g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g518(.A(G15gat), .B1(new_n714), .B2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n716), .A2(new_n720), .ZN(G1326gat));
  NAND2_X1  g520(.A1(new_n699), .A2(new_n474), .ZN(new_n722));
  XNOR2_X1  g521(.A(KEYINPUT43), .B(G22gat), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n722), .B(new_n723), .ZN(G1327gat));
  NAND2_X1  g523(.A1(new_n510), .A2(new_n587), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n622), .A2(new_n623), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n692), .ZN(new_n727));
  NOR3_X1   g526(.A1(new_n725), .A2(new_n658), .A3(new_n727), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n728), .A2(new_n700), .A3(new_n540), .A4(new_n541), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n729), .B(KEYINPUT45), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT44), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n658), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n510), .A2(new_n732), .ZN(new_n733));
  INV_X1    g532(.A(new_n587), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n419), .B1(new_n454), .B2(new_n458), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT89), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n459), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n508), .B1(new_n738), .B2(new_n392), .ZN(new_n739));
  OAI21_X1  g538(.A(KEYINPUT109), .B1(new_n391), .B2(new_n419), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT109), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n473), .A2(new_n741), .A3(new_n474), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n719), .A2(new_n502), .A3(new_n740), .A4(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(new_n658), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n733), .B(new_n735), .C1(new_n744), .C2(KEYINPUT44), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(KEYINPUT110), .ZN(new_n746));
  INV_X1    g545(.A(new_n658), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n470), .A2(new_n509), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n740), .A2(new_n742), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI21_X1  g550(.A(new_n747), .B1(new_n748), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(new_n731), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT110), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n753), .A2(new_n754), .A3(new_n733), .A4(new_n735), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n746), .A2(new_n755), .A3(new_n700), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n756), .B1(new_n524), .B2(new_n526), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n730), .A2(new_n757), .ZN(G1328gat));
  NAND3_X1  g557(.A1(new_n728), .A2(new_n528), .A3(new_n297), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n759), .B(KEYINPUT46), .Z(new_n760));
  NAND3_X1  g559(.A1(new_n746), .A2(new_n755), .A3(new_n297), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G36gat), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(G1329gat));
  OAI21_X1  g562(.A(G43gat), .B1(new_n745), .B2(new_n719), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n728), .A2(new_n518), .A3(new_n468), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n764), .A2(KEYINPUT47), .A3(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n765), .ZN(new_n767));
  INV_X1    g566(.A(new_n719), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n746), .A2(new_n755), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n767), .B1(new_n769), .B2(G43gat), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n766), .B1(new_n770), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g570(.A(G50gat), .B1(new_n745), .B2(new_n419), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n728), .A2(new_n516), .A3(new_n474), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n772), .A2(KEYINPUT48), .A3(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(new_n773), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n746), .A2(new_n755), .A3(new_n474), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(new_n776), .B2(G50gat), .ZN(new_n777));
  XOR2_X1   g576(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n778));
  OAI21_X1  g577(.A(new_n774), .B1(new_n777), .B2(new_n778), .ZN(G1331gat));
  NAND2_X1  g578(.A1(new_n739), .A2(new_n743), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT112), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n726), .A2(new_n747), .A3(new_n587), .A4(new_n692), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n781), .B1(new_n780), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n700), .ZN(new_n786));
  XNOR2_X1  g585(.A(new_n786), .B(G57gat), .ZN(G1332gat));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n780), .A2(new_n782), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT112), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  OAI22_X1  g591(.A1(new_n792), .A2(new_n472), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n793));
  XNOR2_X1  g592(.A(KEYINPUT49), .B(G64gat), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n790), .A2(new_n297), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n788), .B1(new_n793), .B2(new_n795), .ZN(new_n796));
  NOR3_X1   g595(.A1(new_n783), .A2(new_n784), .A3(new_n472), .ZN(new_n797));
  NOR2_X1   g596(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n788), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n796), .A2(new_n800), .ZN(G1333gat));
  OAI21_X1  g600(.A(G71gat), .B1(new_n792), .B2(new_n719), .ZN(new_n802));
  INV_X1    g601(.A(G71gat), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n785), .A2(new_n803), .A3(new_n468), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n802), .A2(new_n804), .A3(KEYINPUT50), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1334gat));
  NAND2_X1  g608(.A1(new_n785), .A2(new_n474), .ZN(new_n810));
  XNOR2_X1  g609(.A(new_n810), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g610(.A1(new_n471), .A2(new_n692), .A3(G85gat), .ZN(new_n812));
  XNOR2_X1  g611(.A(new_n812), .B(KEYINPUT116), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n726), .A2(new_n734), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  OAI211_X1 g614(.A(new_n747), .B(new_n815), .C1(new_n748), .C2(new_n751), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT51), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n744), .A2(KEYINPUT51), .A3(new_n815), .ZN(new_n819));
  AND3_X1   g618(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT115), .ZN(new_n820));
  AOI21_X1  g619(.A(KEYINPUT115), .B1(new_n818), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n813), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n815), .A2(new_n691), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n823), .B(KEYINPUT114), .ZN(new_n824));
  OAI211_X1 g623(.A(new_n824), .B(new_n733), .C1(new_n744), .C2(KEYINPUT44), .ZN(new_n825));
  OAI21_X1  g624(.A(G85gat), .B1(new_n825), .B2(new_n471), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n822), .A2(new_n826), .ZN(G1336gat));
  OR2_X1    g626(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n818), .A2(new_n819), .ZN(new_n829));
  NOR3_X1   g628(.A1(new_n472), .A2(new_n692), .A3(G92gat), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G92gat), .B1(new_n825), .B2(new_n472), .ZN(new_n832));
  NAND2_X1  g631(.A1(KEYINPUT117), .A2(KEYINPUT52), .ZN(new_n833));
  AND4_X1   g632(.A1(new_n828), .A2(new_n831), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  AOI22_X1  g633(.A1(new_n829), .A2(new_n830), .B1(KEYINPUT117), .B2(KEYINPUT52), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n828), .B1(new_n835), .B2(new_n832), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n834), .A2(new_n836), .ZN(G1337gat));
  NOR3_X1   g636(.A1(new_n715), .A2(G99gat), .A3(new_n692), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n838), .B1(new_n820), .B2(new_n821), .ZN(new_n839));
  OAI21_X1  g638(.A(G99gat), .B1(new_n825), .B2(new_n719), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(G1338gat));
  NOR3_X1   g640(.A1(new_n419), .A2(new_n692), .A3(G106gat), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n829), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(G106gat), .B1(new_n825), .B2(new_n419), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g644(.A(new_n845), .B(KEYINPUT53), .ZN(G1339gat));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n661), .B1(new_n680), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n684), .A2(new_n686), .ZN(new_n849));
  OAI21_X1  g648(.A(KEYINPUT54), .B1(new_n683), .B2(new_n670), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT55), .B(new_n848), .C1(new_n849), .C2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT55), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n850), .B1(new_n684), .B2(new_n686), .ZN(new_n853));
  INV_X1    g652(.A(new_n848), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n851), .B(new_n855), .C1(new_n690), .C2(new_n689), .ZN(new_n856));
  INV_X1    g655(.A(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n587), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n583), .A2(new_n515), .A3(new_n576), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n570), .A2(new_n568), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n569), .B1(new_n549), .B2(new_n562), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n566), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  OR2_X1    g661(.A1(new_n578), .A2(new_n579), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT118), .B1(new_n864), .B2(new_n514), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT118), .ZN(new_n866));
  INV_X1    g665(.A(new_n514), .ZN(new_n867));
  AOI211_X1 g666(.A(new_n866), .B(new_n867), .C1(new_n862), .C2(new_n863), .ZN(new_n868));
  OAI211_X1 g667(.A(new_n691), .B(new_n859), .C1(new_n865), .C2(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n747), .B1(new_n858), .B2(new_n869), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n859), .B1(new_n865), .B2(new_n868), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(new_n658), .A3(new_n856), .ZN(new_n872));
  OAI21_X1  g671(.A(new_n726), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n693), .A2(new_n587), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n471), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n738), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n877), .A2(new_n297), .ZN(new_n878));
  INV_X1    g677(.A(new_n878), .ZN(new_n879));
  OR3_X1    g678(.A1(new_n879), .A2(G113gat), .A3(new_n734), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n873), .A2(new_n875), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n419), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(KEYINPUT119), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT119), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n881), .A2(new_n884), .A3(new_n419), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n883), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n471), .A2(new_n297), .ZN(new_n887));
  NAND4_X1  g686(.A1(new_n886), .A2(new_n468), .A3(new_n587), .A4(new_n887), .ZN(new_n888));
  AND3_X1   g687(.A1(new_n888), .A2(KEYINPUT120), .A3(G113gat), .ZN(new_n889));
  AOI21_X1  g688(.A(KEYINPUT120), .B1(new_n888), .B2(G113gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n880), .B1(new_n889), .B2(new_n890), .ZN(G1340gat));
  AOI21_X1  g690(.A(G120gat), .B1(new_n878), .B2(new_n691), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n886), .A2(new_n468), .A3(new_n887), .ZN(new_n893));
  INV_X1    g692(.A(new_n893), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n691), .A2(G120gat), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(G1341gat));
  OAI21_X1  g695(.A(G127gat), .B1(new_n893), .B2(new_n726), .ZN(new_n897));
  OR2_X1    g696(.A1(new_n726), .A2(G127gat), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n879), .B2(new_n898), .ZN(G1342gat));
  NOR4_X1   g698(.A1(new_n877), .A2(G134gat), .A3(new_n297), .A4(new_n658), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(KEYINPUT56), .ZN(new_n901));
  OAI21_X1  g700(.A(G134gat), .B1(new_n893), .B2(new_n658), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1343gat));
  NAND4_X1  g702(.A1(new_n881), .A2(KEYINPUT121), .A3(KEYINPUT57), .A4(new_n474), .ZN(new_n904));
  AND2_X1   g703(.A1(new_n719), .A2(new_n887), .ZN(new_n905));
  INV_X1    g704(.A(new_n869), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n856), .B1(new_n586), .B2(new_n582), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n658), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n871), .A2(new_n658), .A3(new_n856), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n624), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  OAI211_X1 g709(.A(KEYINPUT57), .B(new_n474), .C1(new_n910), .C2(new_n874), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT121), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g712(.A(KEYINPUT57), .B1(new_n881), .B2(new_n474), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n904), .B(new_n905), .C1(new_n913), .C2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G141gat), .B1(new_n915), .B2(new_n734), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT122), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n876), .A2(new_n474), .A3(new_n719), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n919), .A2(new_n297), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n920), .A2(new_n306), .A3(new_n587), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n918), .A2(new_n922), .A3(KEYINPUT58), .ZN(new_n923));
  INV_X1    g722(.A(KEYINPUT58), .ZN(new_n924));
  OAI211_X1 g723(.A(new_n916), .B(new_n921), .C1(new_n917), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(G1344gat));
  NAND2_X1  g725(.A1(new_n308), .A2(KEYINPUT59), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n927), .B1(new_n920), .B2(new_n691), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n915), .A2(new_n692), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n930), .B1(new_n747), .B2(new_n857), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n658), .A2(KEYINPUT123), .A3(new_n856), .ZN(new_n932));
  NOR3_X1   g731(.A1(new_n931), .A2(new_n871), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n726), .B1(new_n933), .B2(new_n870), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n419), .B1(new_n934), .B2(new_n875), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n911), .B1(new_n935), .B2(KEYINPUT57), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n936), .A2(new_n719), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n887), .A2(KEYINPUT59), .A3(new_n691), .ZN(new_n938));
  OAI22_X1  g737(.A1(new_n929), .A2(KEYINPUT59), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n928), .B1(new_n939), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g739(.A(G155gat), .B1(new_n915), .B2(new_n726), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n920), .A2(new_n313), .A3(new_n624), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n941), .A2(new_n942), .ZN(G1346gat));
  OAI21_X1  g742(.A(G162gat), .B1(new_n915), .B2(new_n658), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n747), .A2(new_n314), .A3(new_n472), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n944), .B1(new_n919), .B2(new_n945), .ZN(G1347gat));
  AOI21_X1  g745(.A(new_n700), .B1(new_n873), .B2(new_n875), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n472), .B1(new_n737), .B2(new_n459), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(G169gat), .B1(new_n950), .B2(new_n587), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n700), .A2(new_n472), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n952), .A2(new_n468), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n953), .B1(new_n883), .B2(new_n885), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n734), .A2(new_n224), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n951), .B1(new_n954), .B2(new_n955), .ZN(G1348gat));
  NOR2_X1   g755(.A1(new_n692), .A2(new_n244), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n225), .B1(new_n949), .B2(new_n692), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g759(.A(new_n960), .B(KEYINPUT124), .ZN(G1349gat));
  NAND2_X1  g760(.A1(new_n624), .A2(new_n220), .ZN(new_n962));
  OR3_X1    g761(.A1(new_n949), .A2(KEYINPUT125), .A3(new_n962), .ZN(new_n963));
  OAI21_X1  g762(.A(KEYINPUT125), .B1(new_n949), .B2(new_n962), .ZN(new_n964));
  NAND2_X1  g763(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g764(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g765(.A(new_n233), .B1(new_n954), .B2(new_n624), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT60), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT60), .ZN(new_n969));
  AND2_X1   g768(.A1(new_n954), .A2(new_n624), .ZN(new_n970));
  OAI211_X1 g769(.A(new_n969), .B(new_n965), .C1(new_n970), .C2(new_n233), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n968), .A2(new_n971), .ZN(G1350gat));
  AOI21_X1  g771(.A(new_n221), .B1(new_n954), .B2(new_n747), .ZN(new_n973));
  OR2_X1    g772(.A1(new_n973), .A2(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(KEYINPUT61), .ZN(new_n975));
  NOR3_X1   g774(.A1(new_n949), .A2(G190gat), .A3(new_n658), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT126), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n974), .A2(new_n975), .A3(new_n977), .ZN(G1351gat));
  XNOR2_X1  g777(.A(KEYINPUT127), .B(G197gat), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n936), .A2(new_n719), .A3(new_n952), .ZN(new_n980));
  OAI21_X1  g779(.A(new_n979), .B1(new_n980), .B2(new_n734), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n947), .A2(new_n297), .A3(new_n474), .A4(new_n719), .ZN(new_n982));
  OR2_X1    g781(.A1(new_n734), .A2(new_n979), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(G1352gat));
  NOR3_X1   g783(.A1(new_n982), .A2(G204gat), .A3(new_n692), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT62), .ZN(new_n986));
  OAI21_X1  g785(.A(G204gat), .B1(new_n980), .B2(new_n692), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1353gat));
  OR3_X1    g787(.A1(new_n982), .A2(new_n209), .A3(new_n726), .ZN(new_n989));
  NAND4_X1  g788(.A1(new_n936), .A2(new_n719), .A3(new_n624), .A4(new_n952), .ZN(new_n990));
  AND3_X1   g789(.A1(new_n990), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n991));
  AOI21_X1  g790(.A(KEYINPUT63), .B1(new_n990), .B2(G211gat), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n989), .B1(new_n991), .B2(new_n992), .ZN(G1354gat));
  OAI21_X1  g792(.A(G218gat), .B1(new_n980), .B2(new_n658), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n658), .A2(G218gat), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n994), .B1(new_n982), .B2(new_n995), .ZN(G1355gat));
endmodule


