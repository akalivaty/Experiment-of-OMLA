//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:37 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1260, new_n1261,
    new_n1262, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1318, new_n1319, new_n1320;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  AOI22_X1  g0008(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n210));
  AND2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OR2_X1    g0011(.A1(new_n211), .A2(KEYINPUT66), .ZN(new_n212));
  NAND3_X1  g0012(.A1(new_n209), .A2(new_n210), .A3(KEYINPUT66), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G20), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OR2_X1    g0018(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g0019(.A(KEYINPUT64), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n201), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n222));
  NAND3_X1  g0022(.A1(new_n221), .A2(G50), .A3(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  NAND2_X1  g0024(.A1(G1), .A2(G13), .ZN(new_n225));
  INV_X1    g0025(.A(G20), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n217), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n219), .A2(new_n228), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n218), .ZN(G361));
  XOR2_X1   g0033(.A(G238), .B(G244), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT68), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT67), .B(KEYINPUT2), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  INV_X1    g0044(.A(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(KEYINPUT69), .B(G50), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XOR2_X1   g0049(.A(G107), .B(G116), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n225), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT8), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(G58), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n245), .A2(KEYINPUT8), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT72), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n256), .A2(KEYINPUT72), .A3(G58), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(G20), .A2(G33), .ZN(new_n267));
  AOI22_X1  g0067(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n255), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g0069(.A1(KEYINPUT70), .A2(G1), .ZN(new_n270));
  NOR2_X1   g0070(.A1(KEYINPUT70), .A2(G1), .ZN(new_n271));
  NOR2_X1   g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G20), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n273), .A2(G50), .A3(new_n255), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT70), .ZN(new_n275));
  INV_X1    g0075(.A(G1), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g0077(.A1(KEYINPUT70), .A2(G1), .ZN(new_n278));
  NAND4_X1  g0078(.A1(new_n277), .A2(G13), .A3(G20), .A4(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n274), .B1(G50), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n269), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G41), .ZN(new_n283));
  INV_X1    g0083(.A(G45), .ZN(new_n284));
  AOI21_X1  g0084(.A(G1), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n285), .A2(new_n287), .A3(G274), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n225), .B1(G33), .B2(G41), .ZN(new_n289));
  NOR2_X1   g0089(.A1(G41), .A2(G45), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n272), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n288), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(KEYINPUT3), .B(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(G1698), .ZN(new_n297));
  INV_X1    g0097(.A(G223), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  OAI22_X1  g0099(.A1(new_n297), .A2(new_n298), .B1(new_n299), .B2(new_n296), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  AND3_X1   g0101(.A1(new_n296), .A2(G222), .A3(new_n301), .ZN(new_n302));
  OR2_X1    g0102(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n303), .A2(KEYINPUT71), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n287), .B1(new_n303), .B2(KEYINPUT71), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n282), .B1(new_n306), .B2(G169), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(KEYINPUT73), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT73), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n309), .B(new_n282), .C1(new_n306), .C2(G169), .ZN(new_n310));
  INV_X1    g0110(.A(G179), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n306), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n310), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n282), .A2(KEYINPUT77), .A3(KEYINPUT9), .ZN(new_n314));
  OR2_X1    g0114(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n315));
  NAND2_X1  g0115(.A1(KEYINPUT77), .A2(KEYINPUT9), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n281), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n314), .A2(new_n317), .B1(new_n306), .B2(G190), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT10), .ZN(new_n319));
  INV_X1    g0119(.A(G200), .ZN(new_n320));
  OR2_X1    g0120(.A1(new_n306), .A2(new_n320), .ZN(new_n321));
  AND3_X1   g0121(.A1(new_n318), .A2(new_n319), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n319), .B1(new_n318), .B2(new_n321), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n313), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  AND3_X1   g0124(.A1(new_n285), .A2(new_n287), .A3(G274), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n325), .B1(new_n292), .B2(G232), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G33), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n327), .A2(new_n329), .A3(G223), .A4(new_n301), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n327), .A2(new_n329), .A3(G226), .A4(G1698), .ZN(new_n331));
  NAND2_X1  g0131(.A1(G33), .A2(G87), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(new_n289), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n326), .A2(new_n311), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(G169), .B1(new_n326), .B2(new_n334), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n327), .A2(new_n329), .ZN(new_n338));
  AOI21_X1  g0138(.A(KEYINPUT7), .B1(new_n338), .B2(new_n226), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT7), .ZN(new_n340));
  AOI211_X1 g0140(.A(new_n340), .B(G20), .C1(new_n327), .C2(new_n329), .ZN(new_n341));
  OAI21_X1  g0141(.A(G68), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  XNOR2_X1  g0142(.A(G58), .B(G68), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(G20), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT81), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n267), .A2(new_n345), .A3(G159), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n345), .B1(new_n267), .B2(G159), .ZN(new_n348));
  OAI21_X1  g0148(.A(new_n344), .B1(new_n347), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT16), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n342), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G68), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n340), .B1(new_n296), .B2(G20), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n328), .A2(G33), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n356));
  OAI211_X1 g0156(.A(KEYINPUT7), .B(new_n226), .C1(new_n355), .C2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n353), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  OAI21_X1  g0158(.A(KEYINPUT16), .B1(new_n358), .B2(new_n349), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n255), .B1(new_n352), .B2(new_n359), .ZN(new_n360));
  NOR3_X1   g0160(.A1(new_n270), .A2(new_n271), .A3(new_n226), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n261), .B(new_n260), .C1(new_n361), .C2(new_n254), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n262), .A2(new_n279), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n362), .A2(new_n363), .A3(KEYINPUT82), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT82), .B1(new_n362), .B2(new_n363), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n337), .B1(new_n360), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT18), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT18), .ZN(new_n369));
  OAI211_X1 g0169(.A(new_n337), .B(new_n369), .C1(new_n360), .C2(new_n366), .ZN(new_n370));
  AND2_X1   g0170(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n351), .B1(new_n342), .B2(new_n350), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n358), .A2(KEYINPUT16), .A3(new_n349), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n254), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OR2_X1    g0174(.A1(new_n364), .A2(new_n365), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n326), .A2(new_n376), .A3(new_n334), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n277), .A2(new_n278), .ZN(new_n378));
  OAI211_X1 g0178(.A(G232), .B(new_n287), .C1(new_n378), .C2(new_n290), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n288), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n380), .B1(new_n289), .B2(new_n333), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n377), .B1(new_n381), .B2(G200), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n374), .A2(new_n375), .A3(new_n382), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT83), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT17), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n374), .A2(new_n375), .A3(new_n382), .A4(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n385), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(new_n279), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n299), .ZN(new_n393));
  XNOR2_X1  g0193(.A(new_n393), .B(KEYINPUT75), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n279), .A2(new_n255), .A3(KEYINPUT76), .ZN(new_n395));
  INV_X1    g0195(.A(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(KEYINPUT76), .B1(new_n279), .B2(new_n255), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n398), .A2(G77), .A3(new_n273), .ZN(new_n399));
  NAND2_X1  g0199(.A1(G20), .A2(G77), .ZN(new_n400));
  AND2_X1   g0200(.A1(new_n257), .A2(new_n258), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n226), .A2(new_n264), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n400), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  XNOR2_X1  g0203(.A(KEYINPUT15), .B(G87), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n403), .B1(new_n265), .B2(new_n405), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n394), .B(new_n399), .C1(new_n255), .C2(new_n406), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n296), .A2(G232), .A3(new_n301), .ZN(new_n408));
  INV_X1    g0208(.A(G238), .ZN(new_n409));
  OAI221_X1 g0209(.A(new_n408), .B1(new_n206), .B2(new_n296), .C1(new_n297), .C2(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(new_n289), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n325), .B1(new_n292), .B2(G244), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n411), .A2(new_n311), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n412), .ZN(new_n414));
  INV_X1    g0214(.A(G169), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n407), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n414), .A2(new_n376), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n407), .B1(new_n418), .B2(KEYINPUT74), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT74), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n420), .B1(new_n414), .B2(G200), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n419), .B1(new_n418), .B2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n371), .A2(new_n391), .A3(new_n417), .A4(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n267), .A2(G50), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n353), .A2(G20), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n226), .A2(G33), .ZN(new_n426));
  OAI211_X1 g0226(.A(new_n424), .B(new_n425), .C1(new_n299), .C2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT11), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n427), .A2(new_n428), .A3(new_n254), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n427), .B2(new_n254), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT12), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n392), .B2(new_n353), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n279), .A2(KEYINPUT12), .A3(G68), .ZN(new_n433));
  OAI22_X1  g0233(.A1(new_n429), .A2(new_n430), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(new_n397), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n435), .A2(G68), .A3(new_n273), .A4(new_n395), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n436), .A2(KEYINPUT79), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT79), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n398), .A2(new_n438), .A3(G68), .A4(new_n273), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n434), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n325), .B1(new_n292), .B2(G238), .ZN(new_n441));
  INV_X1    g0241(.A(KEYINPUT13), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n327), .A2(new_n329), .A3(G232), .A4(G1698), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n327), .A2(new_n329), .A3(G226), .A4(new_n301), .ZN(new_n444));
  AND3_X1   g0244(.A1(KEYINPUT78), .A2(G33), .A3(G97), .ZN(new_n445));
  AOI21_X1  g0245(.A(KEYINPUT78), .B1(G33), .B2(G97), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n443), .A2(new_n444), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n289), .ZN(new_n449));
  AND3_X1   g0249(.A1(new_n441), .A2(new_n442), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n442), .B1(new_n441), .B2(new_n449), .ZN(new_n451));
  NOR3_X1   g0251(.A1(new_n450), .A2(new_n451), .A3(G190), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n441), .A2(new_n449), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT13), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n441), .A2(new_n442), .A3(new_n449), .ZN(new_n455));
  AOI21_X1  g0255(.A(G200), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n440), .B1(new_n452), .B2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT80), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n320), .B1(new_n450), .B2(new_n451), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n454), .A2(new_n455), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(G190), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT80), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n461), .A2(new_n462), .A3(new_n440), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g0264(.A(G169), .B1(new_n450), .B2(new_n451), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(KEYINPUT14), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT14), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n460), .A2(new_n467), .A3(G169), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n454), .A2(G179), .A3(new_n455), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n466), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  INV_X1    g0270(.A(new_n440), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n464), .A2(new_n472), .ZN(new_n473));
  NOR3_X1   g0273(.A1(new_n324), .A2(new_n423), .A3(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n327), .A2(new_n329), .A3(G238), .A4(new_n301), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(KEYINPUT87), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT87), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n296), .A2(new_n478), .A3(G238), .A4(new_n301), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n296), .A2(G244), .A3(G1698), .ZN(new_n480));
  NAND2_X1  g0280(.A1(G33), .A2(G116), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n477), .A2(new_n479), .A3(new_n480), .A4(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n289), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n277), .A2(G45), .A3(new_n278), .ZN(new_n484));
  OR2_X1    g0284(.A1(new_n484), .A2(G274), .ZN(new_n485));
  INV_X1    g0285(.A(G250), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n289), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND3_X1   g0288(.A1(new_n483), .A2(G190), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n320), .B1(new_n483), .B2(new_n488), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n279), .A2(new_n255), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT84), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n492), .B1(new_n378), .B2(new_n264), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n272), .A2(KEYINPUT84), .A3(G33), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n491), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n495), .A2(G87), .ZN(new_n496));
  OAI21_X1  g0296(.A(KEYINPUT19), .B1(new_n445), .B2(new_n446), .ZN(new_n497));
  INV_X1    g0297(.A(G87), .ZN(new_n498));
  INV_X1    g0298(.A(new_n207), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n497), .A2(new_n226), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n296), .A2(new_n226), .A3(G68), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT19), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n426), .B2(new_n205), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n254), .B1(new_n500), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n405), .A2(new_n279), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n496), .A2(new_n505), .A3(new_n507), .ZN(new_n508));
  NOR3_X1   g0308(.A1(new_n489), .A2(new_n490), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n483), .A2(new_n488), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n510), .A2(G179), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT88), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n493), .A2(new_n494), .ZN(new_n513));
  INV_X1    g0313(.A(new_n491), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n513), .A2(new_n514), .A3(new_n405), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n505), .A2(new_n515), .A3(new_n507), .ZN(new_n516));
  AOI22_X1  g0316(.A1(new_n482), .A2(new_n289), .B1(new_n485), .B2(new_n487), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(G169), .B2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT88), .B1(new_n517), .B2(new_n311), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n509), .B1(new_n512), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n279), .A2(G97), .ZN(new_n522));
  AOI21_X1  g0322(.A(new_n522), .B1(new_n495), .B2(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n267), .A2(G77), .ZN(new_n524));
  INV_X1    g0324(.A(KEYINPUT6), .ZN(new_n525));
  NOR3_X1   g0325(.A1(new_n525), .A2(new_n205), .A3(G107), .ZN(new_n526));
  XNOR2_X1  g0326(.A(G97), .B(G107), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n526), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n524), .B1(new_n528), .B2(new_n226), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n206), .B1(new_n354), .B2(new_n357), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n254), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g0331(.A1(new_n523), .A2(new_n531), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n327), .A2(new_n329), .A3(G244), .A4(new_n301), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT85), .ZN(new_n534));
  OR2_X1    g0334(.A1(new_n534), .A2(KEYINPUT4), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n533), .A2(new_n536), .ZN(new_n537));
  NAND4_X1  g0337(.A1(new_n296), .A2(G244), .A3(new_n535), .A4(new_n301), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n296), .A2(G250), .A3(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G283), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n537), .A2(new_n538), .A3(new_n539), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n289), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n270), .A2(new_n271), .A3(new_n284), .ZN(new_n543));
  XNOR2_X1  g0343(.A(KEYINPUT5), .B(G41), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(G274), .A3(new_n287), .A4(new_n544), .ZN(new_n545));
  AND2_X1   g0345(.A1(KEYINPUT5), .A2(G41), .ZN(new_n546));
  NOR2_X1   g0346(.A1(KEYINPUT5), .A2(G41), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(G257), .B(new_n287), .C1(new_n484), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n545), .A2(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n542), .A2(new_n376), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(G200), .B1(new_n542), .B2(new_n551), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n532), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n542), .A2(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n415), .ZN(new_n556));
  AOI21_X1  g0356(.A(new_n550), .B1(new_n289), .B2(new_n541), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(new_n311), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n523), .A2(new_n531), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n554), .A2(KEYINPUT86), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g0361(.A(KEYINPUT86), .B1(new_n554), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n521), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n327), .A2(new_n329), .A3(new_n226), .A4(G87), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n564), .A2(KEYINPUT22), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT22), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n296), .A2(new_n566), .A3(new_n226), .A4(G87), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n226), .B2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n265), .A2(G116), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g0374(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT90), .ZN(new_n577));
  INV_X1    g0377(.A(KEYINPUT24), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n574), .B1(new_n565), .B2(new_n567), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT90), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(KEYINPUT24), .B1(new_n580), .B2(KEYINPUT90), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n254), .B(new_n579), .C1(new_n582), .C2(new_n583), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n327), .A2(new_n329), .A3(G257), .A4(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n327), .A2(new_n329), .A3(G250), .A4(new_n301), .ZN(new_n586));
  INV_X1    g0386(.A(G294), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n264), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n289), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n289), .B1(new_n543), .B2(new_n544), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(G264), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n591), .A3(new_n545), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n320), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n289), .A2(new_n588), .B1(new_n590), .B2(G264), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n594), .A2(new_n376), .A3(new_n545), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n279), .A2(G107), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n597), .B(KEYINPUT25), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n495), .A2(G107), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n584), .A2(new_n596), .A3(new_n601), .ZN(new_n602));
  NOR2_X1   g0402(.A1(new_n580), .A2(KEYINPUT90), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n255), .B1(new_n603), .B2(new_n578), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n576), .A2(new_n577), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n605), .A2(KEYINPUT24), .A3(new_n581), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n600), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n592), .A2(new_n415), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n594), .A2(new_n311), .A3(new_n545), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n602), .B1(new_n607), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(G116), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n361), .A2(G13), .A3(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n253), .A2(new_n225), .B1(G20), .B2(new_n612), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n540), .B(new_n226), .C1(G33), .C2(new_n205), .ZN(new_n615));
  AND3_X1   g0415(.A1(new_n614), .A2(KEYINPUT20), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(KEYINPUT20), .B1(new_n614), .B2(new_n615), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n612), .B1(new_n493), .B2(new_n494), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n618), .B1(new_n398), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(G270), .B(new_n287), .C1(new_n484), .C2(new_n548), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n545), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n327), .A2(new_n329), .A3(G264), .A4(G1698), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n327), .A2(new_n329), .A3(G257), .A4(new_n301), .ZN(new_n624));
  INV_X1    g0424(.A(G303), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n296), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(new_n289), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(G179), .A3(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(KEYINPUT89), .B1(new_n620), .B2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n619), .A2(new_n435), .A3(new_n395), .ZN(new_n630));
  INV_X1    g0430(.A(new_n617), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n614), .A2(KEYINPUT20), .A3(new_n615), .ZN(new_n632));
  AOI22_X1  g0432(.A1(new_n631), .A2(new_n632), .B1(new_n612), .B2(new_n392), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n630), .A2(new_n633), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT89), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n545), .A2(new_n621), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n636), .B1(new_n289), .B2(new_n626), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n634), .A2(new_n635), .A3(new_n637), .A4(G179), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n629), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT21), .ZN(new_n640));
  INV_X1    g0440(.A(new_n627), .ZN(new_n641));
  OAI21_X1  g0441(.A(G169), .B1(new_n641), .B2(new_n636), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n640), .B1(new_n642), .B2(new_n620), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n622), .A2(new_n627), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n634), .A2(new_n644), .A3(KEYINPUT21), .A4(G169), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(G200), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n646), .B(new_n620), .C1(new_n376), .C2(new_n644), .ZN(new_n647));
  NAND4_X1  g0447(.A1(new_n639), .A2(new_n643), .A3(new_n645), .A4(new_n647), .ZN(new_n648));
  NOR4_X1   g0448(.A1(new_n475), .A2(new_n563), .A3(new_n611), .A4(new_n648), .ZN(G372));
  INV_X1    g0449(.A(new_n313), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n322), .A2(new_n323), .ZN(new_n651));
  INV_X1    g0451(.A(new_n417), .ZN(new_n652));
  AOI22_X1  g0452(.A1(new_n471), .A2(new_n470), .B1(new_n652), .B2(new_n457), .ZN(new_n653));
  AND2_X1   g0453(.A1(new_n385), .A2(new_n390), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n371), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g0455(.A(new_n650), .B1(new_n651), .B2(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n518), .A2(new_n511), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n610), .B1(new_n584), .B2(new_n601), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n643), .A2(new_n645), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  AOI21_X1  g0462(.A(KEYINPUT92), .B1(new_n662), .B2(new_n639), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n629), .A2(new_n638), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT92), .ZN(new_n665));
  NOR3_X1   g0465(.A1(new_n664), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n660), .B1(new_n663), .B2(new_n666), .ZN(new_n667));
  AND3_X1   g0467(.A1(new_n556), .A2(new_n559), .A3(new_n558), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n555), .A2(new_n320), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n557), .A2(new_n376), .ZN(new_n670));
  AOI21_X1  g0470(.A(new_n559), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n489), .A2(new_n490), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT91), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n505), .A2(new_n507), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n674), .B1(new_n675), .B2(new_n496), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n508), .A2(KEYINPUT91), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n673), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  AND4_X1   g0478(.A1(new_n672), .A2(new_n602), .A3(new_n657), .A4(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n658), .B1(new_n667), .B2(new_n679), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n657), .A3(new_n668), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT26), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(KEYINPUT93), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n521), .A2(KEYINPUT26), .A3(new_n668), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT93), .ZN(new_n686));
  NAND3_X1  g0486(.A1(new_n681), .A2(new_n686), .A3(new_n682), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n685), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n656), .B1(new_n475), .B2(new_n690), .ZN(G369));
  NAND3_X1  g0491(.A1(new_n662), .A2(KEYINPUT92), .A3(new_n639), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n665), .B1(new_n664), .B2(new_n661), .ZN(new_n693));
  INV_X1    g0493(.A(G13), .ZN(new_n694));
  NOR2_X1   g0494(.A1(new_n694), .A2(G20), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n272), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(G213), .B1(new_n696), .B2(KEYINPUT27), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n696), .A2(KEYINPUT27), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT94), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g0500(.A1(new_n696), .A2(KEYINPUT94), .A3(KEYINPUT27), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n697), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  XOR2_X1   g0502(.A(KEYINPUT95), .B(G343), .Z(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n702), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n620), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n692), .A2(new_n693), .A3(new_n706), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n707), .B1(new_n648), .B2(new_n706), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n584), .A2(new_n596), .A3(new_n601), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n711), .A2(new_n659), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n712), .B1(new_n607), .B2(new_n705), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n713), .B1(new_n660), .B2(new_n705), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n710), .A2(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n705), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n716), .B1(new_n662), .B2(new_n639), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n717), .A2(new_n712), .B1(new_n659), .B2(new_n705), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n715), .A2(new_n718), .ZN(G399));
  INV_X1    g0519(.A(new_n229), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(G41), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n499), .A2(new_n498), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n723), .A2(G116), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n722), .A2(G1), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n224), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n722), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n660), .A2(new_n662), .A3(new_n639), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n658), .B1(new_n679), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n520), .A2(new_n512), .ZN(new_n731));
  INV_X1    g0531(.A(new_n509), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n731), .A2(new_n732), .A3(new_n668), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n682), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n734), .B1(new_n682), .B2(new_n681), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n730), .A2(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n736), .A2(KEYINPUT29), .A3(new_n705), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n716), .B1(new_n680), .B2(new_n688), .ZN(new_n738));
  XNOR2_X1  g0538(.A(KEYINPUT96), .B(KEYINPUT29), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n737), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n648), .A2(new_n611), .ZN(new_n742));
  INV_X1    g0542(.A(KEYINPUT86), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n743), .B1(new_n668), .B2(new_n671), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n554), .A2(KEYINPUT86), .A3(new_n560), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND4_X1  g0546(.A1(new_n742), .A2(new_n521), .A3(new_n746), .A4(new_n705), .ZN(new_n747));
  INV_X1    g0547(.A(KEYINPUT30), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n557), .A2(new_n637), .A3(G179), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n517), .A2(new_n594), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n748), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n555), .A2(new_n628), .ZN(new_n752));
  AND3_X1   g0552(.A1(new_n594), .A2(new_n483), .A3(new_n488), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(KEYINPUT30), .A3(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(G179), .B1(new_n622), .B2(new_n627), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n510), .A2(new_n755), .A3(new_n555), .A4(new_n592), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n751), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(new_n716), .ZN(new_n758));
  INV_X1    g0558(.A(KEYINPUT31), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n757), .A2(KEYINPUT31), .A3(new_n716), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n747), .A2(new_n760), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n762), .A2(G330), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n741), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n728), .B1(new_n765), .B2(G1), .ZN(new_n766));
  XOR2_X1   g0566(.A(new_n766), .B(KEYINPUT97), .Z(G364));
  XNOR2_X1  g0567(.A(new_n695), .B(KEYINPUT98), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(G45), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G1), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n721), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n708), .A2(G330), .ZN(new_n772));
  NOR3_X1   g0572(.A1(new_n710), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n773), .B(KEYINPUT99), .ZN(new_n774));
  NOR2_X1   g0574(.A1(G13), .A2(G33), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(G20), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n708), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(G20), .B1(KEYINPUT100), .B2(G169), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g0581(.A1(KEYINPUT100), .A2(G169), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n225), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n783), .A2(new_n777), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n248), .A2(G45), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n720), .A2(new_n296), .ZN(new_n787));
  OAI211_X1 g0587(.A(new_n786), .B(new_n787), .C1(G45), .C2(new_n726), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n720), .A2(new_n338), .ZN(new_n789));
  AOI22_X1  g0589(.A1(new_n789), .A2(G355), .B1(new_n612), .B2(new_n720), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n785), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  INV_X1    g0591(.A(new_n783), .ZN(new_n792));
  INV_X1    g0592(.A(KEYINPUT101), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n793), .B1(new_n226), .B2(G190), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n376), .A2(KEYINPUT101), .A3(G20), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n320), .A2(G179), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n794), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G107), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n226), .A2(new_n311), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n800), .A2(G200), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(G190), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n801), .A2(new_n376), .ZN(new_n803));
  AOI22_X1  g0603(.A1(new_n802), .A2(G68), .B1(new_n803), .B2(G50), .ZN(new_n804));
  NAND3_X1  g0604(.A1(new_n800), .A2(G190), .A3(new_n320), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n338), .B1(new_n806), .B2(G58), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n796), .A2(G20), .A3(G190), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  NOR2_X1   g0609(.A1(G190), .A2(G200), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n800), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G87), .A2(new_n809), .B1(new_n812), .B2(G77), .ZN(new_n813));
  AND4_X1   g0613(.A1(new_n799), .A2(new_n804), .A3(new_n807), .A4(new_n813), .ZN(new_n814));
  NOR2_X1   g0614(.A1(G179), .A2(G200), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n226), .B1(new_n815), .B2(G190), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n816), .B(KEYINPUT102), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n794), .A2(new_n815), .A3(new_n795), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G159), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n817), .A2(G97), .B1(new_n820), .B2(KEYINPUT32), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n814), .B(new_n821), .C1(KEYINPUT32), .C2(new_n820), .ZN(new_n822));
  INV_X1    g0622(.A(new_n803), .ZN(new_n823));
  INV_X1    g0623(.A(G326), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n823), .A2(new_n824), .B1(new_n816), .B2(new_n587), .ZN(new_n825));
  XNOR2_X1  g0625(.A(KEYINPUT33), .B(G317), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(new_n802), .B2(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n819), .A2(G329), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n798), .A2(G283), .ZN(new_n829));
  INV_X1    g0629(.A(G322), .ZN(new_n830));
  INV_X1    g0630(.A(G311), .ZN(new_n831));
  OAI22_X1  g0631(.A1(new_n805), .A2(new_n830), .B1(new_n811), .B2(new_n831), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n296), .B(new_n832), .C1(G303), .C2(new_n809), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n827), .A2(new_n828), .A3(new_n829), .A4(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n792), .B1(new_n822), .B2(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n771), .ZN(new_n836));
  NOR4_X1   g0636(.A1(new_n779), .A2(new_n791), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n774), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(G396));
  NAND2_X1  g0639(.A1(new_n417), .A2(KEYINPUT105), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT105), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n407), .A2(new_n841), .A3(new_n416), .A4(new_n413), .ZN(new_n842));
  AND3_X1   g0642(.A1(new_n422), .A2(new_n840), .A3(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n705), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AND3_X1   g0645(.A1(new_n684), .A2(new_n687), .A3(new_n685), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n659), .B1(new_n692), .B2(new_n693), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n678), .A2(new_n657), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n848), .A2(new_n672), .A3(new_n602), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n657), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n845), .B1(new_n846), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n407), .A2(new_n716), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n422), .A2(new_n840), .A3(new_n852), .A4(new_n842), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n652), .A2(new_n716), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n851), .B1(new_n738), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n771), .B1(new_n856), .B2(new_n763), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n763), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n792), .A2(new_n776), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n771), .B1(G77), .B2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n817), .A2(G97), .B1(G294), .B2(new_n806), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n861), .B(KEYINPUT103), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n338), .B1(new_n811), .B2(new_n612), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n863), .B1(G107), .B2(new_n809), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n802), .A2(G283), .B1(new_n803), .B2(G303), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n797), .A2(new_n498), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n866), .B1(G311), .B2(new_n819), .ZN(new_n867));
  NAND4_X1  g0667(.A1(new_n862), .A2(new_n864), .A3(new_n865), .A4(new_n867), .ZN(new_n868));
  AOI22_X1  g0668(.A1(new_n806), .A2(G143), .B1(new_n812), .B2(G159), .ZN(new_n869));
  INV_X1    g0669(.A(new_n802), .ZN(new_n870));
  INV_X1    g0670(.A(G150), .ZN(new_n871));
  INV_X1    g0671(.A(G137), .ZN(new_n872));
  OAI221_X1 g0672(.A(new_n869), .B1(new_n870), .B2(new_n871), .C1(new_n872), .C2(new_n823), .ZN(new_n873));
  XOR2_X1   g0673(.A(new_n873), .B(KEYINPUT34), .Z(new_n874));
  NOR2_X1   g0674(.A1(new_n797), .A2(new_n353), .ZN(new_n875));
  OAI22_X1  g0675(.A1(new_n808), .A2(new_n202), .B1(new_n816), .B2(new_n245), .ZN(new_n876));
  INV_X1    g0676(.A(G132), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n296), .B1(new_n818), .B2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n875), .B(new_n876), .C1(KEYINPUT104), .C2(new_n878), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(KEYINPUT104), .B2(new_n878), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n868), .B1(new_n874), .B2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n860), .B1(new_n881), .B2(new_n783), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n776), .B2(new_n855), .ZN(new_n883));
  AND2_X1   g0683(.A1(new_n858), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(G384));
  NOR2_X1   g0685(.A1(new_n768), .A2(new_n272), .ZN(new_n886));
  INV_X1    g0686(.A(G330), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n440), .A2(new_n705), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n888), .B1(new_n461), .B2(new_n440), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n472), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n470), .B1(new_n458), .B2(new_n463), .ZN(new_n891));
  INV_X1    g0691(.A(new_n888), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  AND4_X1   g0693(.A1(new_n639), .A2(new_n643), .A3(new_n645), .A4(new_n647), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n712), .A3(new_n705), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n895), .A2(new_n563), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n760), .A2(new_n761), .ZN(new_n897));
  OAI211_X1 g0697(.A(new_n893), .B(new_n855), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT108), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n762), .A2(KEYINPUT108), .A3(new_n855), .A4(new_n893), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT40), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT38), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n702), .B1(new_n360), .B2(new_n366), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n904), .B1(new_n371), .B2(new_n391), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n367), .A2(new_n383), .A3(new_n904), .ZN(new_n906));
  INV_X1    g0706(.A(KEYINPUT37), .ZN(new_n907));
  XNOR2_X1  g0707(.A(new_n906), .B(new_n907), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n903), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n907), .B1(new_n904), .B2(KEYINPUT107), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(new_n906), .ZN(new_n911));
  INV_X1    g0711(.A(new_n702), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n912), .B1(new_n374), .B2(new_n375), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n368), .A2(new_n370), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n913), .B1(new_n654), .B2(new_n914), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n911), .A2(new_n915), .A3(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n902), .B1(new_n909), .B2(new_n916), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n900), .A2(new_n901), .A3(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n367), .A2(new_n383), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n919), .A2(new_n910), .A3(new_n904), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT107), .ZN(new_n921));
  OAI21_X1  g0721(.A(KEYINPUT37), .B1(new_n913), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n906), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR3_X1   g0724(.A1(new_n905), .A2(new_n924), .A3(new_n903), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT38), .B1(new_n911), .B2(new_n915), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n902), .B1(new_n927), .B2(new_n898), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n918), .A2(new_n928), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n474), .A2(new_n762), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n887), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  XNOR2_X1  g0732(.A(new_n932), .B(KEYINPUT109), .ZN(new_n933));
  INV_X1    g0733(.A(new_n893), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n840), .A2(new_n842), .ZN(new_n935));
  NOR2_X1   g0735(.A1(new_n935), .A2(new_n716), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n934), .B1(new_n851), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n925), .B2(new_n926), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n914), .A2(new_n912), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n909), .A2(new_n916), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n470), .A2(new_n471), .A3(new_n705), .ZN(new_n944));
  INV_X1    g0744(.A(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n926), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(KEYINPUT39), .A3(new_n916), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n943), .A2(new_n945), .A3(new_n947), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n939), .A2(new_n940), .A3(new_n948), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n737), .B(new_n474), .C1(new_n738), .C2(new_n740), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n656), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n949), .B(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n886), .B1(new_n933), .B2(new_n952), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n953), .B1(new_n933), .B2(new_n952), .ZN(new_n954));
  INV_X1    g0754(.A(new_n528), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(KEYINPUT35), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(KEYINPUT35), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n956), .A2(G116), .A3(new_n227), .A4(new_n957), .ZN(new_n958));
  XOR2_X1   g0758(.A(KEYINPUT106), .B(KEYINPUT36), .Z(new_n959));
  XNOR2_X1  g0759(.A(new_n958), .B(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(G77), .B1(new_n245), .B2(new_n353), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n726), .A2(new_n961), .B1(G50), .B2(new_n353), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n962), .A2(new_n694), .A3(new_n378), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n954), .A2(new_n960), .A3(new_n963), .ZN(G367));
  NAND2_X1  g0764(.A1(new_n242), .A2(new_n787), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n785), .B1(new_n720), .B2(new_n405), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n836), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OR3_X1    g0767(.A1(new_n676), .A2(new_n677), .A3(new_n705), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n848), .A2(new_n968), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(new_n657), .B2(new_n968), .ZN(new_n970));
  OAI22_X1  g0770(.A1(new_n805), .A2(new_n871), .B1(new_n811), .B2(new_n202), .ZN(new_n971));
  AOI211_X1 g0771(.A(new_n338), .B(new_n971), .C1(G58), .C2(new_n809), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n817), .A2(G68), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n802), .A2(G159), .B1(new_n803), .B2(G143), .ZN(new_n974));
  AOI22_X1  g0774(.A1(G77), .A2(new_n798), .B1(new_n819), .B2(G137), .ZN(new_n975));
  NAND4_X1  g0775(.A1(new_n972), .A2(new_n973), .A3(new_n974), .A4(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(G283), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n338), .B1(new_n811), .B2(new_n977), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n823), .A2(new_n831), .B1(new_n816), .B2(new_n206), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(G303), .C2(new_n806), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n797), .A2(new_n205), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G317), .B2(new_n819), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n809), .A2(KEYINPUT46), .A3(G116), .ZN(new_n983));
  INV_X1    g0783(.A(KEYINPUT46), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n984), .B1(new_n808), .B2(new_n612), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n983), .B(new_n985), .C1(new_n870), .C2(new_n587), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n980), .B(new_n982), .C1(KEYINPUT111), .C2(new_n986), .ZN(new_n987));
  AND2_X1   g0787(.A1(new_n986), .A2(KEYINPUT111), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n976), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT47), .Z(new_n990));
  OAI221_X1 g0790(.A(new_n967), .B1(new_n778), .B2(new_n970), .C1(new_n990), .C2(new_n792), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n672), .B1(new_n532), .B2(new_n705), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n668), .A2(new_n716), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n718), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n995), .A2(KEYINPUT110), .ZN(new_n999));
  OR3_X1    g0799(.A1(new_n997), .A2(new_n998), .A3(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n998), .B1(new_n997), .B2(new_n999), .ZN(new_n1001));
  NOR2_X1   g0801(.A1(new_n718), .A2(new_n994), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT44), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1000), .A2(new_n1001), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n715), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n717), .A2(new_n712), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n714), .B2(new_n717), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1010), .B(new_n709), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n765), .B1(new_n1008), .B2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g0812(.A(new_n721), .B(KEYINPUT41), .Z(new_n1013));
  INV_X1    g0813(.A(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n770), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n994), .A2(new_n712), .A3(new_n717), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1016), .A2(KEYINPUT42), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n560), .B1(new_n992), .B2(new_n660), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n1016), .A2(KEYINPUT42), .B1(new_n705), .B2(new_n1018), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n1017), .A2(new_n1019), .B1(KEYINPUT43), .B2(new_n970), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1020), .B(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1005), .A2(new_n994), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n1022), .B(new_n1023), .Z(new_n1024));
  OAI21_X1  g0824(.A(new_n991), .B1(new_n1015), .B2(new_n1024), .ZN(G387));
  NOR2_X1   g0825(.A1(new_n764), .A2(new_n1011), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n764), .A2(new_n1011), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n1027), .A2(new_n721), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1011), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n714), .A2(new_n778), .ZN(new_n1031));
  INV_X1    g0831(.A(new_n789), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1032), .A2(new_n724), .B1(G107), .B2(new_n229), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n239), .A2(G45), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n724), .ZN(new_n1035));
  AOI211_X1 g0835(.A(G45), .B(new_n1035), .C1(G68), .C2(G77), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n401), .A2(G50), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT50), .ZN(new_n1038));
  AOI211_X1 g0838(.A(new_n720), .B(new_n296), .C1(new_n1036), .C2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1033), .B1(new_n1034), .B2(new_n1039), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n771), .B1(new_n1040), .B2(new_n785), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n808), .A2(new_n587), .B1(new_n816), .B2(new_n977), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n806), .A2(G317), .B1(new_n812), .B2(G303), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n870), .B2(new_n831), .C1(new_n830), .C2(new_n823), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  AND2_X1   g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI221_X1 g0850(.A(new_n338), .B1(new_n818), .B2(new_n824), .C1(new_n612), .C2(new_n797), .ZN(new_n1051));
  OR3_X1    g0851(.A1(new_n1049), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n296), .B1(new_n805), .B2(new_n202), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n809), .A2(G77), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(new_n353), .B2(new_n811), .ZN(new_n1055));
  AOI211_X1 g0855(.A(new_n1053), .B(new_n1055), .C1(G159), .C2(new_n803), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n818), .A2(new_n871), .ZN(new_n1057));
  AOI211_X1 g0857(.A(new_n981), .B(new_n1057), .C1(new_n263), .C2(new_n802), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n817), .A2(new_n405), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1056), .A2(new_n1058), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1052), .A2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1041), .B1(new_n1061), .B2(new_n783), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1030), .A2(new_n770), .B1(new_n1031), .B2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1029), .A2(new_n1063), .ZN(G393));
  INV_X1    g0864(.A(new_n1008), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n722), .B1(new_n1065), .B2(new_n1026), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1008), .A2(new_n1027), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1065), .A2(new_n770), .ZN(new_n1069));
  AND2_X1   g0869(.A1(new_n251), .A2(new_n787), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n784), .B1(new_n205), .B2(new_n229), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n771), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n338), .B1(new_n811), .B2(new_n587), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n870), .A2(new_n625), .B1(new_n816), .B2(new_n612), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1073), .B(new_n1074), .C1(G283), .C2(new_n809), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1075), .B(new_n799), .C1(new_n830), .C2(new_n818), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G317), .A2(new_n803), .B1(new_n806), .B2(G311), .ZN(new_n1077));
  XNOR2_X1  g0877(.A(new_n1077), .B(KEYINPUT52), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n1079), .A2(KEYINPUT112), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1079), .A2(KEYINPUT112), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n338), .B1(new_n809), .B2(G68), .ZN(new_n1082));
  OAI221_X1 g0882(.A(new_n1082), .B1(new_n401), .B2(new_n811), .C1(new_n870), .C2(new_n202), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n866), .B(new_n1083), .C1(G143), .C2(new_n819), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n806), .A2(G159), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n823), .B2(new_n871), .ZN(new_n1086));
  INV_X1    g0886(.A(KEYINPUT51), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n1086), .A2(new_n1087), .B1(G77), .B2(new_n817), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1084), .B(new_n1088), .C1(new_n1087), .C2(new_n1086), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1080), .A2(new_n1081), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1072), .B1(new_n1090), .B2(new_n783), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1091), .B1(new_n994), .B2(new_n778), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1068), .A2(new_n1069), .A3(new_n1092), .ZN(G390));
  OAI21_X1  g0893(.A(new_n771), .B1(new_n263), .B2(new_n859), .ZN(new_n1094));
  OAI22_X1  g0894(.A1(new_n805), .A2(new_n612), .B1(new_n811), .B2(new_n205), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n296), .B(new_n1095), .C1(G87), .C2(new_n809), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n817), .A2(G77), .ZN(new_n1097));
  AOI22_X1  g0897(.A1(new_n802), .A2(G107), .B1(new_n803), .B2(G283), .ZN(new_n1098));
  AOI21_X1  g0898(.A(new_n875), .B1(G294), .B2(new_n819), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1096), .A2(new_n1097), .A3(new_n1098), .A4(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n808), .A2(new_n871), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(new_n1101), .B(KEYINPUT53), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n819), .A2(G125), .ZN(new_n1103));
  OAI211_X1 g0903(.A(new_n1102), .B(new_n1103), .C1(new_n202), .C2(new_n797), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n817), .A2(G159), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n802), .A2(G137), .B1(new_n803), .B2(G128), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n812), .A2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n338), .B1(new_n806), .B2(G132), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  OAI21_X1  g0911(.A(new_n1100), .B1(new_n1104), .B2(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1094), .B1(new_n1112), .B2(new_n783), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n943), .A2(new_n947), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1113), .B1(new_n1115), .B2(new_n776), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n855), .ZN(new_n1117));
  NOR3_X1   g0917(.A1(new_n763), .A2(new_n934), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n844), .B1(new_n680), .B2(new_n688), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n893), .B1(new_n1119), .B2(new_n936), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1120), .A2(new_n944), .B1(new_n943), .B2(new_n947), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n944), .B(KEYINPUT113), .Z(new_n1122));
  NAND2_X1  g0922(.A1(new_n941), .A2(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n716), .B1(new_n730), .B2(new_n735), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n843), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1125), .A2(new_n937), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1123), .B1(new_n1126), .B2(new_n893), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1118), .B1(new_n1121), .B2(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n1114), .B1(new_n938), .B2(new_n945), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n897), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n887), .B1(new_n1130), .B2(new_n747), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1131), .A2(new_n855), .A3(new_n893), .ZN(new_n1132));
  AOI21_X1  g0932(.A(new_n936), .B1(new_n1124), .B2(new_n843), .ZN(new_n1133));
  OAI211_X1 g0933(.A(new_n941), .B(new_n1122), .C1(new_n1133), .C2(new_n934), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1129), .A2(new_n1132), .A3(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(new_n770), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1116), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n474), .A2(new_n1131), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n950), .A2(new_n656), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT114), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n893), .B1(new_n1131), .B2(new_n855), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n1118), .A2(new_n1142), .B1(new_n1119), .B2(new_n936), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n934), .B1(new_n763), .B2(new_n1117), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1144), .A2(new_n1133), .A3(new_n1132), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT114), .ZN(new_n1147));
  NAND4_X1  g0947(.A1(new_n950), .A2(new_n1147), .A3(new_n656), .A4(new_n1139), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1141), .A2(new_n1146), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1149), .A2(KEYINPUT115), .ZN(new_n1150));
  AND2_X1   g0950(.A1(new_n1128), .A2(new_n1135), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n722), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1136), .A2(KEYINPUT115), .A3(new_n1149), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1138), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(G378));
  NAND3_X1  g0955(.A1(new_n1128), .A2(new_n1135), .A3(new_n1146), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1141), .A2(new_n1148), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1157), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1156), .A2(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n918), .A2(new_n928), .A3(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT120), .ZN(new_n1161));
  NAND2_X1  g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n918), .A2(new_n928), .A3(KEYINPUT120), .A4(G330), .ZN(new_n1163));
  XOR2_X1   g0963(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n651), .A2(new_n313), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n324), .A2(new_n1164), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n281), .A2(new_n912), .ZN(new_n1169));
  XNOR2_X1  g0969(.A(new_n1169), .B(KEYINPUT119), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1168), .A2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1166), .A2(new_n1170), .A3(new_n1167), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1162), .A2(new_n1163), .A3(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(new_n1160), .ZN(new_n1176));
  INV_X1    g0976(.A(new_n1174), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1176), .A2(KEYINPUT120), .A3(new_n1177), .ZN(new_n1178));
  AND3_X1   g0978(.A1(new_n1175), .A2(new_n949), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n949), .B1(new_n1175), .B2(new_n1178), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1159), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT57), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n722), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n949), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1162), .A2(new_n1163), .A3(new_n1174), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1160), .A2(new_n1174), .A3(new_n1161), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1184), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT121), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1175), .A2(new_n949), .A3(new_n1178), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1179), .B1(new_n1180), .B2(KEYINPUT121), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1182), .B1(new_n1156), .B2(new_n1158), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n1190), .A2(new_n1191), .A3(new_n1192), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1183), .A2(new_n1193), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n770), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1177), .A2(new_n775), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n771), .B1(G50), .B2(new_n859), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1054), .A2(new_n283), .A3(new_n338), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n1198), .B(KEYINPUT116), .Z(new_n1199));
  NAND2_X1  g0999(.A1(new_n798), .A2(G58), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n1200), .B1(new_n977), .B2(new_n818), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n803), .A2(G116), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n802), .A2(G97), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n806), .A2(G107), .B1(new_n812), .B2(new_n405), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n973), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(new_n1199), .A2(new_n1201), .A3(new_n1205), .ZN(new_n1206));
  XOR2_X1   g1006(.A(new_n1206), .B(KEYINPUT58), .Z(new_n1207));
  AOI21_X1  g1007(.A(G50), .B1(new_n264), .B2(new_n283), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1208), .B1(new_n296), .B2(G41), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n817), .A2(G150), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n802), .A2(G132), .B1(new_n803), .B2(G125), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n812), .A2(G137), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n806), .B1(new_n809), .B2(new_n1108), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1212), .A4(new_n1213), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1214), .A2(KEYINPUT59), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(KEYINPUT117), .B(G124), .ZN(new_n1217));
  OAI211_X1 g1017(.A(new_n264), .B(new_n283), .C1(new_n818), .C2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1218), .B1(G159), .B2(new_n798), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1207), .B(new_n1209), .C1(new_n1215), .C2(new_n1220), .ZN(new_n1221));
  INV_X1    g1021(.A(KEYINPUT118), .ZN(new_n1222));
  OR2_X1    g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n792), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1197), .B1(new_n1223), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1196), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1195), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1194), .A2(new_n1228), .ZN(G375));
  INV_X1    g1029(.A(new_n1146), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1157), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1231), .A2(new_n1014), .A3(new_n1149), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n934), .A2(new_n775), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n771), .B1(G68), .B2(new_n859), .ZN(new_n1234));
  OAI22_X1  g1034(.A1(new_n205), .A2(new_n808), .B1(new_n811), .B2(new_n206), .ZN(new_n1235));
  AOI211_X1 g1035(.A(new_n296), .B(new_n1235), .C1(G283), .C2(new_n806), .ZN(new_n1236));
  AOI22_X1  g1036(.A1(new_n802), .A2(G116), .B1(new_n803), .B2(G294), .ZN(new_n1237));
  AOI22_X1  g1037(.A1(G77), .A2(new_n798), .B1(new_n819), .B2(G303), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1236), .A2(new_n1059), .A3(new_n1237), .A4(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n819), .A2(G128), .B1(new_n809), .B2(G159), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT122), .Z(new_n1241));
  OAI21_X1  g1041(.A(new_n296), .B1(new_n805), .B2(new_n872), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1242), .B1(G150), .B2(new_n812), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n817), .A2(G50), .ZN(new_n1244));
  AOI22_X1  g1044(.A1(G132), .A2(new_n803), .B1(new_n802), .B2(new_n1108), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1243), .A2(new_n1244), .A3(new_n1245), .A4(new_n1200), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1241), .B2(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1234), .B1(new_n1247), .B2(new_n783), .ZN(new_n1248));
  AOI22_X1  g1048(.A1(new_n1146), .A2(new_n770), .B1(new_n1233), .B2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1232), .A2(new_n1249), .ZN(G381));
  OR2_X1    g1050(.A1(new_n1015), .A2(new_n1024), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1069), .A2(new_n1092), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n991), .A3(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1254), .ZN(new_n1255));
  INV_X1    g1055(.A(G375), .ZN(new_n1256));
  NOR4_X1   g1056(.A1(G381), .A2(G396), .A3(G384), .A4(G393), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1255), .A2(new_n1256), .A3(new_n1154), .A4(new_n1257), .ZN(new_n1258));
  XOR2_X1   g1058(.A(new_n1258), .B(KEYINPUT123), .Z(G407));
  AND2_X1   g1059(.A1(new_n703), .A2(G213), .ZN(new_n1260));
  XOR2_X1   g1060(.A(new_n1260), .B(KEYINPUT124), .Z(new_n1261));
  NAND2_X1  g1061(.A1(new_n1154), .A2(new_n1261), .ZN(new_n1262));
  OAI211_X1 g1062(.A(G407), .B(G213), .C1(G375), .C2(new_n1262), .ZN(G409));
  NAND2_X1  g1063(.A1(G390), .A2(G387), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(G393), .A2(G396), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n838), .B1(new_n1029), .B2(new_n1063), .ZN(new_n1266));
  OAI21_X1  g1066(.A(KEYINPUT126), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1254), .A2(new_n1264), .A3(new_n1267), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1265), .A2(new_n1266), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT126), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1268), .A2(new_n1272), .ZN(new_n1273));
  NAND4_X1  g1073(.A1(new_n1254), .A2(new_n1271), .A3(new_n1264), .A4(new_n1267), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1194), .A2(G378), .A3(new_n1228), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1190), .A2(new_n1191), .A3(new_n770), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1277), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1226), .B1(new_n1181), .B2(new_n1013), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1154), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1260), .B1(new_n1276), .B2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1231), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1157), .A2(KEYINPUT60), .A3(new_n1230), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(new_n721), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n1249), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1286), .A2(new_n884), .ZN(new_n1287));
  NAND3_X1  g1087(.A1(new_n1285), .A2(G384), .A3(new_n1249), .ZN(new_n1288));
  AND2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(KEYINPUT62), .B1(new_n1281), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1261), .ZN(new_n1291));
  AOI211_X1 g1091(.A(new_n1154), .B(new_n1227), .C1(new_n1183), .C2(new_n1193), .ZN(new_n1292));
  AOI22_X1  g1092(.A1(new_n1187), .A2(new_n1189), .B1(new_n1158), .B2(new_n1156), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n1293), .A2(new_n1014), .B1(new_n1196), .B2(new_n1225), .ZN(new_n1294));
  AOI21_X1  g1094(.A(G378), .B1(new_n1294), .B2(new_n1277), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1291), .B1(new_n1292), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(KEYINPUT127), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT127), .ZN(new_n1298));
  OAI211_X1 g1098(.A(new_n1298), .B(new_n1291), .C1(new_n1292), .C2(new_n1295), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1289), .A2(KEYINPUT62), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1290), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  NAND4_X1  g1102(.A1(new_n1287), .A2(G2897), .A3(new_n1260), .A4(new_n1288), .ZN(new_n1303));
  AND2_X1   g1103(.A1(new_n1261), .A2(G2897), .ZN(new_n1304));
  OAI21_X1  g1104(.A(new_n1303), .B1(new_n1289), .B2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1297), .A2(new_n1299), .A3(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(KEYINPUT61), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1275), .B1(new_n1302), .B2(new_n1308), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT63), .B1(new_n1281), .B2(new_n1289), .ZN(new_n1310));
  NOR3_X1   g1110(.A1(new_n1275), .A2(new_n1310), .A3(KEYINPUT61), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1300), .A2(KEYINPUT63), .A3(new_n1289), .ZN(new_n1312));
  AND2_X1   g1112(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1281), .A2(KEYINPUT125), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1305), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1311), .A2(new_n1312), .A3(new_n1315), .ZN(new_n1316));
  NAND2_X1  g1116(.A1(new_n1309), .A2(new_n1316), .ZN(G405));
  NAND2_X1  g1117(.A1(G375), .A2(new_n1154), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n1276), .ZN(new_n1319));
  XNOR2_X1  g1119(.A(new_n1319), .B(new_n1289), .ZN(new_n1320));
  XNOR2_X1  g1120(.A(new_n1320), .B(new_n1275), .ZN(G402));
endmodule


