//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 1 0 0 0 0 1 0 0 1 0 1 0 1 0 0 1 0 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:38 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1125, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1279, new_n1280, new_n1281, new_n1282, new_n1283,
    new_n1284, new_n1285, new_n1286, new_n1287, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1298, new_n1299, new_n1300, new_n1301, new_n1302,
    new_n1303, new_n1304, new_n1305, new_n1307, new_n1308, new_n1309,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1361, new_n1362, new_n1363, new_n1364, new_n1365,
    new_n1366, new_n1367, new_n1368, new_n1369, new_n1370;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  INV_X1    g0005(.A(G244), .ZN(new_n206));
  INV_X1    g0006(.A(G107), .ZN(new_n207));
  INV_X1    g0007(.A(G264), .ZN(new_n208));
  OAI221_X1 g0008(.A(new_n204), .B1(new_n205), .B2(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n210));
  INV_X1    g0010(.A(G58), .ZN(new_n211));
  INV_X1    g0011(.A(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G97), .ZN(new_n213));
  INV_X1    g0013(.A(G257), .ZN(new_n214));
  OAI221_X1 g0014(.A(new_n210), .B1(new_n211), .B2(new_n212), .C1(new_n213), .C2(new_n214), .ZN(new_n215));
  OAI21_X1  g0015(.A(new_n203), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  OR2_X1    g0016(.A1(new_n216), .A2(KEYINPUT1), .ZN(new_n217));
  OAI21_X1  g0017(.A(G50), .B1(G58), .B2(G68), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT64), .ZN(new_n219));
  NAND2_X1  g0019(.A1(G1), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(G20), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n203), .A2(G13), .ZN(new_n224));
  OAI211_X1 g0024(.A(new_n224), .B(G250), .C1(G257), .C2(G264), .ZN(new_n225));
  XNOR2_X1  g0025(.A(new_n225), .B(KEYINPUT0), .ZN(new_n226));
  NAND3_X1  g0026(.A1(new_n217), .A2(new_n223), .A3(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n216), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(new_n212), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G68), .B(G77), .Z(new_n237));
  XOR2_X1   g0037(.A(G50), .B(G58), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  NAND2_X1  g0043(.A1(G33), .A2(G41), .ZN(new_n244));
  NAND3_X1  g0044(.A1(new_n244), .A2(G1), .A3(G13), .ZN(new_n245));
  INV_X1    g0045(.A(G1), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n246), .B1(G41), .B2(G45), .ZN(new_n247));
  AND3_X1   g0047(.A1(new_n245), .A2(KEYINPUT65), .A3(new_n247), .ZN(new_n248));
  AOI21_X1  g0048(.A(KEYINPUT65), .B1(new_n245), .B2(new_n247), .ZN(new_n249));
  OAI21_X1  g0049(.A(G226), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT3), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G33), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n205), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n220), .B1(G33), .B2(G41), .ZN(new_n257));
  MUX2_X1   g0057(.A(G222), .B(G223), .S(G1698), .Z(new_n258));
  OAI211_X1 g0058(.A(new_n256), .B(new_n257), .C1(new_n255), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n247), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(new_n245), .A3(G274), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n250), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  OR2_X1    g0062(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(KEYINPUT66), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G169), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND3_X1  g0068(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(new_n220), .ZN(new_n270));
  XNOR2_X1  g0070(.A(KEYINPUT8), .B(G58), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n221), .A2(G33), .ZN(new_n272));
  INV_X1    g0072(.A(G150), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n221), .A2(new_n253), .ZN(new_n274));
  OAI22_X1  g0074(.A1(new_n271), .A2(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G50), .A2(G58), .ZN(new_n276));
  INV_X1    g0076(.A(G68), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n221), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n270), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g0079(.A1(new_n246), .A2(G13), .A3(G20), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n281), .A2(new_n270), .ZN(new_n282));
  INV_X1    g0082(.A(G50), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n246), .B2(G20), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n282), .A2(new_n284), .B1(new_n283), .B2(new_n281), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n287), .B1(new_n265), .B2(new_n288), .ZN(new_n289));
  AND2_X1   g0089(.A1(new_n268), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g0092(.A1(KEYINPUT71), .A2(KEYINPUT9), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XOR2_X1   g0094(.A(new_n294), .B(KEYINPUT72), .Z(new_n295));
  INV_X1    g0095(.A(KEYINPUT10), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n266), .A2(G200), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n265), .A2(G190), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n295), .A2(new_n296), .A3(new_n297), .A4(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n297), .A2(new_n294), .A3(new_n298), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT10), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n290), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT18), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n211), .A2(new_n277), .ZN(new_n304));
  NOR2_X1   g0104(.A1(G58), .A2(G68), .ZN(new_n305));
  OAI21_X1  g0105(.A(G20), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(G20), .A2(G33), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n307), .A2(G159), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n253), .A2(KEYINPUT74), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT74), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n312), .A2(G33), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n311), .A2(new_n313), .A3(KEYINPUT3), .ZN(new_n314));
  AOI21_X1  g0114(.A(G20), .B1(new_n314), .B2(new_n252), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT7), .ZN(new_n316));
  OAI21_X1  g0116(.A(G68), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n252), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT74), .B(G33), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n320));
  NOR3_X1   g0120(.A1(new_n320), .A2(KEYINPUT7), .A3(G20), .ZN(new_n321));
  OAI211_X1 g0121(.A(KEYINPUT16), .B(new_n310), .C1(new_n317), .C2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT16), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n316), .A2(G20), .ZN(new_n324));
  AOI21_X1  g0124(.A(KEYINPUT3), .B1(new_n311), .B2(new_n313), .ZN(new_n325));
  INV_X1    g0125(.A(new_n254), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT3), .B(G33), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n316), .B1(new_n328), .B2(G20), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n277), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n323), .B1(new_n330), .B2(new_n309), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n322), .A2(new_n331), .A3(new_n270), .ZN(new_n332));
  INV_X1    g0132(.A(new_n271), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n246), .A2(G20), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n282), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n271), .A2(new_n281), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n337), .B(KEYINPUT75), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  MUX2_X1   g0139(.A(G223), .B(G226), .S(G1698), .Z(new_n340));
  NAND3_X1  g0140(.A1(new_n340), .A2(new_n314), .A3(new_n252), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G87), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n245), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n245), .A2(new_n247), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n261), .B1(new_n212), .B2(new_n344), .ZN(new_n345));
  NOR2_X1   g0145(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G179), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n347), .B1(new_n267), .B2(new_n346), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n303), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT17), .ZN(new_n351));
  XNOR2_X1  g0151(.A(KEYINPUT76), .B(G190), .ZN(new_n352));
  NOR4_X1   g0152(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT77), .A4(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G200), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n343), .B2(new_n345), .ZN(new_n355));
  INV_X1    g0155(.A(KEYINPUT77), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(new_n352), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n346), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n353), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n351), .B1(new_n339), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n357), .A2(new_n359), .ZN(new_n362));
  INV_X1    g0162(.A(new_n353), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n364), .A2(KEYINPUT17), .A3(new_n332), .A4(new_n338), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n339), .A2(new_n303), .A3(new_n348), .ZN(new_n366));
  NAND4_X1  g0166(.A1(new_n350), .A2(new_n361), .A3(new_n365), .A4(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n280), .A2(KEYINPUT68), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT68), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n370), .A2(new_n246), .A3(G13), .A4(G20), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n270), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(G68), .A3(new_n334), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n221), .A2(G33), .A3(G77), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n374), .B1(new_n221), .B2(G68), .C1(new_n274), .C2(new_n283), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT11), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n375), .A2(new_n376), .A3(new_n270), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n376), .B1(new_n375), .B2(new_n270), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n246), .A2(G13), .ZN(new_n380));
  NOR4_X1   g0180(.A1(new_n380), .A2(KEYINPUT12), .A3(new_n221), .A4(G68), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n369), .A2(new_n371), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n277), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n381), .B1(new_n384), .B2(KEYINPUT12), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(G33), .A2(G97), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g0189(.A1(G226), .A2(G1698), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n212), .B2(G1698), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n389), .B1(new_n391), .B2(new_n328), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n261), .B1(new_n392), .B2(new_n245), .ZN(new_n393));
  INV_X1    g0193(.A(G238), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT65), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n344), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n245), .A2(KEYINPUT65), .A3(new_n247), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(KEYINPUT13), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  OAI21_X1  g0199(.A(G238), .B1(new_n248), .B2(new_n249), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n212), .A2(G1698), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n401), .B1(G226), .B2(G1698), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n388), .B1(new_n402), .B2(new_n255), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n403), .A2(new_n257), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT13), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n400), .A2(new_n404), .A3(new_n405), .A4(new_n261), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n399), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT14), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(G169), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n399), .A2(G179), .A3(new_n406), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n408), .B1(new_n407), .B2(G169), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n387), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT69), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n414), .B1(new_n382), .B2(G77), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n369), .A2(KEYINPUT69), .A3(new_n205), .A4(new_n371), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n372), .A2(G77), .A3(new_n334), .ZN(new_n418));
  NAND2_X1  g0218(.A1(G20), .A2(G77), .ZN(new_n419));
  XNOR2_X1  g0219(.A(KEYINPUT15), .B(G87), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n419), .B1(new_n420), .B2(new_n272), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n271), .A2(new_n274), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n270), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n417), .A2(new_n418), .A3(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n394), .A2(G1698), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n426), .B1(G232), .B2(G1698), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n245), .B1(new_n427), .B2(new_n328), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n255), .A2(new_n207), .ZN(new_n429));
  INV_X1    g0229(.A(G274), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n257), .A2(new_n430), .ZN(new_n431));
  AOI22_X1  g0231(.A1(new_n428), .A2(new_n429), .B1(new_n431), .B2(new_n260), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT67), .ZN(new_n433));
  OAI21_X1  g0233(.A(G244), .B1(new_n248), .B2(new_n249), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n432), .A2(new_n433), .A3(G190), .A4(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n427), .A2(new_n328), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n429), .A3(new_n257), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n434), .A2(new_n261), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(KEYINPUT67), .B1(new_n438), .B2(G200), .ZN(new_n439));
  INV_X1    g0239(.A(G190), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n425), .B(new_n435), .C1(new_n439), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n438), .A2(new_n267), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n432), .A2(new_n288), .A3(new_n434), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n443), .A2(new_n424), .A3(new_n444), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT70), .ZN(new_n447));
  OR2_X1    g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n399), .A2(G190), .A3(new_n406), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n449), .A2(new_n386), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n354), .B1(new_n399), .B2(new_n406), .ZN(new_n451));
  OAI21_X1  g0251(.A(KEYINPUT73), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n407), .A2(G200), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT73), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n453), .A2(new_n454), .A3(new_n386), .A4(new_n449), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n446), .A2(new_n447), .ZN(new_n457));
  AND4_X1   g0257(.A1(new_n413), .A2(new_n448), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n302), .A2(new_n368), .A3(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT80), .ZN(new_n460));
  NOR2_X1   g0260(.A1(G238), .A2(G1698), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n461), .B1(new_n206), .B2(G1698), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n462), .A2(new_n314), .A3(new_n252), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n464), .B1(new_n311), .B2(new_n313), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n245), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(G45), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G1), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n430), .ZN(new_n470));
  INV_X1    g0270(.A(G250), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n471), .B1(new_n468), .B2(G1), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n470), .A2(new_n245), .A3(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n460), .B1(new_n467), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g0275(.A(new_n465), .B1(new_n320), .B2(new_n462), .ZN(new_n476));
  OAI211_X1 g0276(.A(KEYINPUT80), .B(new_n473), .C1(new_n476), .C2(new_n245), .ZN(new_n477));
  AOI21_X1  g0277(.A(G169), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n477), .A3(new_n288), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n246), .A2(G33), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n282), .A2(new_n480), .ZN(new_n481));
  INV_X1    g0281(.A(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(new_n420), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NOR2_X1   g0284(.A1(new_n382), .A2(new_n483), .ZN(new_n485));
  INV_X1    g0285(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n320), .A2(new_n221), .A3(G68), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT19), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n221), .B1(new_n388), .B2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(G87), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n490), .A2(new_n213), .A3(new_n207), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n221), .A2(G33), .A3(G97), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n489), .A2(new_n491), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  AND2_X1   g0293(.A1(new_n487), .A2(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(new_n270), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n484), .B(new_n486), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n479), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n475), .A2(new_n477), .A3(G190), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n495), .B1(new_n487), .B2(new_n493), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n481), .A2(new_n490), .ZN(new_n500));
  NOR3_X1   g0300(.A1(new_n499), .A2(new_n500), .A3(new_n485), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n354), .B1(new_n475), .B2(new_n477), .ZN(new_n503));
  OAI22_X1  g0303(.A1(new_n478), .A2(new_n497), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT81), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n463), .A2(new_n466), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n257), .ZN(new_n508));
  AOI21_X1  g0308(.A(KEYINPUT80), .B1(new_n508), .B2(new_n473), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n467), .A2(new_n460), .A3(new_n474), .ZN(new_n510));
  OAI21_X1  g0310(.A(new_n267), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n511), .A2(new_n479), .A3(new_n496), .ZN(new_n512));
  OAI21_X1  g0312(.A(G200), .B1(new_n509), .B2(new_n510), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(new_n498), .A3(new_n501), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT81), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n506), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(G257), .A2(G1698), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n517), .B1(new_n208), .B2(G1698), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n518), .A2(new_n314), .A3(new_n252), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n255), .A2(G303), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n245), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g0321(.A(KEYINPUT5), .B(G41), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(G274), .A3(new_n245), .A4(new_n469), .ZN(new_n523));
  AND2_X1   g0323(.A1(KEYINPUT5), .A2(G41), .ZN(new_n524));
  NOR2_X1   g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n469), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n245), .ZN(new_n527));
  INV_X1    g0327(.A(G270), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n523), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NOR3_X1   g0329(.A1(new_n521), .A2(new_n529), .A3(new_n288), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n464), .A2(G20), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n270), .A2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(KEYINPUT84), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n270), .A2(KEYINPUT84), .A3(new_n531), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(G33), .A2(G283), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n537), .B(new_n221), .C1(G33), .C2(new_n213), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT20), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  AOI221_X4 g0339(.A(new_n533), .B1(new_n464), .B2(G20), .C1(new_n269), .C2(new_n220), .ZN(new_n540));
  AOI21_X1  g0340(.A(KEYINPUT84), .B1(new_n270), .B2(new_n531), .ZN(new_n541));
  OAI211_X1 g0341(.A(KEYINPUT20), .B(new_n538), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n539), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g0344(.A(KEYINPUT83), .B1(new_n382), .B2(G116), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n369), .A2(new_n546), .A3(new_n464), .A4(new_n371), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n464), .B1(new_n246), .B2(G33), .ZN(new_n549));
  AND3_X1   g0349(.A1(new_n372), .A2(KEYINPUT82), .A3(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(KEYINPUT82), .B1(new_n372), .B2(new_n549), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n548), .B1(new_n550), .B2(new_n551), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n530), .B1(new_n544), .B2(new_n552), .ZN(new_n553));
  OAI21_X1  g0353(.A(G169), .B1(new_n521), .B2(new_n529), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n382), .A2(new_n495), .A3(new_n549), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT82), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n372), .A2(KEYINPUT82), .A3(new_n549), .ZN(new_n558));
  AOI22_X1  g0358(.A1(new_n557), .A2(new_n558), .B1(new_n545), .B2(new_n547), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n538), .B1(new_n540), .B2(new_n541), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n542), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n554), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n553), .B1(new_n564), .B2(KEYINPUT21), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT21), .ZN(new_n566));
  AOI211_X1 g0366(.A(new_n566), .B(new_n554), .C1(new_n563), .C2(new_n559), .ZN(new_n567));
  NOR2_X1   g0367(.A1(new_n521), .A2(new_n529), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n352), .ZN(new_n569));
  OAI21_X1  g0369(.A(G200), .B1(new_n521), .B2(new_n529), .ZN(new_n570));
  AND4_X1   g0370(.A1(new_n563), .A2(new_n569), .A3(new_n559), .A4(new_n570), .ZN(new_n571));
  NOR3_X1   g0371(.A1(new_n565), .A2(new_n567), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G250), .A2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n214), .B2(G1698), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n574), .A2(new_n314), .A3(new_n252), .ZN(new_n575));
  INV_X1    g0375(.A(G294), .ZN(new_n576));
  OR2_X1    g0376(.A1(new_n319), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n245), .B1(new_n575), .B2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n523), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n527), .A2(new_n208), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n582), .A2(G169), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(G179), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT22), .ZN(new_n586));
  NOR3_X1   g0386(.A1(new_n586), .A2(new_n490), .A3(G20), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n314), .A2(new_n587), .A3(new_n252), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n252), .A2(new_n254), .A3(new_n221), .A4(G87), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n586), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n465), .A2(new_n221), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT23), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n592), .B1(new_n221), .B2(G107), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n207), .A2(KEYINPUT23), .A3(G20), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(KEYINPUT85), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n589), .A2(new_n586), .B1(new_n593), .B2(new_n594), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT85), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n598), .A2(new_n599), .A3(new_n588), .A4(new_n591), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n597), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(KEYINPUT24), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n597), .A2(new_n603), .A3(new_n600), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n495), .B1(new_n602), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n281), .A2(new_n207), .ZN(new_n606));
  XNOR2_X1  g0406(.A(new_n606), .B(KEYINPUT25), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n481), .A2(new_n207), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n585), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  INV_X1    g0411(.A(KEYINPUT79), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n523), .B1(new_n527), .B2(new_n214), .ZN(new_n613));
  INV_X1    g0413(.A(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n206), .A2(G1698), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n537), .B1(new_n616), .B2(new_n255), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT4), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n314), .A2(new_n252), .A3(new_n615), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(new_n612), .B(new_n614), .C1(new_n620), .C2(new_n245), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n618), .ZN(new_n622));
  INV_X1    g0422(.A(G1698), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(G244), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n624), .A2(new_n618), .B1(new_n471), .B2(new_n623), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n625), .A2(new_n328), .B1(G33), .B2(G283), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n245), .B1(new_n622), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT79), .B1(new_n627), .B2(new_n613), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n621), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(new_n267), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n627), .A2(new_n613), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n207), .B1(new_n327), .B2(new_n329), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n307), .A2(G77), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT78), .ZN(new_n634));
  INV_X1    g0434(.A(KEYINPUT6), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n635), .A2(new_n213), .A3(G107), .ZN(new_n636));
  XNOR2_X1  g0436(.A(G97), .B(G107), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n636), .B1(new_n635), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n634), .B1(new_n221), .B2(new_n638), .ZN(new_n639));
  OAI21_X1  g0439(.A(new_n270), .B1(new_n632), .B2(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n280), .A2(G97), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n482), .B2(G97), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n288), .A2(new_n631), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  OAI21_X1  g0443(.A(G200), .B1(new_n627), .B2(new_n613), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n644), .A2(new_n640), .A3(new_n642), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n621), .A2(new_n628), .A3(G190), .ZN(new_n646));
  AOI22_X1  g0446(.A1(new_n630), .A2(new_n643), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n581), .A2(new_n354), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(G190), .B2(new_n581), .ZN(new_n649));
  INV_X1    g0449(.A(new_n604), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n603), .B1(new_n597), .B2(new_n600), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n270), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n649), .A2(new_n652), .A3(new_n609), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n572), .A2(new_n611), .A3(new_n647), .A4(new_n653), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n459), .A2(new_n516), .A3(new_n654), .ZN(G372));
  AND3_X1   g0455(.A1(new_n339), .A2(new_n303), .A3(new_n348), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n349), .ZN(new_n657));
  INV_X1    g0457(.A(new_n413), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n453), .A2(new_n386), .A3(new_n449), .ZN(new_n659));
  INV_X1    g0459(.A(new_n445), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n658), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n365), .A2(new_n361), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n657), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n299), .A2(new_n301), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n290), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OR2_X1    g0466(.A1(new_n565), .A2(new_n567), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n611), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n647), .A2(new_n653), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n508), .A2(new_n473), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(new_n267), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n479), .A2(new_n496), .A3(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n671), .A2(G200), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n498), .A2(new_n674), .A3(new_n501), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n670), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n669), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT86), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n673), .A2(new_n679), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n673), .A2(new_n679), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n630), .A2(new_n643), .A3(new_n673), .A4(new_n675), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n680), .B(new_n681), .C1(new_n682), .C2(KEYINPUT26), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n630), .A2(new_n643), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g0485(.A1(new_n506), .A2(new_n515), .A3(new_n685), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n683), .B1(new_n686), .B2(KEYINPUT26), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT87), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n678), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI211_X1 g0489(.A(KEYINPUT87), .B(new_n683), .C1(KEYINPUT26), .C2(new_n686), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n666), .B1(new_n691), .B2(new_n459), .ZN(G369));
  NAND2_X1  g0492(.A1(new_n559), .A2(new_n563), .ZN(new_n693));
  OR3_X1    g0493(.A1(new_n380), .A2(KEYINPUT27), .A3(G20), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT27), .B1(new_n380), .B2(G20), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G213), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(G343), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n667), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n693), .A2(new_n698), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n572), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(G330), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(new_n698), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT88), .B1(new_n611), .B2(new_n706), .ZN(new_n707));
  AOI22_X1  g0507(.A1(new_n652), .A2(new_n609), .B1(new_n583), .B2(new_n584), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT88), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n708), .A2(new_n709), .A3(new_n698), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n698), .B1(new_n605), .B2(new_n610), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n611), .A2(new_n712), .A3(new_n653), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n705), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n611), .A2(new_n698), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n667), .A2(new_n706), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n716), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n715), .A2(new_n719), .ZN(G399));
  INV_X1    g0520(.A(new_n224), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(G41), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n491), .A2(G116), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G1), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n219), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n725), .B1(new_n726), .B2(new_n723), .ZN(new_n727));
  XNOR2_X1  g0527(.A(new_n727), .B(KEYINPUT28), .ZN(new_n728));
  AND3_X1   g0528(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT81), .ZN(new_n729));
  AOI21_X1  g0529(.A(KEYINPUT81), .B1(new_n512), .B2(new_n514), .ZN(new_n730));
  NOR3_X1   g0530(.A1(new_n729), .A2(new_n730), .A3(new_n684), .ZN(new_n731));
  OAI21_X1  g0531(.A(KEYINPUT90), .B1(new_n731), .B2(KEYINPUT26), .ZN(new_n732));
  INV_X1    g0532(.A(KEYINPUT90), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT26), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n686), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n682), .A2(new_n734), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n732), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n667), .A2(new_n708), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n739), .A2(new_n670), .A3(new_n676), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n673), .B(new_n679), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n698), .B1(new_n738), .B2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(KEYINPUT29), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n706), .B1(new_n689), .B2(new_n690), .ZN(new_n745));
  INV_X1    g0545(.A(KEYINPUT29), .ZN(new_n746));
  AND3_X1   g0546(.A1(new_n745), .A2(KEYINPUT89), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(KEYINPUT89), .B1(new_n745), .B2(new_n746), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n744), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT30), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n578), .A2(new_n580), .ZN(new_n751));
  NAND4_X1  g0551(.A1(new_n530), .A2(new_n475), .A3(new_n477), .A4(new_n751), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n750), .B1(new_n629), .B2(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n631), .A2(new_n581), .ZN(new_n754));
  INV_X1    g0554(.A(new_n568), .ZN(new_n755));
  NAND4_X1  g0555(.A1(new_n754), .A2(new_n288), .A3(new_n671), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n629), .A2(new_n752), .A3(new_n750), .ZN(new_n758));
  OAI21_X1  g0558(.A(new_n698), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT31), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  OR3_X1    g0561(.A1(new_n629), .A2(new_n752), .A3(new_n750), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(new_n756), .A3(new_n753), .ZN(new_n763));
  AOI21_X1  g0563(.A(KEYINPUT31), .B1(new_n763), .B2(new_n698), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n670), .A2(new_n708), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n729), .A2(new_n730), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n766), .A2(new_n767), .A3(new_n572), .A4(new_n706), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(new_n704), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n749), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n728), .B1(new_n773), .B2(G1), .ZN(G364));
  INV_X1    g0574(.A(G13), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G20), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n246), .B1(new_n776), .B2(G45), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n722), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n702), .A2(G330), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n705), .B2(new_n781), .ZN(new_n782));
  NOR2_X1   g0582(.A1(G13), .A2(G33), .ZN(new_n783));
  INV_X1    g0583(.A(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(G20), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n703), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n267), .A2(KEYINPUT93), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n221), .B1(KEYINPUT93), .B2(new_n267), .ZN(new_n789));
  AOI21_X1  g0589(.A(new_n220), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n790), .A2(new_n785), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n239), .A2(G45), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n793), .B(KEYINPUT92), .Z(new_n794));
  NOR2_X1   g0594(.A1(new_n320), .A2(new_n721), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n794), .B(new_n795), .C1(G45), .C2(new_n726), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n721), .A2(new_n255), .ZN(new_n797));
  XNOR2_X1  g0597(.A(new_n797), .B(KEYINPUT91), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n798), .A2(G355), .B1(new_n464), .B2(new_n721), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n792), .B1(new_n796), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g0600(.A1(G20), .A2(G179), .ZN(new_n801));
  XNOR2_X1  g0601(.A(new_n801), .B(KEYINPUT94), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n802), .A2(G200), .A3(new_n352), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n804));
  INV_X1    g0604(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n803), .A2(KEYINPUT95), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n808), .A2(G326), .ZN(new_n809));
  NOR2_X1   g0609(.A1(new_n354), .A2(G179), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n810), .A2(G20), .A3(G190), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n255), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT99), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n221), .A2(G190), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n815), .A2(new_n810), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(G179), .A2(G200), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n815), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(new_n817), .A2(G283), .B1(new_n820), .B2(G329), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n221), .B1(new_n818), .B2(G190), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n821), .B1(new_n576), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n813), .A2(KEYINPUT99), .ZN(new_n824));
  NOR2_X1   g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  INV_X1    g0625(.A(G311), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n802), .A2(new_n440), .A3(new_n354), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n802), .A2(new_n354), .A3(new_n352), .ZN(new_n828));
  INV_X1    g0628(.A(G322), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n826), .A2(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n802), .A2(new_n440), .A3(G200), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  XNOR2_X1  g0632(.A(KEYINPUT33), .B(G317), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n830), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n809), .A2(new_n814), .A3(new_n825), .A4(new_n834), .ZN(new_n835));
  INV_X1    g0635(.A(new_n811), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(G87), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n837), .B(new_n328), .C1(new_n207), .C2(new_n816), .ZN(new_n838));
  XNOR2_X1  g0638(.A(new_n838), .B(KEYINPUT96), .ZN(new_n839));
  INV_X1    g0639(.A(new_n828), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(G58), .B2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n820), .A2(G159), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT32), .ZN(new_n843));
  INV_X1    g0643(.A(new_n827), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n843), .B1(G77), .B2(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n841), .B(new_n845), .C1(new_n283), .C2(new_n807), .ZN(new_n846));
  XNOR2_X1  g0646(.A(new_n822), .B(KEYINPUT97), .ZN(new_n847));
  AOI22_X1  g0647(.A1(new_n832), .A2(G68), .B1(new_n847), .B2(G97), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n848), .B(KEYINPUT98), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n835), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n800), .B1(new_n850), .B2(new_n790), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n786), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n782), .B1(new_n852), .B2(new_n780), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT100), .Z(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(G396));
  AND3_X1   g0655(.A1(new_n424), .A2(KEYINPUT101), .A3(new_n698), .ZN(new_n856));
  AOI21_X1  g0656(.A(KEYINPUT101), .B1(new_n424), .B2(new_n698), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n660), .B1(new_n858), .B2(new_n442), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n445), .A2(new_n698), .ZN(new_n860));
  OAI21_X1  g0660(.A(KEYINPUT102), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n424), .A2(new_n698), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT101), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n424), .A2(KEYINPUT101), .A3(new_n698), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n442), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n866), .A2(new_n445), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT102), .ZN(new_n868));
  INV_X1    g0668(.A(new_n860), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n861), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n871), .A2(new_n706), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n873), .B1(new_n689), .B2(new_n690), .ZN(new_n874));
  INV_X1    g0674(.A(new_n745), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n871), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n779), .B1(new_n876), .B2(new_n772), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n877), .B1(new_n772), .B2(new_n876), .ZN(new_n878));
  INV_X1    g0678(.A(new_n790), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n832), .A2(G150), .B1(new_n840), .B2(G143), .ZN(new_n880));
  INV_X1    g0680(.A(G159), .ZN(new_n881));
  INV_X1    g0681(.A(G137), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n880), .B1(new_n881), .B2(new_n827), .C1(new_n807), .C2(new_n882), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT34), .ZN(new_n884));
  INV_X1    g0684(.A(G132), .ZN(new_n885));
  OAI22_X1  g0685(.A1(new_n811), .A2(new_n283), .B1(new_n819), .B2(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n320), .B1(new_n211), .B2(new_n822), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n886), .B(new_n887), .C1(G68), .C2(new_n817), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n328), .B1(new_n836), .B2(G107), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n817), .A2(G87), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n890), .B(new_n891), .C1(new_n826), .C2(new_n819), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n892), .B1(G97), .B2(new_n847), .ZN(new_n893));
  OAI22_X1  g0693(.A1(new_n464), .A2(new_n827), .B1(new_n828), .B2(new_n576), .ZN(new_n894));
  AOI21_X1  g0694(.A(new_n894), .B1(G283), .B2(new_n832), .ZN(new_n895));
  OAI211_X1 g0695(.A(new_n893), .B(new_n895), .C1(new_n812), .C2(new_n807), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n879), .B1(new_n889), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n790), .A2(new_n783), .ZN(new_n898));
  AOI211_X1 g0698(.A(new_n780), .B(new_n897), .C1(new_n205), .C2(new_n898), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n784), .B2(new_n871), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n878), .A2(new_n900), .ZN(G384));
  INV_X1    g0701(.A(new_n638), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(KEYINPUT35), .ZN(new_n904));
  NAND4_X1  g0704(.A1(new_n903), .A2(G116), .A3(new_n222), .A4(new_n904), .ZN(new_n905));
  XNOR2_X1  g0705(.A(new_n905), .B(KEYINPUT36), .ZN(new_n906));
  NOR3_X1   g0706(.A1(new_n726), .A2(new_n205), .A3(new_n304), .ZN(new_n907));
  OAI22_X1  g0707(.A1(new_n907), .A2(KEYINPUT103), .B1(G50), .B2(new_n277), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(KEYINPUT103), .B2(new_n907), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n775), .A2(G1), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n906), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  XNOR2_X1  g0711(.A(new_n911), .B(KEYINPUT104), .ZN(new_n912));
  AOI21_X1  g0712(.A(new_n459), .B1(new_n743), .B2(KEYINPUT29), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n747), .B2(new_n748), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(new_n666), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n322), .A2(new_n270), .ZN(new_n917));
  OAI21_X1  g0717(.A(KEYINPUT7), .B1(new_n320), .B2(G20), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n315), .A2(new_n316), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n918), .A2(new_n919), .A3(G68), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT16), .B1(new_n920), .B2(new_n310), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n338), .B1(new_n917), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(new_n348), .ZN(new_n923));
  INV_X1    g0723(.A(new_n696), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n355), .A2(new_n356), .B1(new_n346), .B2(new_n358), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n332), .B(new_n338), .C1(new_n926), .C2(new_n353), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n925), .A3(new_n927), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n928), .A2(KEYINPUT37), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT105), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n339), .A2(new_n348), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n339), .A2(new_n924), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT37), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n931), .A2(new_n932), .A3(new_n933), .A4(new_n927), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n929), .A2(new_n930), .A3(new_n934), .ZN(new_n935));
  INV_X1    g0735(.A(new_n925), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n367), .A2(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n935), .A2(new_n937), .ZN(new_n938));
  AOI21_X1  g0738(.A(new_n930), .B1(new_n929), .B2(new_n934), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n916), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  AND2_X1   g0740(.A1(new_n332), .A2(new_n338), .ZN(new_n941));
  AOI22_X1  g0741(.A1(new_n941), .A2(new_n364), .B1(new_n922), .B2(new_n924), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n933), .B1(new_n942), .B2(new_n923), .ZN(new_n943));
  INV_X1    g0743(.A(new_n934), .ZN(new_n944));
  OAI21_X1  g0744(.A(KEYINPUT105), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n945), .A2(KEYINPUT38), .A3(new_n937), .A4(new_n935), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n387), .A2(new_n698), .ZN(new_n948));
  AND3_X1   g0748(.A1(new_n413), .A2(new_n659), .A3(new_n948), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n411), .A2(new_n412), .ZN(new_n950));
  AOI21_X1  g0750(.A(new_n948), .B1(new_n456), .B2(new_n950), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  INV_X1    g0752(.A(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(new_n683), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n731), .B2(new_n734), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n740), .B1(new_n955), .B2(KEYINPUT87), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n687), .A2(new_n688), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n872), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  OAI211_X1 g0758(.A(new_n947), .B(new_n953), .C1(new_n958), .C2(new_n860), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n696), .B1(new_n656), .B2(new_n349), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n931), .A2(new_n932), .A3(new_n927), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(new_n933), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n932), .B1(new_n662), .B2(new_n657), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n916), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n946), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(KEYINPUT39), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n940), .A2(KEYINPUT39), .A3(new_n946), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n658), .A2(new_n706), .ZN(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n967), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n959), .A2(new_n960), .A3(new_n971), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n915), .B(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n456), .A2(new_n950), .ZN(new_n974));
  INV_X1    g0774(.A(new_n948), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n413), .A2(new_n659), .A3(new_n948), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n976), .A2(new_n977), .B1(new_n870), .B2(new_n861), .ZN(new_n978));
  NOR3_X1   g0778(.A1(new_n654), .A2(new_n516), .A3(new_n698), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n759), .A2(new_n760), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n763), .A2(KEYINPUT31), .A3(new_n698), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n978), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(new_n940), .B2(new_n946), .ZN(new_n984));
  OR2_X1    g0784(.A1(new_n984), .A2(KEYINPUT40), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n868), .B1(new_n867), .B2(new_n869), .ZN(new_n986));
  AOI211_X1 g0786(.A(KEYINPUT102), .B(new_n860), .C1(new_n866), .C2(new_n445), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n949), .A2(new_n951), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(new_n988), .B1(new_n765), .B2(new_n768), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n965), .A2(KEYINPUT40), .A3(new_n989), .ZN(new_n990));
  AND2_X1   g0790(.A1(new_n985), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n459), .A2(new_n770), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n704), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(new_n992), .B2(new_n991), .ZN(new_n994));
  AND2_X1   g0794(.A1(new_n973), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(KEYINPUT106), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n246), .B2(new_n776), .C1(new_n973), .C2(new_n994), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n995), .A2(KEYINPUT106), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n912), .B1(new_n997), .B2(new_n998), .ZN(G367));
  INV_X1    g0799(.A(new_n795), .ZN(new_n1000));
  OAI221_X1 g0800(.A(new_n791), .B1(new_n224), .B2(new_n420), .C1(new_n1000), .C2(new_n235), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n255), .B1(new_n820), .B2(G137), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n211), .B2(new_n811), .C1(new_n205), .C2(new_n816), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n847), .A2(G68), .ZN(new_n1004));
  OAI221_X1 g0804(.A(new_n1004), .B1(new_n283), .B2(new_n827), .C1(new_n881), .C2(new_n831), .ZN(new_n1005));
  AOI211_X1 g0805(.A(new_n1003), .B(new_n1005), .C1(G150), .C2(new_n840), .ZN(new_n1006));
  INV_X1    g0806(.A(G143), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n807), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G283), .A2(new_n844), .B1(new_n832), .B2(G294), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n1009), .B1(new_n812), .B2(new_n828), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n320), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n817), .A2(G97), .ZN(new_n1012));
  INV_X1    g0812(.A(G317), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1011), .B(new_n1012), .C1(new_n1013), .C2(new_n819), .ZN(new_n1014));
  AOI21_X1  g0814(.A(KEYINPUT46), .B1(new_n836), .B2(G116), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n836), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n207), .B2(new_n822), .ZN(new_n1017));
  NOR4_X1   g0817(.A1(new_n1010), .A2(new_n1014), .A3(new_n1015), .A4(new_n1017), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n826), .B2(new_n807), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1008), .A2(new_n1019), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT47), .Z(new_n1021));
  OAI211_X1 g0821(.A(new_n779), .B(new_n1001), .C1(new_n1021), .C2(new_n879), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n501), .A2(new_n706), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n676), .A2(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1024), .B1(new_n741), .B2(new_n1023), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1022), .B1(new_n785), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n714), .B(new_n718), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(new_n705), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n645), .A2(new_n646), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n684), .A2(new_n1030), .ZN(new_n1031));
  AOI21_X1  g0831(.A(new_n706), .B1(new_n640), .B2(new_n642), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1031), .A2(new_n1032), .B1(new_n684), .B2(new_n706), .ZN(new_n1033));
  INV_X1    g0833(.A(KEYINPUT108), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT44), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1033), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n717), .B1(new_n711), .B2(new_n713), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1036), .B1(new_n1037), .B2(new_n716), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1036), .B1(new_n1034), .B2(new_n1035), .C1(new_n1037), .C2(new_n716), .ZN(new_n1041));
  AOI21_X1  g0841(.A(KEYINPUT45), .B1(new_n719), .B2(new_n1033), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1033), .ZN(new_n1043));
  INV_X1    g0843(.A(KEYINPUT45), .ZN(new_n1044));
  NOR4_X1   g0844(.A1(new_n1037), .A2(new_n1043), .A3(new_n1044), .A4(new_n716), .ZN(new_n1045));
  OAI211_X1 g0845(.A(new_n1040), .B(new_n1041), .C1(new_n1042), .C2(new_n1045), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1046), .A2(KEYINPUT109), .A3(new_n715), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n715), .B1(new_n1046), .B2(KEYINPUT109), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n1029), .B1(new_n1047), .B2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1049), .A2(new_n773), .ZN(new_n1050));
  XOR2_X1   g0850(.A(new_n722), .B(KEYINPUT41), .Z(new_n1051));
  INV_X1    g0851(.A(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n778), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n708), .A2(new_n1030), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n698), .B1(new_n1054), .B2(new_n684), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  AND2_X1   g0856(.A1(new_n1037), .A2(new_n1033), .ZN(new_n1057));
  INV_X1    g0857(.A(KEYINPUT42), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n1056), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(KEYINPUT107), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n1059), .A2(new_n1060), .B1(new_n1058), .B2(new_n1057), .ZN(new_n1061));
  INV_X1    g0861(.A(KEYINPUT43), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1037), .A2(new_n1033), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1055), .B1(new_n1063), .B2(KEYINPUT42), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n1064), .A2(KEYINPUT107), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1061), .A2(new_n1062), .A3(new_n1025), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1025), .A2(new_n1062), .ZN(new_n1067));
  OR2_X1    g0867(.A1(new_n1025), .A2(new_n1062), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1065), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n1064), .A2(KEYINPUT107), .B1(KEYINPUT42), .B2(new_n1063), .ZN(new_n1070));
  OAI211_X1 g0870(.A(new_n1067), .B(new_n1068), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1066), .A2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n715), .A2(new_n1043), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1072), .B(new_n1074), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n1027), .B1(new_n1053), .B2(new_n1075), .ZN(G387));
  NAND3_X1  g0876(.A1(new_n711), .A2(new_n713), .A3(new_n785), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n798), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1078), .A2(new_n724), .B1(G107), .B2(new_n224), .ZN(new_n1079));
  OR2_X1    g0879(.A1(new_n232), .A2(new_n468), .ZN(new_n1080));
  OAI211_X1 g0880(.A(new_n724), .B(new_n468), .C1(new_n277), .C2(new_n205), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT110), .B(KEYINPUT50), .Z(new_n1082));
  NOR3_X1   g0882(.A1(new_n1082), .A2(G50), .A3(new_n271), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1082), .B1(G50), .B2(new_n271), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1000), .B1(new_n1084), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1079), .B1(new_n1080), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n779), .B1(new_n1087), .B2(new_n792), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n847), .A2(new_n483), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n283), .B2(new_n828), .ZN(new_n1090));
  OAI22_X1  g0890(.A1(new_n811), .A2(new_n205), .B1(new_n819), .B2(new_n273), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(KEYINPUT111), .ZN(new_n1092));
  NAND3_X1  g0892(.A1(new_n1092), .A2(new_n320), .A3(new_n1012), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n277), .A2(new_n827), .B1(new_n831), .B2(new_n271), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1091), .A2(KEYINPUT111), .ZN(new_n1095));
  NOR4_X1   g0895(.A1(new_n1090), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AND3_X1   g0896(.A1(new_n808), .A2(KEYINPUT112), .A3(G159), .ZN(new_n1097));
  AOI21_X1  g0897(.A(KEYINPUT112), .B1(new_n808), .B2(G159), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1096), .B1(new_n1097), .B2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n817), .A2(G116), .B1(new_n820), .B2(G326), .ZN(new_n1100));
  INV_X1    g0900(.A(G283), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n811), .A2(new_n576), .B1(new_n822), .B2(new_n1101), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(G303), .A2(new_n844), .B1(new_n832), .B2(G311), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n1013), .B2(new_n828), .C1(new_n807), .C2(new_n829), .ZN(new_n1104));
  INV_X1    g0904(.A(KEYINPUT48), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1102), .B1(new_n1104), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1105), .B2(new_n1104), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT49), .ZN(new_n1108));
  OAI211_X1 g0908(.A(new_n1011), .B(new_n1100), .C1(new_n1107), .C2(new_n1108), .ZN(new_n1109));
  AND2_X1   g0909(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1099), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1088), .B1(new_n1111), .B2(new_n790), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1029), .A2(new_n778), .B1(new_n1077), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n749), .A2(new_n772), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1029), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1116), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n722), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1113), .B1(new_n1117), .B2(new_n1118), .ZN(G393));
  NAND2_X1  g0919(.A1(new_n773), .A2(new_n1029), .ZN(new_n1120));
  OR4_X1    g0920(.A1(new_n723), .A2(new_n1120), .A3(new_n1048), .A4(new_n1047), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1118), .A2(new_n777), .ZN(new_n1122));
  XNOR2_X1  g0922(.A(new_n1046), .B(new_n715), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n807), .A2(new_n273), .B1(new_n881), .B2(new_n828), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1125), .B(KEYINPUT115), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(new_n1126), .B(new_n1127), .ZN(new_n1128));
  OAI21_X1  g0928(.A(new_n891), .B1(new_n1007), .B2(new_n819), .ZN(new_n1129));
  AOI211_X1 g0929(.A(new_n1011), .B(new_n1129), .C1(G68), .C2(new_n836), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n844), .A2(new_n333), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n832), .A2(G50), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n847), .A2(G77), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1128), .A2(new_n1134), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n811), .A2(new_n1101), .B1(new_n819), .B2(new_n829), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n328), .B(new_n1136), .C1(G107), .C2(new_n817), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n464), .B2(new_n822), .C1(new_n576), .C2(new_n827), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n807), .A2(new_n1013), .B1(new_n826), .B2(new_n828), .ZN(new_n1139));
  XOR2_X1   g0939(.A(new_n1139), .B(KEYINPUT52), .Z(new_n1140));
  AOI211_X1 g0940(.A(new_n1138), .B(new_n1140), .C1(G303), .C2(new_n832), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n790), .B1(new_n1135), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1043), .A2(new_n785), .ZN(new_n1143));
  OAI221_X1 g0943(.A(new_n791), .B1(new_n213), .B2(new_n224), .C1(new_n1000), .C2(new_n242), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT113), .Z(new_n1145));
  NAND4_X1  g0945(.A1(new_n1142), .A2(new_n779), .A3(new_n1143), .A4(new_n1145), .ZN(new_n1146));
  NAND3_X1  g0946(.A1(new_n1121), .A2(new_n1124), .A3(new_n1146), .ZN(G390));
  XNOR2_X1  g0947(.A(new_n969), .B(KEYINPUT116), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1148), .B1(new_n946), .B2(new_n964), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n860), .B1(new_n743), .B2(new_n871), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1149), .B1(new_n1150), .B2(new_n952), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n967), .A2(new_n968), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n952), .B1(new_n874), .B2(new_n869), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1152), .B1(new_n1153), .B2(new_n970), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n769), .A2(G330), .A3(new_n871), .A4(new_n953), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1155), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AND3_X1   g0958(.A1(new_n686), .A2(new_n733), .A3(new_n734), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n733), .B1(new_n686), .B2(new_n734), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1159), .A2(new_n1160), .A3(new_n736), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n741), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n678), .A2(new_n1162), .ZN(new_n1163));
  OAI211_X1 g0963(.A(new_n706), .B(new_n871), .C1(new_n1161), .C2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n871), .B(G330), .C1(new_n979), .C2(new_n982), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(new_n952), .ZN(new_n1166));
  NAND4_X1  g0966(.A1(new_n1164), .A2(new_n869), .A3(new_n1155), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1155), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n874), .A2(new_n869), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1167), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n459), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n771), .A2(new_n1172), .ZN(new_n1173));
  NAND4_X1  g0973(.A1(new_n914), .A2(new_n1171), .A3(new_n666), .A4(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n723), .B1(new_n1158), .B2(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT117), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1155), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1151), .A2(new_n1154), .A3(new_n1155), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1177), .B1(new_n1182), .B2(new_n1174), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1177), .B(new_n1174), .C1(new_n1156), .C2(new_n1157), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1184), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1176), .B1(new_n1183), .B2(new_n1185), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1152), .A2(new_n783), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n808), .A2(G128), .B1(G132), .B2(new_n840), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT118), .Z(new_n1189));
  INV_X1    g0989(.A(G125), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n328), .B1(new_n819), .B2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1191), .B1(G50), .B2(new_n817), .ZN(new_n1192));
  AOI21_X1  g0992(.A(KEYINPUT53), .B1(new_n836), .B2(G150), .ZN(new_n1193));
  AND3_X1   g0993(.A1(new_n836), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1194));
  OAI221_X1 g0994(.A(new_n1192), .B1(new_n882), .B2(new_n831), .C1(new_n1193), .C2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n847), .A2(G159), .ZN(new_n1196));
  XNOR2_X1  g0996(.A(KEYINPUT54), .B(G143), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n827), .B2(new_n1197), .ZN(new_n1198));
  NOR3_X1   g0998(.A1(new_n1189), .A2(new_n1195), .A3(new_n1198), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(new_n817), .A2(G68), .B1(new_n820), .B2(G294), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1133), .A2(new_n255), .A3(new_n837), .A4(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n844), .A2(G97), .B1(new_n840), .B2(G116), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n207), .B2(new_n831), .ZN(new_n1203));
  AOI211_X1 g1003(.A(new_n1201), .B(new_n1203), .C1(G283), .C2(new_n808), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n790), .B1(new_n1199), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n780), .B1(new_n898), .B2(new_n271), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1187), .A2(new_n1205), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1158), .B2(new_n778), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1186), .A2(new_n1208), .ZN(G378));
  INV_X1    g1009(.A(KEYINPUT57), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n914), .A2(new_n666), .A3(new_n1173), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n1211), .B1(new_n1158), .B2(new_n1175), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n302), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1213), .A2(new_n286), .A3(new_n924), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n302), .B1(new_n287), .B2(new_n696), .ZN(new_n1215));
  XNOR2_X1  g1015(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1216));
  AND3_X1   g1016(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1216), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1218));
  OR2_X1    g1018(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n990), .B(G330), .C1(new_n984), .C2(KEYINPUT40), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT120), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1224));
  AND2_X1   g1024(.A1(new_n1224), .A2(new_n972), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1224), .A2(new_n972), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1223), .B1(new_n1225), .B2(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n971), .A2(new_n960), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1228), .B(new_n959), .C1(new_n1221), .C2(new_n1220), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1224), .A2(new_n972), .ZN(new_n1230));
  NAND4_X1  g1030(.A1(new_n1229), .A2(new_n1222), .A3(new_n1219), .A4(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1210), .B1(new_n1212), .B2(new_n1232), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1211), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n1182), .B2(new_n1174), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1235), .A2(KEYINPUT57), .A3(new_n1231), .A4(new_n1227), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1233), .A2(new_n722), .A3(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1219), .A2(new_n784), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n780), .B1(new_n898), .B2(new_n283), .ZN(new_n1239));
  NOR2_X1   g1039(.A1(new_n831), .A2(new_n885), .ZN(new_n1240));
  AND2_X1   g1040(.A1(new_n847), .A2(G150), .ZN(new_n1241));
  AOI211_X1 g1041(.A(new_n1240), .B(new_n1241), .C1(G128), .C2(new_n840), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1197), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n844), .A2(G137), .B1(new_n836), .B2(new_n1243), .ZN(new_n1244));
  OAI211_X1 g1044(.A(new_n1242), .B(new_n1244), .C1(new_n1190), .C2(new_n807), .ZN(new_n1245));
  OR2_X1    g1045(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(KEYINPUT59), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n817), .A2(G159), .ZN(new_n1248));
  AOI211_X1 g1048(.A(G33), .B(G41), .C1(new_n820), .C2(G124), .ZN(new_n1249));
  AND4_X1   g1049(.A1(new_n1246), .A2(new_n1247), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  OAI22_X1  g1050(.A1(new_n811), .A2(new_n205), .B1(new_n819), .B2(new_n1101), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(G58), .B2(new_n817), .ZN(new_n1252));
  NOR2_X1   g1052(.A1(new_n320), .A2(G41), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1252), .A2(new_n1004), .A3(new_n1253), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(new_n832), .A2(G97), .B1(new_n840), .B2(G107), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n420), .B2(new_n827), .ZN(new_n1256));
  AOI211_X1 g1056(.A(new_n1254), .B(new_n1256), .C1(G116), .C2(new_n808), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n283), .B1(G33), .B2(G41), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1257), .A2(KEYINPUT58), .B1(new_n1253), .B2(new_n1258), .ZN(new_n1259));
  XNOR2_X1  g1059(.A(new_n1259), .B(KEYINPUT119), .ZN(new_n1260));
  AOI211_X1 g1060(.A(new_n1250), .B(new_n1260), .C1(KEYINPUT58), .C2(new_n1257), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1239), .B1(new_n1261), .B2(new_n879), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1238), .A2(new_n1262), .ZN(new_n1263));
  AND2_X1   g1063(.A1(new_n1227), .A2(new_n1231), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1264), .B2(new_n778), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1237), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT121), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT121), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1237), .A2(new_n1268), .A3(new_n1265), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1267), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(new_n1270), .ZN(G375));
  INV_X1    g1071(.A(new_n1171), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1211), .A2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1052), .A3(new_n1174), .ZN(new_n1274));
  OAI22_X1  g1074(.A1(new_n207), .A2(new_n827), .B1(new_n831), .B2(new_n464), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(new_n808), .B2(G294), .ZN(new_n1276));
  XNOR2_X1  g1076(.A(new_n1276), .B(KEYINPUT122), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n840), .A2(G283), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n328), .B1(new_n817), .B2(G77), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n836), .A2(G97), .B1(new_n820), .B2(G303), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1278), .A2(new_n1089), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  AOI22_X1  g1081(.A1(new_n832), .A2(new_n1243), .B1(new_n840), .B2(G137), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n1282), .B1(new_n807), .B2(new_n885), .ZN(new_n1283));
  NOR2_X1   g1083(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1283), .A2(KEYINPUT123), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n811), .A2(new_n881), .B1(new_n816), .B2(new_n211), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1286), .B1(G128), .B2(new_n820), .ZN(new_n1287));
  OAI211_X1 g1087(.A(new_n1287), .B(new_n320), .C1(new_n273), .C2(new_n827), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1288), .B1(G50), .B2(new_n847), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1285), .A2(new_n1289), .ZN(new_n1290));
  OAI22_X1  g1090(.A1(new_n1277), .A2(new_n1281), .B1(new_n1284), .B2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(new_n790), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n780), .B1(new_n898), .B2(new_n277), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1292), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n783), .B2(new_n952), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n1171), .B2(new_n778), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1274), .A2(new_n1296), .ZN(G381));
  INV_X1    g1097(.A(new_n1208), .ZN(new_n1298));
  OAI21_X1  g1098(.A(KEYINPUT117), .B1(new_n1158), .B2(new_n1175), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1299), .A2(new_n1184), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1300), .B2(new_n1176), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(G387), .A2(G384), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1120), .A2(new_n722), .A3(new_n1116), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1303), .A2(new_n854), .A3(new_n1113), .ZN(new_n1304));
  NOR3_X1   g1104(.A1(G390), .A2(G381), .A3(new_n1304), .ZN(new_n1305));
  NAND4_X1  g1105(.A1(new_n1270), .A2(new_n1301), .A3(new_n1302), .A4(new_n1305), .ZN(G407));
  NAND2_X1  g1106(.A1(new_n697), .A2(G213), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1270), .A2(new_n1301), .A3(new_n1308), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(G407), .A2(G213), .A3(new_n1309), .ZN(G409));
  NAND3_X1  g1110(.A1(new_n1237), .A2(G378), .A3(new_n1265), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1264), .A2(new_n1052), .A3(new_n1235), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1265), .A2(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n1301), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1311), .A2(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1174), .A2(KEYINPUT60), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1316), .A2(new_n1273), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1211), .A2(KEYINPUT60), .A3(new_n1272), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1318), .A2(new_n722), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1296), .B1(new_n1317), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI211_X1 g1122(.A(new_n1296), .B(G384), .C1(new_n1317), .C2(new_n1319), .ZN(new_n1323));
  AND2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1315), .A2(new_n1307), .A3(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1325), .A2(KEYINPUT63), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1308), .B1(new_n1311), .B2(new_n1314), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT63), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1327), .A2(new_n1328), .A3(new_n1324), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1326), .A2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(G390), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(G393), .A2(G396), .ZN(new_n1332));
  AND3_X1   g1132(.A1(G387), .A2(new_n1304), .A3(new_n1332), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  AOI22_X1  g1134(.A1(G387), .A2(new_n1334), .B1(new_n1332), .B2(new_n1304), .ZN(new_n1335));
  OAI21_X1  g1135(.A(new_n1331), .B1(new_n1333), .B2(new_n1335), .ZN(new_n1336));
  NAND3_X1  g1136(.A1(G387), .A2(new_n1304), .A3(new_n1332), .ZN(new_n1337));
  AND2_X1   g1137(.A1(G387), .A2(new_n1334), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1332), .A2(new_n1304), .ZN(new_n1339));
  OAI211_X1 g1139(.A(new_n1337), .B(G390), .C1(new_n1338), .C2(new_n1339), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1336), .A2(new_n1340), .ZN(new_n1341));
  INV_X1    g1141(.A(KEYINPUT61), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1308), .A2(KEYINPUT124), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1322), .A2(new_n1323), .A3(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1308), .A2(G2897), .ZN(new_n1345));
  INV_X1    g1145(.A(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1344), .A2(new_n1346), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1322), .A2(new_n1323), .A3(new_n1345), .A4(new_n1343), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  OAI211_X1 g1149(.A(new_n1341), .B(new_n1342), .C1(new_n1327), .C2(new_n1349), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1330), .A2(new_n1351), .ZN(new_n1352));
  XNOR2_X1  g1152(.A(KEYINPUT126), .B(KEYINPUT62), .ZN(new_n1353));
  AND3_X1   g1153(.A1(new_n1327), .A2(new_n1324), .A3(new_n1353), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1342), .B1(new_n1327), .B2(new_n1349), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT126), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(KEYINPUT62), .ZN(new_n1357));
  AOI21_X1  g1157(.A(new_n1357), .B1(new_n1327), .B2(new_n1324), .ZN(new_n1358));
  NOR3_X1   g1158(.A1(new_n1354), .A2(new_n1355), .A3(new_n1358), .ZN(new_n1359));
  OAI21_X1  g1159(.A(new_n1352), .B1(new_n1359), .B2(new_n1341), .ZN(G405));
  NOR2_X1   g1160(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1361));
  AND2_X1   g1161(.A1(new_n1341), .A2(new_n1361), .ZN(new_n1362));
  NOR2_X1   g1162(.A1(new_n1341), .A2(new_n1361), .ZN(new_n1363));
  NOR2_X1   g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  NOR2_X1   g1164(.A1(new_n1270), .A2(G378), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1324), .A2(KEYINPUT127), .ZN(new_n1366));
  NAND2_X1  g1166(.A1(new_n1366), .A2(new_n1311), .ZN(new_n1367));
  NOR2_X1   g1167(.A1(new_n1365), .A2(new_n1367), .ZN(new_n1368));
  NAND2_X1  g1168(.A1(new_n1364), .A2(new_n1368), .ZN(new_n1369));
  OAI22_X1  g1169(.A1(new_n1362), .A2(new_n1363), .B1(new_n1365), .B2(new_n1367), .ZN(new_n1370));
  NAND2_X1  g1170(.A1(new_n1369), .A2(new_n1370), .ZN(G402));
endmodule


