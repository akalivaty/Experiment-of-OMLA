

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X1 U552 ( .A1(n688), .A2(n798), .ZN(n733) );
  NAND2_X1 U553 ( .A1(n733), .A2(G8), .ZN(n689) );
  INV_X1 U554 ( .A(KEYINPUT66), .ZN(n552) );
  XNOR2_X2 U555 ( .A(n526), .B(KEYINPUT65), .ZN(n548) );
  XOR2_X1 U556 ( .A(KEYINPUT100), .B(n733), .Z(n709) );
  INV_X1 U557 ( .A(KEYINPUT28), .ZN(n706) );
  INV_X1 U558 ( .A(KEYINPUT31), .ZN(n701) );
  INV_X1 U559 ( .A(KEYINPUT32), .ZN(n741) );
  XNOR2_X1 U560 ( .A(n742), .B(n741), .ZN(n750) );
  XOR2_X1 U561 ( .A(KEYINPUT99), .B(n689), .Z(n754) );
  INV_X1 U562 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U563 ( .A1(G2104), .A2(G2105), .ZN(n524) );
  NAND2_X1 U564 ( .A1(n827), .A2(n820), .ZN(n821) );
  OR2_X1 U565 ( .A1(n822), .A2(n821), .ZN(n834) );
  NOR2_X1 U566 ( .A1(n542), .A2(G651), .ZN(n652) );
  XNOR2_X1 U567 ( .A(n553), .B(n552), .ZN(n555) );
  AND2_X1 U568 ( .A1(G2105), .A2(G2104), .ZN(n884) );
  NAND2_X1 U569 ( .A1(G114), .A2(n884), .ZN(n522) );
  NOR2_X1 U570 ( .A1(n525), .A2(G2104), .ZN(n520) );
  XNOR2_X1 U571 ( .A(n520), .B(KEYINPUT64), .ZN(n885) );
  NAND2_X1 U572 ( .A1(G126), .A2(n885), .ZN(n521) );
  NAND2_X1 U573 ( .A1(n522), .A2(n521), .ZN(n523) );
  XNOR2_X1 U574 ( .A(KEYINPUT90), .B(n523), .ZN(n531) );
  XOR2_X2 U575 ( .A(KEYINPUT17), .B(n524), .Z(n881) );
  NAND2_X1 U576 ( .A1(G138), .A2(n881), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n525), .A2(G2104), .ZN(n526) );
  NAND2_X1 U578 ( .A1(G102), .A2(n548), .ZN(n527) );
  NAND2_X1 U579 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U580 ( .A(KEYINPUT91), .B(n529), .Z(n530) );
  NOR2_X1 U581 ( .A1(n531), .A2(n530), .ZN(G164) );
  INV_X1 U582 ( .A(G651), .ZN(n541) );
  NOR2_X1 U583 ( .A1(G543), .A2(n541), .ZN(n532) );
  XOR2_X1 U584 ( .A(KEYINPUT1), .B(n532), .Z(n651) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n542) );
  NAND2_X1 U586 ( .A1(G49), .A2(n652), .ZN(n534) );
  NAND2_X1 U587 ( .A1(G74), .A2(G651), .ZN(n533) );
  NAND2_X1 U588 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U589 ( .A1(n651), .A2(n535), .ZN(n536) );
  XNOR2_X1 U590 ( .A(n536), .B(KEYINPUT84), .ZN(n538) );
  NAND2_X1 U591 ( .A1(G87), .A2(n542), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n538), .A2(n537), .ZN(G288) );
  NOR2_X1 U593 ( .A1(G543), .A2(G651), .ZN(n647) );
  NAND2_X1 U594 ( .A1(G91), .A2(n647), .ZN(n540) );
  NAND2_X1 U595 ( .A1(G65), .A2(n651), .ZN(n539) );
  NAND2_X1 U596 ( .A1(n540), .A2(n539), .ZN(n545) );
  NOR2_X1 U597 ( .A1(n542), .A2(n541), .ZN(n648) );
  NAND2_X1 U598 ( .A1(n648), .A2(G78), .ZN(n543) );
  XOR2_X1 U599 ( .A(KEYINPUT70), .B(n543), .Z(n544) );
  NOR2_X1 U600 ( .A1(n545), .A2(n544), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n652), .A2(G53), .ZN(n546) );
  NAND2_X1 U602 ( .A1(n547), .A2(n546), .ZN(G299) );
  NAND2_X1 U603 ( .A1(n548), .A2(G101), .ZN(n549) );
  XOR2_X1 U604 ( .A(KEYINPUT23), .B(n549), .Z(n551) );
  NAND2_X1 U605 ( .A1(G125), .A2(n885), .ZN(n550) );
  NAND2_X1 U606 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n884), .A2(G113), .ZN(n554) );
  AND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n796) );
  NAND2_X1 U609 ( .A1(G137), .A2(n881), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT67), .B(n556), .Z(n687) );
  AND2_X1 U611 ( .A1(n796), .A2(n687), .ZN(G160) );
  NAND2_X1 U612 ( .A1(G64), .A2(n651), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G52), .A2(n652), .ZN(n557) );
  NAND2_X1 U614 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U615 ( .A1(G90), .A2(n647), .ZN(n560) );
  NAND2_X1 U616 ( .A1(G77), .A2(n648), .ZN(n559) );
  NAND2_X1 U617 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U618 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U619 ( .A1(n563), .A2(n562), .ZN(G171) );
  INV_X1 U620 ( .A(G108), .ZN(G238) );
  NAND2_X1 U621 ( .A1(G88), .A2(n647), .ZN(n565) );
  NAND2_X1 U622 ( .A1(G75), .A2(n648), .ZN(n564) );
  NAND2_X1 U623 ( .A1(n565), .A2(n564), .ZN(n569) );
  NAND2_X1 U624 ( .A1(G62), .A2(n651), .ZN(n567) );
  NAND2_X1 U625 ( .A1(G50), .A2(n652), .ZN(n566) );
  NAND2_X1 U626 ( .A1(n567), .A2(n566), .ZN(n568) );
  NOR2_X1 U627 ( .A1(n569), .A2(n568), .ZN(G166) );
  NAND2_X1 U628 ( .A1(n647), .A2(G89), .ZN(n570) );
  XNOR2_X1 U629 ( .A(n570), .B(KEYINPUT4), .ZN(n572) );
  NAND2_X1 U630 ( .A1(G76), .A2(n648), .ZN(n571) );
  NAND2_X1 U631 ( .A1(n572), .A2(n571), .ZN(n573) );
  XNOR2_X1 U632 ( .A(KEYINPUT5), .B(n573), .ZN(n580) );
  XNOR2_X1 U633 ( .A(KEYINPUT80), .B(KEYINPUT6), .ZN(n578) );
  NAND2_X1 U634 ( .A1(n652), .A2(G51), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n651), .A2(G63), .ZN(n574) );
  XOR2_X1 U636 ( .A(KEYINPUT79), .B(n574), .Z(n575) );
  NAND2_X1 U637 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U638 ( .A(n578), .B(n577), .Z(n579) );
  NAND2_X1 U639 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U640 ( .A(KEYINPUT7), .B(n581), .ZN(G168) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G94), .A2(G452), .ZN(n582) );
  XNOR2_X1 U643 ( .A(n582), .B(KEYINPUT69), .ZN(G173) );
  NAND2_X1 U644 ( .A1(G7), .A2(G661), .ZN(n583) );
  XNOR2_X1 U645 ( .A(n583), .B(KEYINPUT10), .ZN(G223) );
  XOR2_X1 U646 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n585) );
  XNOR2_X1 U647 ( .A(G223), .B(KEYINPUT71), .ZN(n836) );
  NAND2_X1 U648 ( .A1(G567), .A2(n836), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G234) );
  NAND2_X1 U650 ( .A1(G81), .A2(n647), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(KEYINPUT74), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(KEYINPUT12), .ZN(n589) );
  NAND2_X1 U653 ( .A1(G68), .A2(n648), .ZN(n588) );
  NAND2_X1 U654 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U655 ( .A(n590), .B(KEYINPUT13), .ZN(n592) );
  NAND2_X1 U656 ( .A1(G43), .A2(n652), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U658 ( .A1(G56), .A2(n651), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n593), .B(KEYINPUT14), .ZN(n594) );
  XNOR2_X1 U660 ( .A(n594), .B(KEYINPUT73), .ZN(n595) );
  NOR2_X1 U661 ( .A1(n596), .A2(n595), .ZN(n978) );
  INV_X1 U662 ( .A(n978), .ZN(n617) );
  XNOR2_X1 U663 ( .A(G860), .B(KEYINPUT75), .ZN(n612) );
  OR2_X1 U664 ( .A1(n617), .A2(n612), .ZN(G153) );
  INV_X1 U665 ( .A(G171), .ZN(G301) );
  NAND2_X1 U666 ( .A1(G79), .A2(n648), .ZN(n598) );
  NAND2_X1 U667 ( .A1(G54), .A2(n652), .ZN(n597) );
  NAND2_X1 U668 ( .A1(n598), .A2(n597), .ZN(n604) );
  NAND2_X1 U669 ( .A1(n647), .A2(G92), .ZN(n599) );
  XNOR2_X1 U670 ( .A(n599), .B(KEYINPUT76), .ZN(n601) );
  NAND2_X1 U671 ( .A1(G66), .A2(n651), .ZN(n600) );
  NAND2_X1 U672 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U673 ( .A(n602), .B(KEYINPUT77), .Z(n603) );
  NOR2_X1 U674 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT15), .B(n605), .Z(n606) );
  XOR2_X1 U676 ( .A(KEYINPUT78), .B(n606), .Z(n983) );
  NOR2_X1 U677 ( .A1(n983), .A2(G868), .ZN(n608) );
  INV_X1 U678 ( .A(G868), .ZN(n668) );
  NOR2_X1 U679 ( .A1(n668), .A2(G301), .ZN(n607) );
  NOR2_X1 U680 ( .A1(n608), .A2(n607), .ZN(G284) );
  INV_X1 U681 ( .A(G299), .ZN(n971) );
  NAND2_X1 U682 ( .A1(n971), .A2(n668), .ZN(n609) );
  XNOR2_X1 U683 ( .A(n609), .B(KEYINPUT81), .ZN(n611) );
  NOR2_X1 U684 ( .A1(n668), .A2(G286), .ZN(n610) );
  NOR2_X1 U685 ( .A1(n611), .A2(n610), .ZN(G297) );
  NAND2_X1 U686 ( .A1(n612), .A2(G559), .ZN(n613) );
  INV_X1 U687 ( .A(n983), .ZN(n636) );
  NAND2_X1 U688 ( .A1(n613), .A2(n636), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n614), .B(KEYINPUT16), .ZN(n615) );
  XNOR2_X1 U690 ( .A(KEYINPUT82), .B(n615), .ZN(G148) );
  NAND2_X1 U691 ( .A1(G868), .A2(n636), .ZN(n616) );
  NOR2_X1 U692 ( .A1(G559), .A2(n616), .ZN(n619) );
  NOR2_X1 U693 ( .A1(G868), .A2(n617), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(G282) );
  NAND2_X1 U695 ( .A1(G111), .A2(n884), .ZN(n621) );
  NAND2_X1 U696 ( .A1(G135), .A2(n881), .ZN(n620) );
  NAND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n885), .A2(G123), .ZN(n622) );
  XOR2_X1 U699 ( .A(KEYINPUT18), .B(n622), .Z(n623) );
  NOR2_X1 U700 ( .A1(n624), .A2(n623), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n548), .A2(G99), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n1013) );
  XNOR2_X1 U703 ( .A(n1013), .B(G2096), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n627), .B(KEYINPUT83), .ZN(n629) );
  INV_X1 U705 ( .A(G2100), .ZN(n628) );
  NAND2_X1 U706 ( .A1(n629), .A2(n628), .ZN(G156) );
  NAND2_X1 U707 ( .A1(G93), .A2(n647), .ZN(n631) );
  NAND2_X1 U708 ( .A1(G80), .A2(n648), .ZN(n630) );
  NAND2_X1 U709 ( .A1(n631), .A2(n630), .ZN(n635) );
  NAND2_X1 U710 ( .A1(G67), .A2(n651), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G55), .A2(n652), .ZN(n632) );
  NAND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  OR2_X1 U713 ( .A1(n635), .A2(n634), .ZN(n669) );
  NAND2_X1 U714 ( .A1(G559), .A2(n636), .ZN(n665) );
  XOR2_X1 U715 ( .A(n978), .B(n665), .Z(n637) );
  NOR2_X1 U716 ( .A1(G860), .A2(n637), .ZN(n638) );
  XOR2_X1 U717 ( .A(n669), .B(n638), .Z(G145) );
  NAND2_X1 U718 ( .A1(G86), .A2(n647), .ZN(n640) );
  NAND2_X1 U719 ( .A1(G61), .A2(n651), .ZN(n639) );
  NAND2_X1 U720 ( .A1(n640), .A2(n639), .ZN(n644) );
  NAND2_X1 U721 ( .A1(G73), .A2(n648), .ZN(n641) );
  XNOR2_X1 U722 ( .A(n641), .B(KEYINPUT85), .ZN(n642) );
  XNOR2_X1 U723 ( .A(n642), .B(KEYINPUT2), .ZN(n643) );
  NOR2_X1 U724 ( .A1(n644), .A2(n643), .ZN(n646) );
  NAND2_X1 U725 ( .A1(n652), .A2(G48), .ZN(n645) );
  NAND2_X1 U726 ( .A1(n646), .A2(n645), .ZN(G305) );
  NAND2_X1 U727 ( .A1(G85), .A2(n647), .ZN(n650) );
  NAND2_X1 U728 ( .A1(G72), .A2(n648), .ZN(n649) );
  NAND2_X1 U729 ( .A1(n650), .A2(n649), .ZN(n656) );
  NAND2_X1 U730 ( .A1(G60), .A2(n651), .ZN(n654) );
  NAND2_X1 U731 ( .A1(G47), .A2(n652), .ZN(n653) );
  NAND2_X1 U732 ( .A1(n654), .A2(n653), .ZN(n655) );
  NOR2_X1 U733 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U734 ( .A(KEYINPUT68), .B(n657), .Z(G290) );
  XOR2_X1 U735 ( .A(KEYINPUT19), .B(KEYINPUT86), .Z(n659) );
  XNOR2_X1 U736 ( .A(n978), .B(G166), .ZN(n658) );
  XNOR2_X1 U737 ( .A(n659), .B(n658), .ZN(n660) );
  INV_X1 U738 ( .A(G288), .ZN(n975) );
  XOR2_X1 U739 ( .A(n660), .B(n975), .Z(n662) );
  XNOR2_X1 U740 ( .A(G290), .B(n971), .ZN(n661) );
  XNOR2_X1 U741 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U742 ( .A(n669), .B(n663), .ZN(n664) );
  XNOR2_X1 U743 ( .A(G305), .B(n664), .ZN(n903) );
  XNOR2_X1 U744 ( .A(n903), .B(KEYINPUT87), .ZN(n666) );
  XNOR2_X1 U745 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U746 ( .A1(n667), .A2(G868), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U748 ( .A1(n671), .A2(n670), .ZN(G295) );
  NAND2_X1 U749 ( .A1(G2078), .A2(G2084), .ZN(n672) );
  XOR2_X1 U750 ( .A(KEYINPUT20), .B(n672), .Z(n673) );
  NAND2_X1 U751 ( .A1(G2090), .A2(n673), .ZN(n674) );
  XNOR2_X1 U752 ( .A(KEYINPUT21), .B(n674), .ZN(n675) );
  NAND2_X1 U753 ( .A1(n675), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G69), .A2(G120), .ZN(n676) );
  XOR2_X1 U756 ( .A(KEYINPUT89), .B(n676), .Z(n677) );
  NOR2_X1 U757 ( .A1(G238), .A2(n677), .ZN(n678) );
  NAND2_X1 U758 ( .A1(G57), .A2(n678), .ZN(n842) );
  NAND2_X1 U759 ( .A1(n842), .A2(G567), .ZN(n684) );
  NAND2_X1 U760 ( .A1(G132), .A2(G82), .ZN(n679) );
  XNOR2_X1 U761 ( .A(n679), .B(KEYINPUT22), .ZN(n680) );
  XNOR2_X1 U762 ( .A(n680), .B(KEYINPUT88), .ZN(n681) );
  NOR2_X1 U763 ( .A1(G218), .A2(n681), .ZN(n682) );
  NAND2_X1 U764 ( .A1(G96), .A2(n682), .ZN(n843) );
  NAND2_X1 U765 ( .A1(n843), .A2(G2106), .ZN(n683) );
  NAND2_X1 U766 ( .A1(n684), .A2(n683), .ZN(n844) );
  NAND2_X1 U767 ( .A1(G483), .A2(G661), .ZN(n685) );
  NOR2_X1 U768 ( .A1(n844), .A2(n685), .ZN(n840) );
  NAND2_X1 U769 ( .A1(n840), .A2(G36), .ZN(G176) );
  INV_X1 U770 ( .A(G166), .ZN(G303) );
  NOR2_X1 U771 ( .A1(G1981), .A2(G305), .ZN(n686) );
  XNOR2_X1 U772 ( .A(KEYINPUT24), .B(n686), .ZN(n690) );
  AND2_X1 U773 ( .A1(n687), .A2(G40), .ZN(n795) );
  AND2_X1 U774 ( .A1(n796), .A2(n795), .ZN(n688) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n798) );
  INV_X1 U776 ( .A(n754), .ZN(n771) );
  NAND2_X1 U777 ( .A1(n690), .A2(n771), .ZN(n756) );
  NOR2_X1 U778 ( .A1(G1966), .A2(n754), .ZN(n746) );
  NOR2_X1 U779 ( .A1(G2084), .A2(n733), .ZN(n743) );
  NOR2_X1 U780 ( .A1(n746), .A2(n743), .ZN(n691) );
  XNOR2_X1 U781 ( .A(n691), .B(KEYINPUT102), .ZN(n692) );
  NAND2_X1 U782 ( .A1(n692), .A2(G8), .ZN(n693) );
  XNOR2_X1 U783 ( .A(n693), .B(KEYINPUT30), .ZN(n694) );
  NOR2_X1 U784 ( .A1(G168), .A2(n694), .ZN(n700) );
  XOR2_X1 U785 ( .A(G2078), .B(KEYINPUT25), .Z(n931) );
  INV_X1 U786 ( .A(n709), .ZN(n695) );
  NOR2_X1 U787 ( .A1(n931), .A2(n695), .ZN(n696) );
  XNOR2_X1 U788 ( .A(n696), .B(KEYINPUT101), .ZN(n698) );
  INV_X1 U789 ( .A(n733), .ZN(n714) );
  OR2_X1 U790 ( .A1(G1961), .A2(n714), .ZN(n697) );
  NAND2_X1 U791 ( .A1(n698), .A2(n697), .ZN(n727) );
  NOR2_X1 U792 ( .A1(G171), .A2(n727), .ZN(n699) );
  NOR2_X1 U793 ( .A1(n700), .A2(n699), .ZN(n702) );
  XNOR2_X1 U794 ( .A(n702), .B(n701), .ZN(n731) );
  NAND2_X1 U795 ( .A1(G2072), .A2(n709), .ZN(n703) );
  XNOR2_X1 U796 ( .A(n703), .B(KEYINPUT27), .ZN(n705) );
  INV_X1 U797 ( .A(G1956), .ZN(n945) );
  NOR2_X1 U798 ( .A1(n709), .A2(n945), .ZN(n704) );
  NOR2_X1 U799 ( .A1(n705), .A2(n704), .ZN(n708) );
  NOR2_X1 U800 ( .A1(n708), .A2(n971), .ZN(n707) );
  XNOR2_X1 U801 ( .A(n707), .B(n706), .ZN(n725) );
  NAND2_X1 U802 ( .A1(n708), .A2(n971), .ZN(n723) );
  NAND2_X1 U803 ( .A1(G2067), .A2(n709), .ZN(n711) );
  NAND2_X1 U804 ( .A1(G1348), .A2(n733), .ZN(n710) );
  NAND2_X1 U805 ( .A1(n711), .A2(n710), .ZN(n719) );
  NAND2_X1 U806 ( .A1(n983), .A2(n719), .ZN(n713) );
  NAND2_X1 U807 ( .A1(G1341), .A2(n733), .ZN(n712) );
  NAND2_X1 U808 ( .A1(n713), .A2(n712), .ZN(n718) );
  NAND2_X1 U809 ( .A1(n714), .A2(G1996), .ZN(n715) );
  XNOR2_X1 U810 ( .A(n715), .B(KEYINPUT26), .ZN(n716) );
  NAND2_X1 U811 ( .A1(n716), .A2(n978), .ZN(n717) );
  NOR2_X1 U812 ( .A1(n718), .A2(n717), .ZN(n721) );
  NOR2_X1 U813 ( .A1(n983), .A2(n719), .ZN(n720) );
  NOR2_X1 U814 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U815 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U816 ( .A1(n725), .A2(n724), .ZN(n726) );
  XOR2_X1 U817 ( .A(KEYINPUT29), .B(n726), .Z(n729) );
  NAND2_X1 U818 ( .A1(n727), .A2(G171), .ZN(n728) );
  NAND2_X1 U819 ( .A1(n729), .A2(n728), .ZN(n730) );
  NAND2_X1 U820 ( .A1(n731), .A2(n730), .ZN(n744) );
  AND2_X1 U821 ( .A1(G286), .A2(G8), .ZN(n732) );
  NAND2_X1 U822 ( .A1(n744), .A2(n732), .ZN(n740) );
  INV_X1 U823 ( .A(G8), .ZN(n738) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n754), .ZN(n735) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U826 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U827 ( .A1(n736), .A2(G303), .ZN(n737) );
  OR2_X1 U828 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U830 ( .A1(G8), .A2(n743), .ZN(n748) );
  INV_X1 U831 ( .A(n744), .ZN(n745) );
  NOR2_X1 U832 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U833 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U834 ( .A1(n750), .A2(n749), .ZN(n765) );
  NOR2_X1 U835 ( .A1(G2090), .A2(G303), .ZN(n751) );
  NAND2_X1 U836 ( .A1(G8), .A2(n751), .ZN(n752) );
  NAND2_X1 U837 ( .A1(n765), .A2(n752), .ZN(n753) );
  NAND2_X1 U838 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U839 ( .A1(n756), .A2(n755), .ZN(n781) );
  NOR2_X1 U840 ( .A1(G1971), .A2(G303), .ZN(n757) );
  XNOR2_X1 U841 ( .A(KEYINPUT103), .B(n757), .ZN(n763) );
  INV_X1 U842 ( .A(G1976), .ZN(n974) );
  NAND2_X1 U843 ( .A1(n974), .A2(n975), .ZN(n762) );
  NAND2_X1 U844 ( .A1(n975), .A2(KEYINPUT33), .ZN(n758) );
  NOR2_X1 U845 ( .A1(G1976), .A2(n758), .ZN(n759) );
  NAND2_X1 U846 ( .A1(n759), .A2(n771), .ZN(n770) );
  INV_X1 U847 ( .A(n770), .ZN(n761) );
  INV_X1 U848 ( .A(KEYINPUT33), .ZN(n760) );
  OR2_X1 U849 ( .A1(n761), .A2(n760), .ZN(n769) );
  AND2_X1 U850 ( .A1(n762), .A2(n769), .ZN(n766) );
  AND2_X1 U851 ( .A1(n763), .A2(n766), .ZN(n764) );
  NAND2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n779) );
  INV_X1 U853 ( .A(n766), .ZN(n768) );
  NAND2_X1 U854 ( .A1(G288), .A2(G1976), .ZN(n767) );
  NOR2_X1 U855 ( .A1(n768), .A2(n767), .ZN(n777) );
  INV_X1 U856 ( .A(n769), .ZN(n773) );
  AND2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n772) );
  OR2_X1 U858 ( .A1(n773), .A2(n772), .ZN(n775) );
  XNOR2_X1 U859 ( .A(G1981), .B(G305), .ZN(n989) );
  INV_X1 U860 ( .A(n989), .ZN(n774) );
  NAND2_X1 U861 ( .A1(n775), .A2(n774), .ZN(n776) );
  NOR2_X1 U862 ( .A1(n777), .A2(n776), .ZN(n778) );
  AND2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n780) );
  NOR2_X1 U864 ( .A1(n781), .A2(n780), .ZN(n782) );
  XNOR2_X1 U865 ( .A(n782), .B(KEYINPUT104), .ZN(n822) );
  XNOR2_X1 U866 ( .A(KEYINPUT37), .B(G2067), .ZN(n829) );
  NAND2_X1 U867 ( .A1(G140), .A2(n881), .ZN(n784) );
  NAND2_X1 U868 ( .A1(G104), .A2(n548), .ZN(n783) );
  NAND2_X1 U869 ( .A1(n784), .A2(n783), .ZN(n786) );
  XOR2_X1 U870 ( .A(KEYINPUT93), .B(KEYINPUT34), .Z(n785) );
  XNOR2_X1 U871 ( .A(n786), .B(n785), .ZN(n792) );
  NAND2_X1 U872 ( .A1(n884), .A2(G116), .ZN(n787) );
  XNOR2_X1 U873 ( .A(n787), .B(KEYINPUT94), .ZN(n789) );
  NAND2_X1 U874 ( .A1(G128), .A2(n885), .ZN(n788) );
  NAND2_X1 U875 ( .A1(n789), .A2(n788), .ZN(n790) );
  XOR2_X1 U876 ( .A(KEYINPUT35), .B(n790), .Z(n791) );
  NOR2_X1 U877 ( .A1(n792), .A2(n791), .ZN(n793) );
  XOR2_X1 U878 ( .A(n793), .B(KEYINPUT95), .Z(n794) );
  XNOR2_X1 U879 ( .A(KEYINPUT36), .B(n794), .ZN(n897) );
  NOR2_X1 U880 ( .A1(n829), .A2(n897), .ZN(n1021) );
  NAND2_X1 U881 ( .A1(n796), .A2(n795), .ZN(n797) );
  NOR2_X1 U882 ( .A1(n798), .A2(n797), .ZN(n831) );
  NAND2_X1 U883 ( .A1(n1021), .A2(n831), .ZN(n827) );
  NAND2_X1 U884 ( .A1(G107), .A2(n884), .ZN(n800) );
  NAND2_X1 U885 ( .A1(G119), .A2(n885), .ZN(n799) );
  NAND2_X1 U886 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U887 ( .A1(n881), .A2(G131), .ZN(n801) );
  XOR2_X1 U888 ( .A(KEYINPUT96), .B(n801), .Z(n802) );
  NOR2_X1 U889 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U890 ( .A1(n548), .A2(G95), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n899) );
  NAND2_X1 U892 ( .A1(n899), .A2(G1991), .ZN(n816) );
  NAND2_X1 U893 ( .A1(n548), .A2(G105), .ZN(n806) );
  XNOR2_X1 U894 ( .A(n806), .B(KEYINPUT38), .ZN(n808) );
  NAND2_X1 U895 ( .A1(G129), .A2(n885), .ZN(n807) );
  NAND2_X1 U896 ( .A1(n808), .A2(n807), .ZN(n811) );
  NAND2_X1 U897 ( .A1(G117), .A2(n884), .ZN(n809) );
  XNOR2_X1 U898 ( .A(KEYINPUT97), .B(n809), .ZN(n810) );
  NOR2_X1 U899 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U900 ( .A(n812), .B(KEYINPUT98), .ZN(n814) );
  NAND2_X1 U901 ( .A1(G141), .A2(n881), .ZN(n813) );
  NAND2_X1 U902 ( .A1(n814), .A2(n813), .ZN(n896) );
  NAND2_X1 U903 ( .A1(n896), .A2(G1996), .ZN(n815) );
  NAND2_X1 U904 ( .A1(n816), .A2(n815), .ZN(n1012) );
  INV_X1 U905 ( .A(n1012), .ZN(n818) );
  XOR2_X1 U906 ( .A(KEYINPUT92), .B(G1986), .Z(n817) );
  XNOR2_X1 U907 ( .A(G290), .B(n817), .ZN(n986) );
  NAND2_X1 U908 ( .A1(n818), .A2(n986), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n819), .A2(n831), .ZN(n820) );
  NOR2_X1 U910 ( .A1(G1996), .A2(n896), .ZN(n1009) );
  NOR2_X1 U911 ( .A1(G1986), .A2(G290), .ZN(n823) );
  NOR2_X1 U912 ( .A1(G1991), .A2(n899), .ZN(n1016) );
  NOR2_X1 U913 ( .A1(n823), .A2(n1016), .ZN(n824) );
  NOR2_X1 U914 ( .A1(n1012), .A2(n824), .ZN(n825) );
  NOR2_X1 U915 ( .A1(n1009), .A2(n825), .ZN(n826) );
  XNOR2_X1 U916 ( .A(KEYINPUT39), .B(n826), .ZN(n828) );
  NAND2_X1 U917 ( .A1(n828), .A2(n827), .ZN(n830) );
  NAND2_X1 U918 ( .A1(n829), .A2(n897), .ZN(n1025) );
  NAND2_X1 U919 ( .A1(n830), .A2(n1025), .ZN(n832) );
  NAND2_X1 U920 ( .A1(n832), .A2(n831), .ZN(n833) );
  NAND2_X1 U921 ( .A1(n834), .A2(n833), .ZN(n835) );
  XNOR2_X1 U922 ( .A(KEYINPUT40), .B(n835), .ZN(G329) );
  NAND2_X1 U923 ( .A1(n836), .A2(G2106), .ZN(n837) );
  XOR2_X1 U924 ( .A(KEYINPUT105), .B(n837), .Z(G217) );
  AND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n838) );
  NAND2_X1 U926 ( .A1(G661), .A2(n838), .ZN(G259) );
  NAND2_X1 U927 ( .A1(G3), .A2(G1), .ZN(n839) );
  XNOR2_X1 U928 ( .A(KEYINPUT106), .B(n839), .ZN(n841) );
  NAND2_X1 U929 ( .A1(n841), .A2(n840), .ZN(G188) );
  XNOR2_X1 U930 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  INV_X1 U932 ( .A(G132), .ZN(G219) );
  INV_X1 U933 ( .A(G82), .ZN(G220) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n843), .A2(n842), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  INV_X1 U937 ( .A(n844), .ZN(G319) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n846) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n845) );
  XNOR2_X1 U940 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2090), .Z(n848) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n847) );
  XNOR2_X1 U943 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U944 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n851) );
  XNOR2_X1 U946 ( .A(n852), .B(n851), .ZN(G227) );
  XOR2_X1 U947 ( .A(G1981), .B(G1956), .Z(n854) );
  XNOR2_X1 U948 ( .A(G1966), .B(G1961), .ZN(n853) );
  XNOR2_X1 U949 ( .A(n854), .B(n853), .ZN(n855) );
  XOR2_X1 U950 ( .A(n855), .B(G2474), .Z(n857) );
  XNOR2_X1 U951 ( .A(G1991), .B(G1996), .ZN(n856) );
  XNOR2_X1 U952 ( .A(n857), .B(n856), .ZN(n861) );
  XOR2_X1 U953 ( .A(KEYINPUT41), .B(G1976), .Z(n859) );
  XNOR2_X1 U954 ( .A(G1986), .B(G1971), .ZN(n858) );
  XNOR2_X1 U955 ( .A(n859), .B(n858), .ZN(n860) );
  XNOR2_X1 U956 ( .A(n861), .B(n860), .ZN(G229) );
  NAND2_X1 U957 ( .A1(G112), .A2(n884), .ZN(n862) );
  XNOR2_X1 U958 ( .A(n862), .B(KEYINPUT108), .ZN(n869) );
  NAND2_X1 U959 ( .A1(G136), .A2(n881), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G100), .A2(n548), .ZN(n863) );
  NAND2_X1 U961 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U962 ( .A1(n885), .A2(G124), .ZN(n865) );
  XOR2_X1 U963 ( .A(KEYINPUT44), .B(n865), .Z(n866) );
  NOR2_X1 U964 ( .A1(n867), .A2(n866), .ZN(n868) );
  NAND2_X1 U965 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U966 ( .A(KEYINPUT109), .B(n870), .ZN(G162) );
  XOR2_X1 U967 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n871) );
  XNOR2_X1 U968 ( .A(n1013), .B(n871), .ZN(n880) );
  NAND2_X1 U969 ( .A1(G118), .A2(n884), .ZN(n873) );
  NAND2_X1 U970 ( .A1(G130), .A2(n885), .ZN(n872) );
  NAND2_X1 U971 ( .A1(n873), .A2(n872), .ZN(n878) );
  NAND2_X1 U972 ( .A1(G142), .A2(n881), .ZN(n875) );
  NAND2_X1 U973 ( .A1(G106), .A2(n548), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U975 ( .A(KEYINPUT45), .B(n876), .Z(n877) );
  NOR2_X1 U976 ( .A1(n878), .A2(n877), .ZN(n879) );
  XOR2_X1 U977 ( .A(n880), .B(n879), .Z(n893) );
  NAND2_X1 U978 ( .A1(G139), .A2(n881), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G103), .A2(n548), .ZN(n882) );
  NAND2_X1 U980 ( .A1(n883), .A2(n882), .ZN(n890) );
  NAND2_X1 U981 ( .A1(G115), .A2(n884), .ZN(n887) );
  NAND2_X1 U982 ( .A1(G127), .A2(n885), .ZN(n886) );
  NAND2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U984 ( .A(KEYINPUT47), .B(n888), .Z(n889) );
  NOR2_X1 U985 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U986 ( .A(KEYINPUT110), .B(n891), .Z(n1004) );
  XNOR2_X1 U987 ( .A(n1004), .B(G162), .ZN(n892) );
  XNOR2_X1 U988 ( .A(n893), .B(n892), .ZN(n894) );
  XOR2_X1 U989 ( .A(G160), .B(n894), .Z(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n901) );
  XOR2_X1 U991 ( .A(G164), .B(n897), .Z(n898) );
  XNOR2_X1 U992 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U993 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U994 ( .A1(G37), .A2(n902), .ZN(G395) );
  XOR2_X1 U995 ( .A(n903), .B(G286), .Z(n905) );
  XNOR2_X1 U996 ( .A(G171), .B(n983), .ZN(n904) );
  XNOR2_X1 U997 ( .A(n905), .B(n904), .ZN(n906) );
  NOR2_X1 U998 ( .A1(G37), .A2(n906), .ZN(n907) );
  XOR2_X1 U999 ( .A(KEYINPUT111), .B(n907), .Z(G397) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2430), .Z(n909) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2443), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(n909), .B(n908), .ZN(n915) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n911) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n910) );
  XNOR2_X1 U1005 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2427), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  XOR2_X1 U1008 ( .A(n915), .B(n914), .Z(n916) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n916), .ZN(n922) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n922), .ZN(n919) );
  NOR2_X1 U1011 ( .A1(G227), .A2(G229), .ZN(n917) );
  XNOR2_X1 U1012 ( .A(KEYINPUT49), .B(n917), .ZN(n918) );
  NOR2_X1 U1013 ( .A1(n919), .A2(n918), .ZN(n921) );
  NOR2_X1 U1014 ( .A1(G395), .A2(G397), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(n921), .A2(n920), .ZN(G225) );
  INV_X1 U1016 ( .A(G225), .ZN(G308) );
  INV_X1 U1017 ( .A(G96), .ZN(G221) );
  INV_X1 U1018 ( .A(G57), .ZN(G237) );
  INV_X1 U1019 ( .A(n922), .ZN(G401) );
  XNOR2_X1 U1020 ( .A(G1991), .B(G25), .ZN(n924) );
  XNOR2_X1 U1021 ( .A(G33), .B(G2072), .ZN(n923) );
  NOR2_X1 U1022 ( .A1(n924), .A2(n923), .ZN(n930) );
  XOR2_X1 U1023 ( .A(G1996), .B(G32), .Z(n925) );
  NAND2_X1 U1024 ( .A1(n925), .A2(G28), .ZN(n928) );
  XNOR2_X1 U1025 ( .A(KEYINPUT116), .B(G2067), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G26), .B(n926), .ZN(n927) );
  NOR2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n933) );
  XNOR2_X1 U1029 ( .A(G27), .B(n931), .ZN(n932) );
  NOR2_X1 U1030 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n934), .B(KEYINPUT117), .ZN(n935) );
  XNOR2_X1 U1032 ( .A(n935), .B(KEYINPUT53), .ZN(n938) );
  XOR2_X1 U1033 ( .A(G2084), .B(G34), .Z(n936) );
  XNOR2_X1 U1034 ( .A(KEYINPUT54), .B(n936), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n940) );
  XNOR2_X1 U1036 ( .A(G35), .B(G2090), .ZN(n939) );
  NOR2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1038 ( .A(KEYINPUT55), .B(n941), .Z(n943) );
  XNOR2_X1 U1039 ( .A(G29), .B(KEYINPUT118), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n1002) );
  XNOR2_X1 U1041 ( .A(G5), .B(G1961), .ZN(n944) );
  XNOR2_X1 U1042 ( .A(n944), .B(KEYINPUT121), .ZN(n967) );
  XOR2_X1 U1043 ( .A(G1966), .B(G21), .Z(n957) );
  XNOR2_X1 U1044 ( .A(n945), .B(G20), .ZN(n953) );
  XOR2_X1 U1045 ( .A(G1341), .B(G19), .Z(n948) );
  XOR2_X1 U1046 ( .A(KEYINPUT122), .B(G6), .Z(n946) );
  XNOR2_X1 U1047 ( .A(G1981), .B(n946), .ZN(n947) );
  NAND2_X1 U1048 ( .A1(n948), .A2(n947), .ZN(n951) );
  XOR2_X1 U1049 ( .A(KEYINPUT59), .B(G1348), .Z(n949) );
  XNOR2_X1 U1050 ( .A(G4), .B(n949), .ZN(n950) );
  NOR2_X1 U1051 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(n953), .A2(n952), .ZN(n954) );
  XNOR2_X1 U1053 ( .A(n954), .B(KEYINPUT60), .ZN(n955) );
  XNOR2_X1 U1054 ( .A(n955), .B(KEYINPUT123), .ZN(n956) );
  NAND2_X1 U1055 ( .A1(n957), .A2(n956), .ZN(n965) );
  XOR2_X1 U1056 ( .A(G1971), .B(G22), .Z(n959) );
  XNOR2_X1 U1057 ( .A(n974), .B(G23), .ZN(n958) );
  NAND2_X1 U1058 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1059 ( .A(G24), .B(G1986), .ZN(n960) );
  NOR2_X1 U1060 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(n962), .Z(n963) );
  XNOR2_X1 U1062 ( .A(KEYINPUT124), .B(n963), .ZN(n964) );
  NOR2_X1 U1063 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1064 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1065 ( .A(n968), .B(KEYINPUT125), .Z(n969) );
  XNOR2_X1 U1066 ( .A(KEYINPUT61), .B(n969), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(G16), .A2(n970), .ZN(n998) );
  XOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .Z(n996) );
  XNOR2_X1 U1069 ( .A(G166), .B(G1971), .ZN(n973) );
  XNOR2_X1 U1070 ( .A(n971), .B(G1956), .ZN(n972) );
  NAND2_X1 U1071 ( .A1(n973), .A2(n972), .ZN(n977) );
  XNOR2_X1 U1072 ( .A(n975), .B(n974), .ZN(n976) );
  NOR2_X1 U1073 ( .A1(n977), .A2(n976), .ZN(n982) );
  XOR2_X1 U1074 ( .A(n978), .B(G1341), .Z(n980) );
  XOR2_X1 U1075 ( .A(G171), .B(G1961), .Z(n979) );
  NOR2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NAND2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(G1348), .B(n983), .ZN(n984) );
  NOR2_X1 U1079 ( .A1(n985), .A2(n984), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n987), .A2(n986), .ZN(n993) );
  XOR2_X1 U1081 ( .A(G168), .B(G1966), .Z(n988) );
  NOR2_X1 U1082 ( .A1(n989), .A2(n988), .ZN(n990) );
  XOR2_X1 U1083 ( .A(KEYINPUT119), .B(n990), .Z(n991) );
  XNOR2_X1 U1084 ( .A(n991), .B(KEYINPUT57), .ZN(n992) );
  NOR2_X1 U1085 ( .A1(n993), .A2(n992), .ZN(n994) );
  XNOR2_X1 U1086 ( .A(n994), .B(KEYINPUT120), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NOR2_X1 U1088 ( .A1(n998), .A2(n997), .ZN(n999) );
  XNOR2_X1 U1089 ( .A(KEYINPUT126), .B(n999), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1000), .A2(G11), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(n1003), .B(KEYINPUT127), .ZN(n1034) );
  INV_X1 U1093 ( .A(G29), .ZN(n1032) );
  XOR2_X1 U1094 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n1028) );
  XOR2_X1 U1095 ( .A(G164), .B(G2078), .Z(n1006) );
  XNOR2_X1 U1096 ( .A(G2072), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XOR2_X1 U1098 ( .A(KEYINPUT50), .B(n1007), .Z(n1024) );
  XOR2_X1 U1099 ( .A(G2090), .B(G162), .Z(n1008) );
  NOR2_X1 U1100 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1101 ( .A(n1010), .B(KEYINPUT51), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1019) );
  XNOR2_X1 U1103 ( .A(G160), .B(G2084), .ZN(n1014) );
  NAND2_X1 U1104 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1105 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  XNOR2_X1 U1106 ( .A(n1017), .B(KEYINPUT112), .ZN(n1018) );
  NAND2_X1 U1107 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT113), .B(n1022), .ZN(n1023) );
  NOR2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1026) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1028), .B(n1027), .ZN(n1029) );
  XNOR2_X1 U1113 ( .A(n1029), .B(KEYINPUT52), .ZN(n1030) );
  NOR2_X1 U1114 ( .A1(KEYINPUT55), .A2(n1030), .ZN(n1031) );
  NOR2_X1 U1115 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1116 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XNOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1035), .ZN(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

