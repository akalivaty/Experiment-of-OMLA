//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n443, new_n447, new_n448, new_n451, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n555, new_n556, new_n557, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156, new_n1157, new_n1158;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XNOR2_X1  g006(.A(KEYINPUT64), .B(G2066), .ZN(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  XNOR2_X1  g013(.A(KEYINPUT65), .B(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT66), .Z(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT68), .ZN(G217));
  OR4_X1    g027(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(KEYINPUT69), .B(KEYINPUT2), .ZN(new_n454));
  XNOR2_X1  g029(.A(new_n453), .B(new_n454), .ZN(new_n455));
  NOR4_X1   g030(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(new_n455), .ZN(new_n459));
  INV_X1    g034(.A(new_n456), .ZN(new_n460));
  AOI22_X1  g035(.A1(new_n459), .A2(G2106), .B1(G567), .B2(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  AND2_X1   g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G101), .ZN(new_n464));
  AND3_X1   g039(.A1(KEYINPUT71), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT3), .B1(KEYINPUT71), .B2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(new_n462), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G137), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n464), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g045(.A(KEYINPUT3), .B(G2104), .ZN(new_n471));
  XNOR2_X1  g046(.A(new_n471), .B(KEYINPUT70), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n472), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n470), .B1(new_n473), .B2(new_n462), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  OAI21_X1  g050(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n462), .A2(G112), .ZN(new_n479));
  OAI21_X1  g054(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n467), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G136), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT72), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n462), .ZN(new_n487));
  INV_X1    g062(.A(G126), .ZN(new_n488));
  OAI21_X1  g063(.A(new_n487), .B1(new_n476), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g064(.A(new_n489), .B(KEYINPUT73), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n472), .A2(new_n462), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(new_n492), .A3(G138), .ZN(new_n493));
  INV_X1    g068(.A(G138), .ZN(new_n494));
  OAI21_X1  g069(.A(KEYINPUT4), .B1(new_n467), .B2(new_n494), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(G164));
  INV_X1    g071(.A(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n498), .B2(KEYINPUT74), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT74), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n501));
  OR2_X1    g076(.A1(KEYINPUT6), .A2(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(KEYINPUT6), .A2(G651), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n499), .A2(new_n501), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G88), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n498), .B1(new_n502), .B2(new_n503), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g083(.A(new_n505), .B1(new_n506), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n499), .A2(new_n501), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n510), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n511));
  INV_X1    g086(.A(G651), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n509), .A2(new_n513), .ZN(G166));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT75), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT7), .ZN(new_n517));
  OR2_X1    g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n504), .A2(G89), .ZN(new_n519));
  AND2_X1   g094(.A1(G63), .A2(G651), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n507), .A2(G51), .B1(new_n510), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n516), .A2(new_n517), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n518), .A2(new_n519), .A3(new_n521), .A4(new_n522), .ZN(G286));
  INV_X1    g098(.A(G286), .ZN(G168));
  AOI22_X1  g099(.A1(new_n504), .A2(G90), .B1(new_n507), .B2(G52), .ZN(new_n525));
  INV_X1    g100(.A(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(G77), .A2(G543), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n527), .B1(new_n510), .B2(G64), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n528), .A2(new_n512), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT76), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(new_n530), .ZN(new_n531));
  OR2_X1    g106(.A1(new_n528), .A2(new_n512), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT76), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n532), .A2(new_n533), .A3(new_n525), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G301));
  INV_X1    g111(.A(G301), .ZN(G171));
  INV_X1    g112(.A(G56), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n538), .B1(new_n499), .B2(new_n501), .ZN(new_n539));
  AND2_X1   g114(.A1(G68), .A2(G543), .ZN(new_n540));
  OAI21_X1  g115(.A(G651), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT77), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT77), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n543), .B(G651), .C1(new_n539), .C2(new_n540), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n504), .A2(G81), .B1(new_n507), .B2(G43), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n542), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(KEYINPUT78), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g123(.A1(new_n542), .A2(KEYINPUT78), .A3(new_n544), .A4(new_n545), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(G860), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT79), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT80), .ZN(G188));
  INV_X1    g133(.A(G65), .ZN(new_n559));
  AND3_X1   g134(.A1(new_n500), .A2(KEYINPUT5), .A3(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(KEYINPUT5), .B1(new_n500), .B2(G543), .ZN(new_n561));
  OAI21_X1  g136(.A(KEYINPUT81), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT81), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n499), .A2(new_n563), .A3(new_n501), .ZN(new_n564));
  AOI21_X1  g139(.A(new_n559), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g140(.A1(G78), .A2(G543), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(new_n567));
  OAI21_X1  g142(.A(KEYINPUT82), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  AND3_X1   g143(.A1(new_n499), .A2(new_n563), .A3(new_n501), .ZN(new_n569));
  AOI21_X1  g144(.A(new_n563), .B1(new_n499), .B2(new_n501), .ZN(new_n570));
  OAI21_X1  g145(.A(G65), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT82), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n571), .A2(new_n572), .A3(new_n566), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n568), .A2(G651), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G53), .ZN(new_n575));
  OR3_X1    g150(.A1(new_n508), .A2(KEYINPUT9), .A3(new_n575), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT9), .B1(new_n508), .B2(new_n575), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n576), .A2(new_n577), .B1(G91), .B2(new_n504), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G166), .ZN(G303));
  AOI22_X1  g155(.A1(new_n504), .A2(G87), .B1(new_n507), .B2(G49), .ZN(new_n581));
  OAI21_X1  g156(.A(G651), .B1(new_n510), .B2(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(G288));
  AOI22_X1  g158(.A1(new_n510), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n512), .ZN(new_n585));
  AOI22_X1  g160(.A1(new_n504), .A2(G86), .B1(new_n507), .B2(G48), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(G305));
  AOI22_X1  g162(.A1(new_n504), .A2(G85), .B1(new_n507), .B2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n510), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n512), .B2(new_n589), .ZN(G290));
  OAI21_X1  g165(.A(G66), .B1(new_n569), .B2(new_n570), .ZN(new_n591));
  NAND2_X1  g166(.A1(G79), .A2(G543), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n512), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g168(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n507), .A2(G54), .ZN(new_n595));
  AOI21_X1  g170(.A(KEYINPUT10), .B1(new_n504), .B2(G92), .ZN(new_n596));
  INV_X1    g171(.A(new_n596), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n595), .A3(new_n599), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(G868), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n601), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g177(.A(new_n601), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g178(.A(G299), .B(G286), .S(G868), .Z(G297));
  XOR2_X1   g179(.A(G297), .B(KEYINPUT83), .Z(G280));
  INV_X1    g180(.A(new_n598), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(new_n596), .ZN(new_n607));
  NOR2_X1   g182(.A1(new_n607), .A2(new_n593), .ZN(new_n608));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n609), .B2(G860), .ZN(G148));
  OAI21_X1  g185(.A(G868), .B1(new_n600), .B2(G559), .ZN(new_n611));
  INV_X1    g186(.A(new_n550), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G868), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n491), .A2(G2104), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT12), .ZN(new_n616));
  XOR2_X1   g191(.A(new_n616), .B(KEYINPUT13), .Z(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2100), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n482), .A2(G135), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT84), .Z(new_n620));
  NAND2_X1  g195(.A1(new_n477), .A2(G123), .ZN(new_n621));
  NOR2_X1   g196(.A1(new_n462), .A2(G111), .ZN(new_n622));
  OAI21_X1  g197(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n623));
  OAI211_X1 g198(.A(new_n620), .B(new_n621), .C1(new_n622), .C2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT85), .ZN(new_n625));
  INV_X1    g200(.A(G2096), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  NOR2_X1   g202(.A1(new_n618), .A2(new_n627), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(KEYINPUT86), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(G2427), .B(G2438), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2430), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT15), .B(G2435), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(G1341), .B(G1348), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n635), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2443), .B(G2446), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n642), .A2(G14), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(G401));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  XNOR2_X1  g221(.A(G2067), .B(G2678), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g223(.A(G2072), .B(G2078), .Z(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  OR2_X1    g225(.A1(new_n646), .A2(new_n647), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(KEYINPUT88), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n653), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(KEYINPUT17), .ZN(new_n655));
  OAI221_X1 g230(.A(new_n648), .B1(new_n650), .B2(new_n651), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  NOR2_X1   g231(.A1(new_n648), .A2(new_n649), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n660), .B(new_n626), .ZN(new_n661));
  XNOR2_X1  g236(.A(KEYINPUT89), .B(G2100), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(G227));
  XNOR2_X1  g238(.A(G1956), .B(G2474), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1961), .B(G1966), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XOR2_X1   g242(.A(new_n667), .B(KEYINPUT19), .Z(new_n668));
  NOR2_X1   g243(.A1(new_n664), .A2(new_n665), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  OAI21_X1  g245(.A(new_n666), .B1(new_n668), .B2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n668), .A2(new_n669), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT20), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n674), .A2(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(G1991), .B(G1996), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n679), .B(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(G1981), .B(G1986), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  NAND2_X1  g258(.A1(new_n625), .A2(G29), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT31), .B(G11), .ZN(new_n685));
  XOR2_X1   g260(.A(KEYINPUT98), .B(G28), .Z(new_n686));
  AOI21_X1  g261(.A(G29), .B1(new_n686), .B2(KEYINPUT30), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT99), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n690), .B1(KEYINPUT30), .B2(new_n686), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n684), .B(new_n685), .C1(new_n689), .C2(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT100), .ZN(new_n693));
  INV_X1    g268(.A(G16), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G5), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G171), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n696), .A2(G1961), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n694), .A2(G21), .ZN(new_n698));
  OAI21_X1  g273(.A(new_n698), .B1(G168), .B2(new_n694), .ZN(new_n699));
  INV_X1    g274(.A(G1966), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n699), .B(new_n700), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n693), .A2(new_n697), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n702), .A2(KEYINPUT101), .ZN(new_n703));
  NOR2_X1   g278(.A1(G29), .A2(G35), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G162), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT29), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(G2090), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n706), .A2(G2090), .ZN(new_n708));
  OR2_X1    g283(.A1(new_n696), .A2(G1961), .ZN(new_n709));
  INV_X1    g284(.A(G29), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(G32), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n482), .A2(G141), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n477), .A2(G129), .ZN(new_n713));
  NAND3_X1  g288(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n714));
  INV_X1    g289(.A(KEYINPUT26), .ZN(new_n715));
  OR2_X1    g290(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n714), .A2(new_n715), .ZN(new_n717));
  AOI22_X1  g292(.A1(new_n716), .A2(new_n717), .B1(G105), .B2(new_n463), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n712), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(KEYINPUT96), .ZN(new_n720));
  OR2_X1    g295(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n719), .A2(new_n720), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n711), .B1(new_n724), .B2(new_n710), .ZN(new_n725));
  XOR2_X1   g300(.A(KEYINPUT27), .B(G1996), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n710), .A2(G27), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n727), .B(KEYINPUT102), .ZN(new_n728));
  OAI21_X1  g303(.A(new_n728), .B1(G164), .B2(new_n710), .ZN(new_n729));
  AOI22_X1  g304(.A1(new_n725), .A2(new_n726), .B1(new_n729), .B2(G2078), .ZN(new_n730));
  NAND3_X1  g305(.A1(new_n708), .A2(new_n709), .A3(new_n730), .ZN(new_n731));
  NOR3_X1   g306(.A1(new_n703), .A2(new_n707), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n694), .A2(G23), .ZN(new_n733));
  INV_X1    g308(.A(G288), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n694), .ZN(new_n735));
  XOR2_X1   g310(.A(new_n735), .B(KEYINPUT92), .Z(new_n736));
  XOR2_X1   g311(.A(KEYINPUT33), .B(G1976), .Z(new_n737));
  OR2_X1    g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n736), .A2(new_n737), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT91), .B(G16), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n741), .A2(G22), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G166), .B2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(G1971), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n743), .B(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G6), .A2(G16), .ZN(new_n746));
  INV_X1    g321(.A(G305), .ZN(new_n747));
  AOI21_X1  g322(.A(new_n746), .B1(new_n747), .B2(G16), .ZN(new_n748));
  XOR2_X1   g323(.A(KEYINPUT32), .B(G1981), .Z(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND4_X1  g325(.A1(new_n738), .A2(new_n739), .A3(new_n745), .A4(new_n750), .ZN(new_n751));
  OR2_X1    g326(.A1(new_n751), .A2(KEYINPUT34), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(KEYINPUT34), .ZN(new_n753));
  OR2_X1    g328(.A1(G95), .A2(G2105), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n754), .B(G2104), .C1(G107), .C2(new_n462), .ZN(new_n755));
  INV_X1    g330(.A(G131), .ZN(new_n756));
  INV_X1    g331(.A(G119), .ZN(new_n757));
  OAI221_X1 g332(.A(new_n755), .B1(new_n467), .B2(new_n756), .C1(new_n757), .C2(new_n476), .ZN(new_n758));
  MUX2_X1   g333(.A(G25), .B(new_n758), .S(G29), .Z(new_n759));
  XOR2_X1   g334(.A(KEYINPUT35), .B(G1991), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  MUX2_X1   g336(.A(G24), .B(G290), .S(new_n741), .Z(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1986), .Z(new_n763));
  NAND4_X1  g338(.A1(new_n752), .A2(new_n753), .A3(new_n761), .A4(new_n763), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT93), .B(KEYINPUT36), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  INV_X1    g341(.A(new_n766), .ZN(new_n767));
  OR2_X1    g342(.A1(G104), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n769));
  INV_X1    g344(.A(G140), .ZN(new_n770));
  INV_X1    g345(.A(G128), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n769), .B1(new_n467), .B2(new_n770), .C1(new_n771), .C2(new_n476), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n772), .A2(G29), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT95), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n710), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(G2067), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(KEYINPUT24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n710), .B1(new_n780), .B2(G34), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n780), .B2(G34), .ZN(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G160), .B2(G29), .ZN(new_n783));
  OAI221_X1 g358(.A(new_n779), .B1(G2078), .B2(new_n729), .C1(G2084), .C2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n740), .A2(G20), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT23), .Z(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(G299), .B2(G16), .ZN(new_n787));
  INV_X1    g362(.A(G1956), .ZN(new_n788));
  XNOR2_X1  g363(.A(new_n787), .B(new_n788), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n741), .A2(G19), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n612), .B2(new_n741), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1341), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n694), .A2(G4), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n608), .B2(new_n694), .ZN(new_n794));
  XOR2_X1   g369(.A(KEYINPUT94), .B(G1348), .Z(new_n795));
  INV_X1    g370(.A(new_n795), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n794), .B(new_n796), .ZN(new_n797));
  NOR4_X1   g372(.A1(new_n784), .A2(new_n789), .A3(new_n792), .A4(new_n797), .ZN(new_n798));
  INV_X1    g373(.A(G2072), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n800));
  INV_X1    g375(.A(KEYINPUT25), .ZN(new_n801));
  OR2_X1    g376(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  AOI22_X1  g378(.A1(new_n482), .A2(G139), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  AOI22_X1  g379(.A1(new_n472), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n805), .B2(new_n462), .ZN(new_n806));
  INV_X1    g381(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n807), .A2(new_n710), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(new_n710), .B2(G33), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n799), .A2(new_n809), .B1(new_n783), .B2(G2084), .ZN(new_n810));
  OAI221_X1 g385(.A(new_n810), .B1(new_n799), .B2(new_n809), .C1(new_n725), .C2(new_n726), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT97), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(new_n702), .B2(KEYINPUT101), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n732), .A2(new_n767), .A3(new_n798), .A4(new_n813), .ZN(G150));
  INV_X1    g389(.A(G150), .ZN(G311));
  NAND2_X1  g390(.A1(new_n504), .A2(G93), .ZN(new_n816));
  INV_X1    g391(.A(G55), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n816), .B1(new_n817), .B2(new_n508), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n510), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n819), .A2(new_n512), .ZN(new_n820));
  NOR2_X1   g395(.A1(new_n818), .A2(new_n820), .ZN(new_n821));
  NOR2_X1   g396(.A1(new_n821), .A2(new_n551), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT37), .ZN(new_n823));
  AOI21_X1  g398(.A(new_n821), .B1(new_n548), .B2(new_n549), .ZN(new_n824));
  NOR3_X1   g399(.A1(new_n546), .A2(new_n820), .A3(new_n818), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT38), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n600), .A2(new_n609), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(KEYINPUT39), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT103), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n551), .B1(new_n829), .B2(new_n830), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n823), .B1(new_n832), .B2(new_n833), .ZN(G145));
  XNOR2_X1  g409(.A(new_n723), .B(new_n772), .ZN(new_n835));
  OAI21_X1  g410(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n836));
  INV_X1    g411(.A(G118), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n836), .B1(new_n837), .B2(G2105), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n477), .A2(G130), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT104), .Z(new_n840));
  AOI211_X1 g415(.A(new_n838), .B(new_n840), .C1(G142), .C2(new_n482), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n835), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n616), .B(new_n758), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n843), .A2(new_n844), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n489), .B1(new_n493), .B2(new_n495), .ZN(new_n847));
  NOR3_X1   g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n842), .B(new_n844), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n493), .A2(new_n495), .ZN(new_n850));
  INV_X1    g425(.A(new_n489), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NOR2_X1   g427(.A1(new_n849), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n806), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n625), .B(new_n474), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n855), .B(G162), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n847), .B1(new_n845), .B2(new_n846), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n849), .A2(new_n852), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n857), .A2(new_n858), .A3(new_n807), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n854), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(G37), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n856), .B1(new_n854), .B2(new_n859), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT40), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n864), .B(new_n865), .ZN(G395));
  XOR2_X1   g441(.A(G305), .B(G290), .Z(new_n867));
  XNOR2_X1  g442(.A(G166), .B(new_n734), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n867), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT42), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(KEYINPUT107), .B2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(KEYINPUT108), .ZN(new_n872));
  NOR2_X1   g447(.A1(new_n600), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n826), .B(new_n873), .ZN(new_n874));
  NAND2_X1  g449(.A1(G299), .A2(new_n600), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n608), .A2(new_n574), .A3(new_n578), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n875), .A2(new_n879), .A3(new_n876), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(KEYINPUT105), .ZN(new_n881));
  INV_X1    g456(.A(KEYINPUT105), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n875), .A2(new_n882), .A3(new_n876), .A4(new_n879), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT106), .ZN(new_n885));
  AOI211_X1 g460(.A(new_n885), .B(new_n879), .C1(new_n875), .C2(new_n876), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n875), .A2(new_n876), .ZN(new_n888));
  OAI21_X1  g463(.A(new_n885), .B1(new_n888), .B2(new_n879), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n884), .A2(new_n887), .A3(new_n889), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n878), .B1(new_n890), .B2(new_n874), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n872), .B(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n870), .A2(KEYINPUT107), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n892), .B(new_n893), .Z(new_n894));
  NAND2_X1  g469(.A1(new_n894), .A2(G868), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(G868), .B2(new_n821), .ZN(G295));
  OAI21_X1  g471(.A(new_n895), .B1(G868), .B2(new_n821), .ZN(G331));
  AND3_X1   g472(.A1(new_n530), .A2(new_n534), .A3(G286), .ZN(new_n898));
  AOI21_X1  g473(.A(G286), .B1(new_n530), .B2(new_n534), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n826), .A2(new_n900), .ZN(new_n901));
  OAI22_X1  g476(.A1(new_n824), .A2(new_n825), .B1(new_n898), .B2(new_n899), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n903), .A2(new_n877), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n904), .B1(new_n890), .B2(new_n903), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n869), .B1(new_n905), .B2(KEYINPUT109), .ZN(new_n906));
  AND2_X1   g481(.A1(new_n901), .A2(new_n902), .ZN(new_n907));
  AOI21_X1  g482(.A(KEYINPUT106), .B1(new_n877), .B2(KEYINPUT41), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n908), .A2(new_n886), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n909), .B2(new_n884), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT109), .ZN(new_n911));
  NOR3_X1   g486(.A1(new_n910), .A2(new_n911), .A3(new_n904), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n861), .B1(new_n906), .B2(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n869), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT110), .B1(new_n905), .B2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT110), .ZN(new_n916));
  NOR4_X1   g491(.A1(new_n910), .A2(new_n916), .A3(new_n869), .A4(new_n904), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g493(.A(KEYINPUT43), .B1(new_n913), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT111), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT111), .ZN(new_n922));
  OAI211_X1 g497(.A(new_n922), .B(KEYINPUT43), .C1(new_n913), .C2(new_n918), .ZN(new_n923));
  INV_X1    g498(.A(new_n918), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT43), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n888), .A2(new_n879), .ZN(new_n926));
  INV_X1    g501(.A(new_n880), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n903), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n877), .B2(new_n903), .ZN(new_n929));
  AOI21_X1  g504(.A(G37), .B1(new_n929), .B2(new_n869), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n924), .A2(new_n925), .A3(new_n930), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n920), .A2(new_n921), .A3(new_n923), .A4(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT112), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n925), .B1(new_n924), .B2(new_n930), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n913), .A2(new_n918), .A3(KEYINPUT43), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT44), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AND3_X1   g511(.A1(new_n932), .A2(new_n933), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n933), .B1(new_n932), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(G397));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n847), .B2(G1384), .ZN(new_n941));
  NAND2_X1  g516(.A1(G160), .A2(G40), .ZN(new_n942));
  OAI21_X1  g517(.A(KEYINPUT113), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1384), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n852), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT113), .ZN(new_n946));
  AND2_X1   g521(.A1(G160), .A2(G40), .ZN(new_n947));
  NAND4_X1  g522(.A1(new_n945), .A2(new_n946), .A3(new_n940), .A4(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n943), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT114), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n943), .A2(new_n948), .A3(KEYINPUT114), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n953), .A2(new_n723), .ZN(new_n954));
  INV_X1    g529(.A(new_n949), .ZN(new_n955));
  INV_X1    g530(.A(G1996), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT46), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n772), .B(new_n778), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n952), .ZN(new_n962));
  AOI21_X1  g537(.A(KEYINPUT114), .B1(new_n943), .B2(new_n948), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n961), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n949), .A2(G1996), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n965), .A2(KEYINPUT46), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n954), .A2(new_n959), .A3(new_n964), .A4(new_n966), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n967), .B(KEYINPUT47), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n954), .A2(new_n957), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n723), .A2(new_n956), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n964), .A2(KEYINPUT115), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT115), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n953), .A2(new_n972), .A3(new_n961), .ZN(new_n973));
  AOI22_X1  g548(.A1(new_n969), .A2(new_n970), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n760), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n758), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n758), .A2(new_n975), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n953), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NOR2_X1   g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n955), .A2(new_n979), .ZN(new_n980));
  XNOR2_X1  g555(.A(new_n980), .B(KEYINPUT48), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n974), .A2(new_n978), .A3(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n953), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n724), .B1(new_n951), .B2(new_n952), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n970), .B1(new_n984), .B2(new_n965), .ZN(new_n985));
  AOI21_X1  g560(.A(new_n972), .B1(new_n953), .B2(new_n961), .ZN(new_n986));
  AOI211_X1 g561(.A(KEYINPUT115), .B(new_n960), .C1(new_n951), .C2(new_n952), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n985), .B(new_n977), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n772), .A2(G2067), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  OAI211_X1 g566(.A(new_n968), .B(new_n982), .C1(new_n991), .C2(KEYINPUT126), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n993));
  OAI21_X1  g568(.A(KEYINPUT127), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  OR2_X1    g569(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n995));
  AND2_X1   g570(.A1(new_n968), .A2(new_n982), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(KEYINPUT126), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n995), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n994), .A2(new_n999), .ZN(new_n1000));
  AND2_X1   g575(.A1(G290), .A2(G1986), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n955), .B1(new_n979), .B2(new_n1001), .ZN(new_n1002));
  AND3_X1   g577(.A1(new_n974), .A2(new_n1002), .A3(new_n978), .ZN(new_n1003));
  INV_X1    g578(.A(G8), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n847), .A2(G1384), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n942), .B1(new_n1005), .B2(KEYINPUT45), .ZN(new_n1006));
  OAI21_X1  g581(.A(new_n940), .B1(G164), .B2(G1384), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT116), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1006), .A2(KEYINPUT116), .A3(new_n1007), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n744), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n947), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1014));
  NOR3_X1   g589(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1015));
  OR3_X1    g590(.A1(new_n1014), .A2(G2090), .A3(new_n1015), .ZN(new_n1016));
  AOI21_X1  g591(.A(new_n1004), .B1(new_n1012), .B2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g592(.A1(G166), .A2(new_n1004), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT55), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  XNOR2_X1  g595(.A(new_n1019), .B(KEYINPUT117), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n942), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1022));
  AND2_X1   g597(.A1(new_n493), .A2(new_n495), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n944), .B1(new_n1023), .B2(new_n490), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(KEYINPUT50), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1022), .A2(new_n1025), .ZN(new_n1026));
  OR2_X1    g601(.A1(new_n1026), .A2(G2090), .ZN(new_n1027));
  AOI211_X1 g602(.A(new_n1004), .B(new_n1021), .C1(new_n1012), .C2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1005), .A2(new_n947), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1029), .A2(G8), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(G1976), .B2(new_n734), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT52), .ZN(new_n1032));
  OR2_X1    g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  OAI211_X1 g608(.A(new_n1031), .B(new_n1032), .C1(G1976), .C2(new_n734), .ZN(new_n1034));
  XNOR2_X1  g609(.A(G305), .B(G1981), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT49), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1036), .A2(G8), .A3(new_n1029), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1034), .A3(new_n1037), .ZN(new_n1038));
  NOR3_X1   g613(.A1(new_n1020), .A2(new_n1028), .A3(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n788), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT56), .B(G2072), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1006), .A2(new_n1007), .A3(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1042), .A2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1046));
  XNOR2_X1  g621(.A(G299), .B(new_n1046), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1041), .B1(new_n1045), .B2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(new_n1047), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1042), .A2(new_n1044), .A3(KEYINPUT120), .A4(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g626(.A(KEYINPUT121), .B1(new_n1029), .B2(G2067), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT121), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1005), .A2(new_n947), .A3(new_n1053), .A4(new_n778), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1052), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n796), .B1(new_n1022), .B2(new_n1025), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n608), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1051), .A2(new_n1059), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT60), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n600), .A2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1062), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1026), .A2(new_n795), .ZN(new_n1064));
  INV_X1    g639(.A(new_n1062), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1064), .A2(new_n1054), .A3(new_n1052), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1063), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n600), .A2(new_n1061), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1048), .A2(new_n1070), .A3(new_n1050), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1005), .A2(KEYINPUT45), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1072), .A2(new_n1007), .A3(new_n956), .A4(new_n947), .ZN(new_n1073));
  XOR2_X1   g648(.A(KEYINPUT58), .B(G1341), .Z(new_n1074));
  NAND2_X1  g649(.A1(new_n1029), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT122), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1073), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1076), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n612), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT59), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT59), .B(new_n612), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n1069), .A2(new_n1071), .A3(new_n1081), .A4(new_n1082), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1042), .A2(new_n1049), .A3(new_n1044), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1058), .A2(KEYINPUT123), .A3(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT123), .ZN(new_n1086));
  NAND4_X1  g661(.A1(new_n1042), .A2(new_n1044), .A3(new_n1086), .A4(new_n1049), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n1070), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1060), .B1(new_n1083), .B2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n942), .B1(new_n945), .B2(new_n940), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1091), .A2(G2078), .ZN(new_n1092));
  AND2_X1   g667(.A1(new_n1072), .A2(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g668(.A(KEYINPUT124), .B(G1961), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1090), .A2(new_n1093), .B1(new_n1026), .B2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(G2078), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1096));
  OAI211_X1 g671(.A(G301), .B(new_n1095), .C1(new_n1096), .C2(KEYINPUT53), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1026), .A2(new_n1094), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1090), .B(new_n1092), .C1(new_n940), .C2(new_n1024), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(G2078), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1011), .ZN(new_n1102));
  AOI21_X1  g677(.A(KEYINPUT116), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g679(.A(new_n1100), .B1(new_n1104), .B2(new_n1091), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1097), .B1(new_n1105), .B2(G301), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1090), .B1(new_n940), .B2(new_n1024), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(new_n700), .ZN(new_n1109));
  INV_X1    g684(.A(G2084), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n1022), .A2(new_n1025), .A3(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1109), .A2(G168), .A3(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(G8), .ZN(new_n1113));
  AOI21_X1  g688(.A(G168), .B1(new_n1109), .B2(new_n1111), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT51), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT51), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1116), .A3(G8), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1106), .A2(new_n1107), .B1(new_n1115), .B2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1095), .B1(new_n1096), .B2(KEYINPUT53), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1107), .B1(new_n1119), .B2(G171), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1121));
  OAI211_X1 g696(.A(new_n1121), .B(G301), .C1(new_n1096), .C2(KEYINPUT53), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1122), .A2(KEYINPUT125), .ZN(new_n1123));
  NOR2_X1   g698(.A1(new_n1122), .A2(KEYINPUT125), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1120), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1089), .A2(new_n1118), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1127), .A2(KEYINPUT62), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1105), .A2(G301), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT62), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1115), .A2(new_n1130), .A3(new_n1117), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1128), .A2(new_n1129), .A3(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1040), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(G1976), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1037), .A2(new_n1134), .A3(new_n734), .ZN(new_n1135));
  INV_X1    g710(.A(G1981), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n747), .A2(new_n1136), .ZN(new_n1137));
  AOI21_X1  g712(.A(new_n1030), .B1(new_n1135), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1038), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1139), .B2(new_n1028), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1012), .A2(new_n1027), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1021), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1141), .A2(G8), .A3(new_n1142), .ZN(new_n1143));
  AOI211_X1 g718(.A(new_n1004), .B(G286), .C1(new_n1109), .C2(new_n1111), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1139), .A2(KEYINPUT63), .A3(new_n1143), .A4(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1141), .A2(G8), .ZN(new_n1146));
  OR2_X1    g721(.A1(new_n1146), .A2(KEYINPUT118), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1019), .B1(new_n1146), .B2(KEYINPUT118), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1145), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(KEYINPUT63), .B1(new_n1039), .B2(new_n1144), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1140), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n1003), .B1(new_n1133), .B2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1000), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g728(.A(G319), .B1(new_n643), .B2(new_n644), .ZN(new_n1155));
  NOR3_X1   g729(.A1(G229), .A2(G227), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g730(.A(new_n1156), .B1(new_n862), .B2(new_n863), .ZN(new_n1157));
  AND2_X1   g731(.A1(new_n920), .A2(new_n931), .ZN(new_n1158));
  AOI21_X1  g732(.A(new_n1157), .B1(new_n923), .B2(new_n1158), .ZN(G308));
  INV_X1    g733(.A(G308), .ZN(G225));
endmodule


