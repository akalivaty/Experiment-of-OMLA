//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 1 0 1 1 1 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n720, new_n722, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n832, new_n833, new_n834, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT11), .ZN(new_n203));
  INV_X1    g002(.A(G169gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G197gat), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n205), .B(new_n206), .ZN(new_n207));
  XOR2_X1   g006(.A(new_n207), .B(KEYINPUT12), .Z(new_n208));
  NOR2_X1   g007(.A1(G29gat), .A2(G36gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(new_n209), .B(KEYINPUT14), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT93), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G43gat), .B(G50gat), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(KEYINPUT15), .ZN(new_n215));
  INV_X1    g014(.A(G36gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT92), .B(G29gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n214), .B(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n216), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(new_n210), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n212), .A2(new_n218), .B1(new_n220), .B2(new_n215), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT94), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(G8gat), .ZN(new_n224));
  XNOR2_X1  g023(.A(G15gat), .B(G22gat), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT16), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n225), .B1(new_n226), .B2(G1gat), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n224), .B1(new_n227), .B2(KEYINPUT95), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(G1gat), .B2(new_n225), .ZN(new_n229));
  XOR2_X1   g028(.A(new_n228), .B(new_n229), .Z(new_n230));
  XNOR2_X1  g029(.A(new_n223), .B(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(G229gat), .A2(G233gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n232), .B(KEYINPUT96), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT98), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n234), .B(KEYINPUT13), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n236), .B(KEYINPUT99), .Z(new_n237));
  NOR2_X1   g036(.A1(new_n223), .A2(new_n230), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n221), .A2(KEYINPUT17), .ZN(new_n239));
  INV_X1    g038(.A(new_n223), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(KEYINPUT17), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n238), .B1(new_n241), .B2(new_n230), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(new_n233), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT18), .ZN(new_n244));
  NOR2_X1   g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n237), .A2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n208), .B1(new_n246), .B2(KEYINPUT97), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n244), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(new_n246), .B(new_n248), .C1(KEYINPUT97), .C2(new_n208), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G8gat), .B(G36gat), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n254), .B(G64gat), .ZN(new_n255));
  INV_X1    g054(.A(G92gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n255), .B(new_n256), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT88), .B(KEYINPUT38), .Z(new_n258));
  INV_X1    g057(.A(new_n258), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT37), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT77), .B(G197gat), .ZN(new_n263));
  INV_X1    g062(.A(G204gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT78), .ZN(new_n266));
  AOI22_X1  g065(.A1(new_n266), .A2(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n267), .B1(new_n266), .B2(KEYINPUT22), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g068(.A(G211gat), .B(G218gat), .Z(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n270), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n265), .A2(new_n272), .A3(new_n268), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(G226gat), .A2(G233gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n204), .A2(new_n276), .A3(KEYINPUT23), .ZN(new_n277));
  NAND2_X1  g076(.A1(G169gat), .A2(G176gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT67), .ZN(new_n280));
  NOR2_X1   g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n280), .B1(new_n281), .B2(KEYINPUT23), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n204), .A2(new_n276), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT23), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n283), .A2(KEYINPUT67), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n279), .B1(new_n282), .B2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G183gat), .A2(G190gat), .ZN(new_n288));
  AND2_X1   g087(.A1(KEYINPUT24), .A2(G183gat), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n292));
  OAI21_X1  g091(.A(KEYINPUT25), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NOR2_X1   g092(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  INV_X1    g095(.A(G183gat), .ZN(new_n297));
  INV_X1    g096(.A(G190gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n300), .C1(new_n292), .C2(new_n301), .ZN(new_n302));
  AND2_X1   g101(.A1(new_n292), .A2(new_n301), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n296), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(G183gat), .A2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT24), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n301), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n290), .A2(new_n308), .A3(KEYINPUT66), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n304), .A2(new_n286), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g110(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n311), .A2(KEYINPUT68), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g112(.A(KEYINPUT68), .B1(new_n311), .B2(new_n312), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n295), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g114(.A(KEYINPUT27), .B(G183gat), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n316), .A2(new_n298), .ZN(new_n317));
  OR2_X1    g116(.A1(new_n317), .A2(KEYINPUT28), .ZN(new_n318));
  AOI22_X1  g117(.A1(new_n317), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n319));
  OR2_X1    g118(.A1(new_n283), .A2(KEYINPUT26), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n283), .A2(KEYINPUT26), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n320), .A2(new_n278), .A3(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n319), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n275), .B1(new_n315), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT29), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n311), .A2(new_n312), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT68), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n311), .A2(KEYINPUT68), .A3(new_n312), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n294), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n323), .B1(new_n330), .B2(KEYINPUT69), .ZN(new_n331));
  OAI211_X1 g130(.A(KEYINPUT69), .B(new_n295), .C1(new_n313), .C2(new_n314), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  XOR2_X1   g133(.A(new_n275), .B(KEYINPUT79), .Z(new_n335));
  INV_X1    g134(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT80), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n324), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n334), .A2(KEYINPUT80), .A3(new_n336), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n274), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT69), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n315), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n343), .A2(new_n332), .A3(new_n323), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n335), .ZN(new_n345));
  INV_X1    g144(.A(new_n323), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n325), .B1(new_n330), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(new_n275), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n345), .A2(new_n274), .A3(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n262), .B1(new_n341), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n346), .B1(new_n315), .B2(new_n342), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n352), .B2(new_n332), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n338), .B1(new_n353), .B2(new_n335), .ZN(new_n354));
  INV_X1    g153(.A(new_n324), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n354), .A2(new_n340), .A3(new_n274), .A4(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n345), .A2(new_n348), .ZN(new_n357));
  INV_X1    g156(.A(new_n274), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n262), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n261), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n354), .A2(new_n340), .A3(new_n355), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n350), .B1(new_n362), .B2(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(new_n257), .ZN(new_n364));
  XNOR2_X1  g163(.A(G1gat), .B(G29gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n365), .B(KEYINPUT0), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(G57gat), .ZN(new_n367));
  INV_X1    g166(.A(G85gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(G141gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(G148gat), .ZN(new_n372));
  INV_X1    g171(.A(G148gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G141gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G155gat), .A2(G162gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n376), .A2(KEYINPUT2), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g177(.A(G155gat), .B(G162gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  OAI21_X1  g179(.A(KEYINPUT82), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n372), .A2(new_n374), .B1(KEYINPUT2), .B2(new_n376), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT82), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n382), .A2(new_n383), .A3(new_n379), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n378), .A2(new_n386), .A3(new_n380), .ZN(new_n387));
  OAI21_X1  g186(.A(KEYINPUT81), .B1(new_n382), .B2(new_n379), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n385), .A2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G113gat), .B(G120gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(KEYINPUT71), .ZN(new_n392));
  NOR2_X1   g191(.A1(G127gat), .A2(G134gat), .ZN(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(G127gat), .A2(G134gat), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT1), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n391), .A2(KEYINPUT1), .ZN(new_n397));
  NOR2_X1   g196(.A1(new_n397), .A2(new_n393), .ZN(new_n398));
  XOR2_X1   g197(.A(KEYINPUT70), .B(G127gat), .Z(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(G134gat), .ZN(new_n400));
  AOI22_X1  g199(.A1(new_n392), .A2(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n390), .B(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(G225gat), .A2(G233gat), .ZN(new_n403));
  OAI21_X1  g202(.A(KEYINPUT5), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n390), .A2(KEYINPUT83), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n385), .A2(new_n389), .A3(new_n406), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n401), .A4(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n390), .A2(KEYINPUT3), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT3), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n385), .A2(new_n389), .A3(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n392), .A2(new_n396), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n398), .A2(new_n400), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n409), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT4), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n416), .B1(new_n414), .B2(new_n390), .ZN(new_n417));
  NAND4_X1  g216(.A1(new_n408), .A2(new_n415), .A3(new_n403), .A4(new_n417), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT84), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n403), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n401), .B1(new_n390), .B2(KEYINPUT3), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n421), .B1(new_n422), .B2(new_n411), .ZN(new_n423));
  NAND4_X1  g222(.A1(new_n423), .A2(KEYINPUT84), .A3(new_n417), .A4(new_n408), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n404), .B1(new_n420), .B2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT4), .B1(new_n414), .B2(new_n390), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n405), .A2(new_n401), .A3(new_n407), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(new_n427), .B2(KEYINPUT4), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT5), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n428), .A2(new_n429), .A3(new_n423), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n370), .B1(new_n425), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n431), .A2(KEYINPUT87), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT6), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n420), .A2(new_n424), .ZN(new_n434));
  INV_X1    g233(.A(new_n404), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n436), .A2(new_n369), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT87), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n438), .B(new_n370), .C1(new_n425), .C2(new_n430), .ZN(new_n439));
  NAND4_X1  g238(.A1(new_n432), .A2(new_n433), .A3(new_n437), .A4(new_n439), .ZN(new_n440));
  OR2_X1    g239(.A1(new_n431), .A2(new_n433), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n364), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT89), .B1(new_n361), .B2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n364), .A2(new_n441), .A3(new_n440), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n363), .A2(KEYINPUT37), .ZN(new_n445));
  INV_X1    g244(.A(new_n360), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n260), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT89), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n444), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n257), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n341), .A2(new_n262), .A3(new_n350), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n450), .B1(new_n451), .B2(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n259), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n443), .A2(new_n449), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n274), .B1(new_n325), .B2(new_n411), .ZN(new_n455));
  NAND2_X1  g254(.A1(G228gat), .A2(G233gat), .ZN(new_n456));
  NOR2_X1   g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(new_n390), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT29), .B1(new_n271), .B2(new_n273), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n458), .B2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n460), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n405), .A2(new_n407), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n455), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(new_n456), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n461), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT85), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g267(.A(G78gat), .B(G106gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n469), .B(KEYINPUT31), .ZN(new_n470));
  XOR2_X1   g269(.A(new_n470), .B(G50gat), .Z(new_n471));
  NAND2_X1  g270(.A1(new_n468), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(G22gat), .ZN(new_n473));
  NOR2_X1   g272(.A1(new_n466), .A2(new_n467), .ZN(new_n474));
  INV_X1    g273(.A(G22gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(new_n475), .A3(new_n471), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n473), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n475), .B1(new_n468), .B2(new_n471), .ZN(new_n478));
  INV_X1    g277(.A(new_n471), .ZN(new_n479));
  AOI211_X1 g278(.A(G22gat), .B(new_n479), .C1(new_n466), .C2(new_n467), .ZN(new_n480));
  OAI22_X1  g279(.A1(new_n478), .A2(new_n480), .B1(new_n467), .B2(new_n466), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT30), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n364), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n450), .B1(new_n341), .B2(new_n350), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n362), .A2(new_n358), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n486), .A2(KEYINPUT30), .A3(new_n349), .A4(new_n257), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n484), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n403), .B1(new_n428), .B2(new_n415), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT39), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  AND2_X1   g290(.A1(new_n402), .A2(new_n403), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n492), .B2(KEYINPUT86), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n493), .B1(KEYINPUT86), .B2(new_n492), .ZN(new_n494));
  OAI211_X1 g293(.A(new_n491), .B(new_n369), .C1(new_n494), .C2(new_n489), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT40), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n496), .ZN(new_n498));
  AND4_X1   g297(.A1(new_n432), .A2(new_n497), .A3(new_n439), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n482), .B1(new_n488), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n454), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT36), .ZN(new_n502));
  XNOR2_X1  g301(.A(G15gat), .B(G43gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(G71gat), .B(G99gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n503), .B(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G227gat), .A2(G233gat), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n352), .A2(new_n401), .A3(new_n332), .ZN(new_n508));
  AOI21_X1  g307(.A(new_n401), .B1(new_n352), .B2(new_n332), .ZN(new_n509));
  OAI21_X1  g308(.A(new_n508), .B1(new_n509), .B2(KEYINPUT72), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT72), .ZN(new_n511));
  AOI211_X1 g310(.A(new_n511), .B(new_n401), .C1(new_n352), .C2(new_n332), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n507), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(new_n505), .B1(new_n513), .B2(KEYINPUT32), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT33), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT32), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n344), .A2(new_n414), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(new_n511), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n509), .A2(KEYINPUT72), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n520), .A2(new_n521), .A3(new_n508), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n518), .B1(new_n522), .B2(new_n507), .ZN(new_n523));
  OR2_X1    g322(.A1(new_n505), .A2(new_n515), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT73), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND4_X1  g324(.A1(new_n513), .A2(KEYINPUT73), .A3(KEYINPUT32), .A4(new_n524), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n517), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT75), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n520), .A2(new_n521), .A3(new_n506), .A4(new_n508), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT74), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT34), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(KEYINPUT34), .B1(new_n530), .B2(new_n529), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n534), .B1(new_n535), .B2(new_n532), .ZN(new_n536));
  NOR2_X1   g335(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n513), .A2(KEYINPUT32), .A3(new_n524), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(new_n526), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n530), .A2(new_n529), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(new_n533), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n530), .A2(new_n531), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n544), .A2(KEYINPUT75), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  AOI22_X1  g345(.A1(new_n541), .A2(new_n517), .B1(new_n546), .B2(new_n534), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n502), .B1(new_n537), .B2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n535), .A2(new_n532), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n529), .B(KEYINPUT34), .C1(new_n530), .C2(new_n531), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI22_X1  g350(.A1(new_n540), .A2(new_n526), .B1(new_n516), .B2(new_n514), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n502), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT76), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(new_n549), .B2(new_n550), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n534), .B(KEYINPUT76), .C1(new_n535), .C2(new_n532), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n555), .A2(new_n528), .A3(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n437), .A2(new_n433), .A3(new_n431), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n441), .ZN(new_n561));
  AOI211_X1 g360(.A(new_n450), .B(new_n350), .C1(new_n362), .C2(new_n358), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n561), .B1(new_n562), .B2(KEYINPUT30), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n485), .A2(new_n487), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n482), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n501), .A2(new_n559), .A3(new_n565), .ZN(new_n566));
  OAI21_X1  g365(.A(KEYINPUT90), .B1(new_n537), .B2(new_n547), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n528), .A2(new_n536), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT90), .ZN(new_n570));
  NAND3_X1  g369(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n440), .A2(new_n441), .ZN(new_n572));
  XOR2_X1   g371(.A(KEYINPUT91), .B(KEYINPUT35), .Z(new_n573));
  NAND4_X1  g372(.A1(new_n572), .A2(new_n477), .A3(new_n481), .A4(new_n573), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n574), .A2(new_n488), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n567), .A2(new_n571), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n482), .B1(new_n551), .B2(new_n552), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n563), .A2(new_n564), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n577), .A2(new_n557), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n579), .A2(KEYINPUT35), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n576), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n253), .B1(new_n566), .B2(new_n581), .ZN(new_n582));
  AND2_X1   g381(.A1(G232gat), .A2(G233gat), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n585), .A2(G85gat), .A3(G92gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT7), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(G99gat), .A2(G106gat), .ZN(new_n589));
  AOI22_X1  g388(.A1(KEYINPUT8), .A2(new_n589), .B1(new_n368), .B2(new_n256), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n585), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n588), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  XOR2_X1   g391(.A(G99gat), .B(G106gat), .Z(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n584), .B1(new_n223), .B2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(new_n241), .B2(new_n594), .ZN(new_n596));
  XNOR2_X1  g395(.A(G134gat), .B(G162gat), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n583), .A2(KEYINPUT41), .ZN(new_n599));
  XNOR2_X1  g398(.A(G190gat), .B(G218gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n598), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n598), .A2(new_n601), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT21), .ZN(new_n605));
  XNOR2_X1  g404(.A(G57gat), .B(G64gat), .ZN(new_n606));
  AOI21_X1  g405(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT100), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(G71gat), .B(G78gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n230), .B1(new_n605), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n611), .B(G183gat), .ZN(new_n612));
  XOR2_X1   g411(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n613));
  NAND2_X1  g412(.A1(G231gat), .A2(G233gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(new_n613), .B(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n612), .B(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n610), .A2(new_n605), .ZN(new_n617));
  XOR2_X1   g416(.A(G127gat), .B(G155gat), .Z(new_n618));
  XNOR2_X1  g417(.A(new_n617), .B(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(G211gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(KEYINPUT10), .ZN(new_n626));
  OR3_X1    g425(.A1(new_n594), .A2(new_n610), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n594), .B(new_n610), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n627), .B1(new_n628), .B2(KEYINPUT10), .ZN(new_n629));
  NAND2_X1  g428(.A1(G230gat), .A2(G233gat), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(KEYINPUT102), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n628), .A2(G230gat), .A3(G233gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(G120gat), .B(G148gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(G176gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(new_n264), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NOR2_X1   g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n630), .B(KEYINPUT103), .Z(new_n640));
  AND2_X1   g439(.A1(new_n629), .A2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n637), .B1(new_n641), .B2(new_n633), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n642), .ZN(new_n643));
  NOR3_X1   g442(.A1(new_n604), .A2(new_n625), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n582), .A2(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n645), .A2(new_n561), .ZN(new_n646));
  XOR2_X1   g445(.A(new_n646), .B(G1gat), .Z(G1324gat));
  INV_X1    g446(.A(new_n488), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n649), .A2(new_n224), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT105), .Z(new_n651));
  XOR2_X1   g450(.A(KEYINPUT16), .B(G8gat), .Z(new_n652));
  AOI21_X1  g451(.A(KEYINPUT104), .B1(new_n649), .B2(new_n652), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT42), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(G1325gat));
  OAI21_X1  g454(.A(G15gat), .B1(new_n645), .B2(new_n559), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n567), .A2(new_n571), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  OR2_X1    g457(.A1(new_n658), .A2(G15gat), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n656), .B1(new_n645), .B2(new_n659), .ZN(G1326gat));
  INV_X1    g459(.A(new_n482), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n645), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  INV_X1    g463(.A(new_n561), .ZN(new_n665));
  INV_X1    g464(.A(new_n604), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n624), .A2(new_n643), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g467(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n582), .A2(new_n665), .A3(new_n217), .A4(new_n669), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(KEYINPUT45), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n565), .A2(KEYINPUT106), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT106), .ZN(new_n673));
  OAI211_X1 g472(.A(new_n673), .B(new_n482), .C1(new_n563), .C2(new_n564), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n501), .A2(new_n559), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n676), .A2(new_n581), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n677), .A2(new_n604), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT44), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n566), .A2(new_n581), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n666), .A2(new_n679), .ZN(new_n681));
  AOI22_X1  g480(.A1(new_n678), .A2(new_n679), .B1(new_n680), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n682), .A2(new_n252), .A3(new_n667), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n683), .A2(new_n561), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n671), .B1(new_n684), .B2(new_n217), .ZN(G1328gat));
  OAI21_X1  g484(.A(G36gat), .B1(new_n683), .B2(new_n648), .ZN(new_n686));
  NAND4_X1  g485(.A1(new_n582), .A2(new_n216), .A3(new_n488), .A4(new_n669), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT46), .Z(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(G1329gat));
  OAI21_X1  g488(.A(G43gat), .B1(new_n683), .B2(new_n559), .ZN(new_n690));
  INV_X1    g489(.A(new_n669), .ZN(new_n691));
  NOR3_X1   g490(.A1(new_n658), .A2(G43gat), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n582), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n690), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT47), .Z(G1330gat));
  OAI21_X1  g494(.A(G50gat), .B1(new_n683), .B2(new_n661), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n691), .A2(new_n661), .A3(G50gat), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n582), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(KEYINPUT107), .ZN(new_n700));
  INV_X1    g499(.A(KEYINPUT107), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n696), .A2(new_n701), .A3(new_n698), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n700), .A2(KEYINPUT48), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(KEYINPUT48), .B1(new_n700), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(G1331gat));
  NOR2_X1   g504(.A1(new_n604), .A2(new_n625), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n253), .A2(new_n706), .A3(new_n643), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT108), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(new_n677), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(new_n665), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g511(.A1(new_n709), .A2(new_n648), .ZN(new_n713));
  NOR2_X1   g512(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n714));
  AND2_X1   g513(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n713), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n716), .B1(new_n713), .B2(new_n714), .ZN(G1333gat));
  OR3_X1    g516(.A1(new_n709), .A2(G71gat), .A3(new_n658), .ZN(new_n718));
  OAI21_X1  g517(.A(G71gat), .B1(new_n709), .B2(new_n559), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(new_n720), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g520(.A1(new_n710), .A2(new_n482), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G78gat), .ZN(G1335gat));
  AOI22_X1  g522(.A1(new_n548), .A2(new_n558), .B1(new_n672), .B2(new_n674), .ZN(new_n724));
  AOI22_X1  g523(.A1(new_n724), .A2(new_n501), .B1(new_n576), .B2(new_n580), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n679), .B1(new_n725), .B2(new_n666), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n680), .A2(new_n681), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n252), .A2(new_n624), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n643), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n726), .A2(new_n727), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(KEYINPUT109), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT109), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n726), .A2(new_n727), .A3(new_n734), .A4(new_n731), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G85gat), .B1(new_n736), .B2(new_n561), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n666), .B1(new_n676), .B2(new_n581), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n728), .B1(new_n738), .B2(KEYINPUT110), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT110), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n740), .A3(new_n666), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT51), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n742), .B1(new_n739), .B2(new_n741), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n561), .A2(G85gat), .A3(new_n730), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT111), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n737), .B1(new_n747), .B2(new_n749), .ZN(G1336gat));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n488), .A3(new_n735), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G92gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT112), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT112), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(new_n754), .A3(G92gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR3_X1   g555(.A1(new_n648), .A2(G92gat), .A3(new_n730), .ZN(new_n757));
  XNOR2_X1  g556(.A(new_n757), .B(KEYINPUT113), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT114), .B1(new_n739), .B2(new_n741), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n738), .A2(KEYINPUT110), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n740), .B1(new_n725), .B2(new_n666), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT114), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n728), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n759), .A2(new_n742), .A3(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n743), .B1(new_n764), .B2(KEYINPUT115), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n759), .A2(new_n766), .A3(new_n742), .A4(new_n763), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n758), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(KEYINPUT52), .B1(new_n756), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n757), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n770), .B1(new_n744), .B2(new_n745), .ZN(new_n771));
  OAI21_X1  g570(.A(G92gat), .B1(new_n732), .B2(new_n648), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT52), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OR3_X1    g573(.A1(new_n771), .A2(KEYINPUT116), .A3(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(KEYINPUT116), .B1(new_n771), .B2(new_n774), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n769), .A2(new_n777), .ZN(G1337gat));
  OAI21_X1  g577(.A(G99gat), .B1(new_n736), .B2(new_n559), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n746), .A2(new_n643), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n658), .A2(G99gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n779), .B1(new_n780), .B2(new_n781), .ZN(G1338gat));
  NAND3_X1  g581(.A1(new_n682), .A2(new_n482), .A3(new_n731), .ZN(new_n783));
  XOR2_X1   g582(.A(KEYINPUT117), .B(G106gat), .Z(new_n784));
  AOI21_X1  g583(.A(KEYINPUT53), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  OR2_X1    g584(.A1(new_n661), .A2(G106gat), .ZN(new_n786));
  OAI21_X1  g585(.A(new_n785), .B1(new_n780), .B2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n765), .A2(new_n767), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n786), .A2(new_n730), .ZN(new_n789));
  NAND3_X1  g588(.A1(new_n733), .A2(new_n482), .A3(new_n735), .ZN(new_n790));
  AOI22_X1  g589(.A1(new_n788), .A2(new_n789), .B1(new_n790), .B2(new_n784), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n787), .B1(new_n791), .B2(new_n792), .ZN(G1339gat));
  OAI211_X1 g592(.A(new_n632), .B(KEYINPUT54), .C1(new_n629), .C2(new_n640), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT54), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n636), .B1(new_n641), .B2(new_n795), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  OR2_X1    g596(.A1(new_n797), .A2(KEYINPUT55), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(KEYINPUT55), .ZN(new_n799));
  NAND3_X1  g598(.A1(new_n798), .A2(new_n639), .A3(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n252), .A2(new_n801), .ZN(new_n802));
  AND2_X1   g601(.A1(new_n246), .A2(new_n248), .ZN(new_n803));
  INV_X1    g602(.A(new_n207), .ZN(new_n804));
  OAI22_X1  g603(.A1(new_n242), .A2(new_n233), .B1(new_n231), .B2(new_n235), .ZN(new_n805));
  AOI22_X1  g604(.A1(new_n803), .A2(new_n208), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n643), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n604), .B1(new_n802), .B2(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n806), .A2(new_n604), .A3(new_n801), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n625), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n253), .A2(new_n706), .A3(new_n730), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  AND2_X1   g611(.A1(new_n577), .A2(new_n557), .ZN(new_n813));
  AND3_X1   g612(.A1(new_n812), .A2(new_n665), .A3(new_n813), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n648), .ZN(new_n815));
  AOI21_X1  g614(.A(G113gat), .B1(new_n815), .B2(new_n252), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n810), .A2(new_n811), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n817), .A2(new_n482), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n488), .A2(new_n561), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n818), .A2(new_n657), .A3(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(G113gat), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n820), .A2(new_n821), .A3(new_n253), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n816), .A2(new_n822), .ZN(G1340gat));
  AOI21_X1  g622(.A(G120gat), .B1(new_n815), .B2(new_n643), .ZN(new_n824));
  INV_X1    g623(.A(G120gat), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n820), .A2(new_n825), .A3(new_n730), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n824), .A2(new_n826), .ZN(G1341gat));
  OAI21_X1  g626(.A(new_n399), .B1(new_n820), .B2(new_n625), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n625), .A2(new_n399), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n815), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n828), .A2(new_n830), .ZN(G1342gat));
  NOR3_X1   g630(.A1(new_n666), .A2(new_n488), .A3(G134gat), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n814), .A2(new_n832), .ZN(new_n833));
  XOR2_X1   g632(.A(new_n833), .B(KEYINPUT56), .Z(new_n834));
  OAI21_X1  g633(.A(G134gat), .B1(new_n820), .B2(new_n666), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(G1343gat));
  AND4_X1   g635(.A1(new_n665), .A2(new_n812), .A3(new_n482), .A4(new_n559), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n837), .A2(new_n371), .A3(new_n252), .A4(new_n648), .ZN(new_n838));
  OR2_X1    g637(.A1(new_n800), .A2(KEYINPUT118), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n800), .A2(KEYINPUT118), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(new_n252), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n604), .B1(new_n841), .B2(new_n807), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n625), .B1(new_n842), .B2(new_n809), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n843), .A2(new_n811), .ZN(new_n844));
  OAI21_X1  g643(.A(KEYINPUT57), .B1(new_n844), .B2(new_n661), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n812), .A2(new_n482), .ZN(new_n846));
  OR2_X1    g645(.A1(new_n846), .A2(KEYINPUT57), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n559), .A2(new_n819), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n845), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(new_n253), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n838), .B1(new_n850), .B2(new_n371), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(KEYINPUT58), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n853), .B(new_n838), .C1(new_n850), .C2(new_n371), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n852), .A2(new_n854), .ZN(G1344gat));
  NOR2_X1   g654(.A1(new_n849), .A2(new_n730), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n856), .A2(KEYINPUT59), .A3(new_n373), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT59), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n811), .B(KEYINPUT119), .Z(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(new_n843), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n661), .A2(KEYINPUT57), .ZN(new_n861));
  AOI22_X1  g660(.A1(new_n860), .A2(new_n861), .B1(new_n846), .B2(KEYINPUT57), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n862), .A2(new_n643), .A3(new_n848), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n858), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n648), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n643), .A2(new_n373), .ZN(new_n866));
  OAI22_X1  g665(.A1(new_n857), .A2(new_n864), .B1(new_n865), .B2(new_n866), .ZN(G1345gat));
  OAI21_X1  g666(.A(G155gat), .B1(new_n849), .B2(new_n625), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n625), .A2(G155gat), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n868), .B1(new_n865), .B2(new_n869), .ZN(G1346gat));
  NOR3_X1   g669(.A1(new_n666), .A2(new_n488), .A3(G162gat), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n837), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT120), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n873), .B1(new_n849), .B2(new_n666), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n874), .A2(G162gat), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n849), .A2(new_n873), .A3(new_n666), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n872), .B1(new_n875), .B2(new_n876), .ZN(G1347gat));
  NOR2_X1   g676(.A1(new_n648), .A2(new_n665), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n657), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n879), .A2(KEYINPUT121), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(KEYINPUT121), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n818), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g681(.A(G169gat), .B1(new_n882), .B2(new_n253), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(KEYINPUT122), .ZN(new_n884));
  AND2_X1   g683(.A1(new_n812), .A2(new_n878), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n885), .A2(new_n813), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n204), .A3(new_n252), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n884), .A2(new_n888), .ZN(G1348gat));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n276), .A3(new_n643), .ZN(new_n890));
  OAI21_X1  g689(.A(G176gat), .B1(new_n882), .B2(new_n730), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1349gat));
  INV_X1    g691(.A(KEYINPUT60), .ZN(new_n893));
  OAI21_X1  g692(.A(G183gat), .B1(new_n882), .B2(new_n625), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT123), .ZN(new_n895));
  NAND4_X1  g694(.A1(new_n885), .A2(new_n316), .A3(new_n813), .A4(new_n624), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n895), .B1(new_n894), .B2(new_n896), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n893), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n894), .A2(new_n896), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT123), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n894), .A2(new_n895), .A3(new_n896), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n901), .A2(KEYINPUT60), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n899), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n887), .A2(new_n298), .A3(new_n604), .ZN(new_n905));
  XNOR2_X1  g704(.A(new_n905), .B(KEYINPUT124), .ZN(new_n906));
  OAI21_X1  g705(.A(G190gat), .B1(new_n882), .B2(new_n666), .ZN(new_n907));
  NOR2_X1   g706(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n908));
  AND2_X1   g707(.A1(KEYINPUT125), .A2(KEYINPUT61), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n907), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n907), .A2(new_n908), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n906), .A2(new_n910), .A3(new_n911), .ZN(G1351gat));
  AND2_X1   g711(.A1(new_n559), .A2(new_n878), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT126), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n862), .A2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(G197gat), .B1(new_n915), .B2(new_n253), .ZN(new_n916));
  INV_X1    g715(.A(new_n846), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(new_n913), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n919), .A2(new_n206), .A3(new_n252), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n916), .A2(new_n920), .ZN(G1352gat));
  NOR3_X1   g720(.A1(new_n918), .A2(G204gat), .A3(new_n730), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT62), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n862), .A2(new_n643), .A3(new_n914), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n264), .B2(new_n924), .ZN(G1353gat));
  NAND3_X1  g724(.A1(new_n919), .A2(new_n620), .A3(new_n624), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n862), .A2(new_n624), .A3(new_n914), .ZN(new_n927));
  AND3_X1   g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT63), .B1(new_n927), .B2(G211gat), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n926), .B1(new_n928), .B2(new_n929), .ZN(G1354gat));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n915), .A2(new_n666), .ZN(new_n932));
  INV_X1    g731(.A(G218gat), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n604), .A2(new_n933), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n918), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n931), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  OAI221_X1 g736(.A(KEYINPUT127), .B1(new_n918), .B2(new_n935), .C1(new_n932), .C2(new_n933), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1355gat));
endmodule


