

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U562 ( .A1(n702), .A2(n807), .ZN(n744) );
  OR2_X1 U563 ( .A1(n774), .A2(n772), .ZN(n761) );
  NOR2_X1 U564 ( .A1(n988), .A2(n707), .ZN(n712) );
  INV_X1 U565 ( .A(n744), .ZN(n728) );
  XNOR2_X1 U566 ( .A(n559), .B(KEYINPUT66), .ZN(n560) );
  XNOR2_X1 U567 ( .A(G2104), .B(KEYINPUT65), .ZN(n562) );
  XNOR2_X1 U568 ( .A(n561), .B(n560), .ZN(n564) );
  NOR2_X1 U569 ( .A1(n650), .A2(G651), .ZN(n661) );
  NOR2_X2 U570 ( .A1(n562), .A2(G2105), .ZN(n897) );
  NOR2_X1 U571 ( .A1(n566), .A2(n565), .ZN(n567) );
  INV_X1 U572 ( .A(G651), .ZN(n532) );
  NOR2_X1 U573 ( .A1(G543), .A2(n532), .ZN(n529) );
  XOR2_X1 U574 ( .A(KEYINPUT1), .B(n529), .Z(n656) );
  NAND2_X1 U575 ( .A1(G64), .A2(n656), .ZN(n531) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n650) );
  NAND2_X1 U577 ( .A1(G52), .A2(n661), .ZN(n530) );
  NAND2_X1 U578 ( .A1(n531), .A2(n530), .ZN(n538) );
  NOR2_X1 U579 ( .A1(n650), .A2(n532), .ZN(n660) );
  NAND2_X1 U580 ( .A1(n660), .A2(G77), .ZN(n533) );
  XOR2_X1 U581 ( .A(KEYINPUT67), .B(n533), .Z(n535) );
  NOR2_X1 U582 ( .A1(G543), .A2(G651), .ZN(n657) );
  NAND2_X1 U583 ( .A1(n657), .A2(G90), .ZN(n534) );
  NAND2_X1 U584 ( .A1(n535), .A2(n534), .ZN(n536) );
  XOR2_X1 U585 ( .A(KEYINPUT9), .B(n536), .Z(n537) );
  NOR2_X1 U586 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U587 ( .A(KEYINPUT68), .B(n539), .ZN(G171) );
  INV_X1 U588 ( .A(G171), .ZN(G301) );
  NAND2_X1 U589 ( .A1(G85), .A2(n657), .ZN(n541) );
  NAND2_X1 U590 ( .A1(G72), .A2(n660), .ZN(n540) );
  NAND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U592 ( .A1(G60), .A2(n656), .ZN(n543) );
  NAND2_X1 U593 ( .A1(G47), .A2(n661), .ZN(n542) );
  NAND2_X1 U594 ( .A1(n543), .A2(n542), .ZN(n544) );
  OR2_X1 U595 ( .A1(n545), .A2(n544), .ZN(G290) );
  XOR2_X1 U596 ( .A(G2435), .B(G2454), .Z(n547) );
  XNOR2_X1 U597 ( .A(G2430), .B(G2438), .ZN(n546) );
  XNOR2_X1 U598 ( .A(n547), .B(n546), .ZN(n554) );
  XOR2_X1 U599 ( .A(G2446), .B(KEYINPUT111), .Z(n549) );
  XNOR2_X1 U600 ( .A(G2451), .B(G2443), .ZN(n548) );
  XNOR2_X1 U601 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U602 ( .A(n550), .B(G2427), .Z(n552) );
  XNOR2_X1 U603 ( .A(G1348), .B(G1341), .ZN(n551) );
  XNOR2_X1 U604 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U605 ( .A(n554), .B(n553), .ZN(n555) );
  AND2_X1 U606 ( .A1(n555), .A2(G14), .ZN(G401) );
  AND2_X1 U607 ( .A1(G2105), .A2(G2104), .ZN(n901) );
  NAND2_X1 U608 ( .A1(G113), .A2(n901), .ZN(n558) );
  NOR2_X1 U609 ( .A1(G2105), .A2(G2104), .ZN(n556) );
  XOR2_X1 U610 ( .A(KEYINPUT17), .B(n556), .Z(n898) );
  NAND2_X1 U611 ( .A1(G137), .A2(n898), .ZN(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n566) );
  NAND2_X1 U613 ( .A1(G101), .A2(n897), .ZN(n561) );
  INV_X1 U614 ( .A(KEYINPUT23), .ZN(n559) );
  AND2_X1 U615 ( .A1(n562), .A2(G2105), .ZN(n902) );
  NAND2_X1 U616 ( .A1(G125), .A2(n902), .ZN(n563) );
  NAND2_X1 U617 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U618 ( .A(KEYINPUT64), .B(n567), .ZN(n701) );
  BUF_X1 U619 ( .A(n701), .Z(G160) );
  AND2_X1 U620 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U621 ( .A(G132), .ZN(G219) );
  INV_X1 U622 ( .A(G82), .ZN(G220) );
  NAND2_X1 U623 ( .A1(n656), .A2(G62), .ZN(n570) );
  NAND2_X1 U624 ( .A1(G50), .A2(n661), .ZN(n568) );
  XOR2_X1 U625 ( .A(KEYINPUT87), .B(n568), .Z(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U627 ( .A1(G88), .A2(n657), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G75), .A2(n660), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U630 ( .A1(n574), .A2(n573), .ZN(G166) );
  NAND2_X1 U631 ( .A1(n657), .A2(G89), .ZN(n575) );
  XNOR2_X1 U632 ( .A(n575), .B(KEYINPUT4), .ZN(n577) );
  NAND2_X1 U633 ( .A1(G76), .A2(n660), .ZN(n576) );
  NAND2_X1 U634 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U635 ( .A(n578), .B(KEYINPUT5), .ZN(n583) );
  NAND2_X1 U636 ( .A1(G63), .A2(n656), .ZN(n580) );
  NAND2_X1 U637 ( .A1(G51), .A2(n661), .ZN(n579) );
  NAND2_X1 U638 ( .A1(n580), .A2(n579), .ZN(n581) );
  XOR2_X1 U639 ( .A(KEYINPUT6), .B(n581), .Z(n582) );
  NAND2_X1 U640 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U641 ( .A(n584), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U642 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U643 ( .A1(G7), .A2(G661), .ZN(n585) );
  XNOR2_X1 U644 ( .A(n585), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U645 ( .A(G223), .ZN(n843) );
  NAND2_X1 U646 ( .A1(n843), .A2(G567), .ZN(n586) );
  XNOR2_X1 U647 ( .A(n586), .B(KEYINPUT11), .ZN(n587) );
  XNOR2_X1 U648 ( .A(KEYINPUT71), .B(n587), .ZN(G234) );
  XOR2_X1 U649 ( .A(G860), .B(KEYINPUT74), .Z(n620) );
  XOR2_X1 U650 ( .A(KEYINPUT14), .B(KEYINPUT72), .Z(n589) );
  NAND2_X1 U651 ( .A1(G56), .A2(n656), .ZN(n588) );
  XNOR2_X1 U652 ( .A(n589), .B(n588), .ZN(n596) );
  NAND2_X1 U653 ( .A1(G81), .A2(n657), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT73), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(n591), .B(KEYINPUT12), .ZN(n593) );
  NAND2_X1 U656 ( .A1(G68), .A2(n660), .ZN(n592) );
  NAND2_X1 U657 ( .A1(n593), .A2(n592), .ZN(n594) );
  XOR2_X1 U658 ( .A(KEYINPUT13), .B(n594), .Z(n595) );
  NOR2_X1 U659 ( .A1(n596), .A2(n595), .ZN(n598) );
  NAND2_X1 U660 ( .A1(n661), .A2(G43), .ZN(n597) );
  NAND2_X1 U661 ( .A1(n598), .A2(n597), .ZN(n988) );
  OR2_X1 U662 ( .A1(n620), .A2(n988), .ZN(G153) );
  NAND2_X1 U663 ( .A1(G301), .A2(G868), .ZN(n609) );
  NAND2_X1 U664 ( .A1(n657), .A2(G92), .ZN(n599) );
  XOR2_X1 U665 ( .A(KEYINPUT75), .B(n599), .Z(n601) );
  NAND2_X1 U666 ( .A1(n656), .A2(G66), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n602) );
  XNOR2_X1 U668 ( .A(KEYINPUT76), .B(n602), .ZN(n606) );
  NAND2_X1 U669 ( .A1(G79), .A2(n660), .ZN(n604) );
  NAND2_X1 U670 ( .A1(G54), .A2(n661), .ZN(n603) );
  NAND2_X1 U671 ( .A1(n604), .A2(n603), .ZN(n605) );
  NOR2_X1 U672 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U673 ( .A(KEYINPUT15), .B(n607), .Z(n972) );
  OR2_X1 U674 ( .A1(n972), .A2(G868), .ZN(n608) );
  NAND2_X1 U675 ( .A1(n609), .A2(n608), .ZN(G284) );
  NAND2_X1 U676 ( .A1(G65), .A2(n656), .ZN(n611) );
  NAND2_X1 U677 ( .A1(G91), .A2(n657), .ZN(n610) );
  NAND2_X1 U678 ( .A1(n611), .A2(n610), .ZN(n614) );
  NAND2_X1 U679 ( .A1(G53), .A2(n661), .ZN(n612) );
  XNOR2_X1 U680 ( .A(KEYINPUT69), .B(n612), .ZN(n613) );
  NOR2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U682 ( .A1(n660), .A2(G78), .ZN(n615) );
  NAND2_X1 U683 ( .A1(n616), .A2(n615), .ZN(G299) );
  INV_X1 U684 ( .A(G299), .ZN(n973) );
  INV_X1 U685 ( .A(G868), .ZN(n672) );
  NAND2_X1 U686 ( .A1(n973), .A2(n672), .ZN(n617) );
  XNOR2_X1 U687 ( .A(n617), .B(KEYINPUT77), .ZN(n619) );
  NOR2_X1 U688 ( .A1(n672), .A2(G286), .ZN(n618) );
  NOR2_X1 U689 ( .A1(n619), .A2(n618), .ZN(G297) );
  NAND2_X1 U690 ( .A1(n620), .A2(G559), .ZN(n621) );
  NAND2_X1 U691 ( .A1(n621), .A2(n972), .ZN(n622) );
  XNOR2_X1 U692 ( .A(n622), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U693 ( .A1(G868), .A2(n988), .ZN(n625) );
  NAND2_X1 U694 ( .A1(G868), .A2(n972), .ZN(n623) );
  NOR2_X1 U695 ( .A1(G559), .A2(n623), .ZN(n624) );
  NOR2_X1 U696 ( .A1(n625), .A2(n624), .ZN(G282) );
  NAND2_X1 U697 ( .A1(G111), .A2(n901), .ZN(n627) );
  NAND2_X1 U698 ( .A1(G99), .A2(n897), .ZN(n626) );
  NAND2_X1 U699 ( .A1(n627), .A2(n626), .ZN(n628) );
  XNOR2_X1 U700 ( .A(KEYINPUT79), .B(n628), .ZN(n634) );
  NAND2_X1 U701 ( .A1(n902), .A2(G123), .ZN(n629) );
  XNOR2_X1 U702 ( .A(n629), .B(KEYINPUT18), .ZN(n631) );
  NAND2_X1 U703 ( .A1(G135), .A2(n898), .ZN(n630) );
  NAND2_X1 U704 ( .A1(n631), .A2(n630), .ZN(n632) );
  XOR2_X1 U705 ( .A(KEYINPUT78), .B(n632), .Z(n633) );
  NAND2_X1 U706 ( .A1(n634), .A2(n633), .ZN(n933) );
  XNOR2_X1 U707 ( .A(G2096), .B(n933), .ZN(n635) );
  NOR2_X1 U708 ( .A1(G2100), .A2(n635), .ZN(n636) );
  XOR2_X1 U709 ( .A(KEYINPUT80), .B(n636), .Z(G156) );
  NAND2_X1 U710 ( .A1(G86), .A2(n657), .ZN(n645) );
  NAND2_X1 U711 ( .A1(G73), .A2(n660), .ZN(n637) );
  XNOR2_X1 U712 ( .A(n637), .B(KEYINPUT84), .ZN(n638) );
  XNOR2_X1 U713 ( .A(n638), .B(KEYINPUT2), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G61), .A2(n656), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G48), .A2(n661), .ZN(n641) );
  XNOR2_X1 U717 ( .A(KEYINPUT85), .B(n641), .ZN(n642) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U719 ( .A1(n645), .A2(n644), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT86), .ZN(G305) );
  NAND2_X1 U721 ( .A1(G49), .A2(n661), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U724 ( .A1(n656), .A2(n649), .ZN(n653) );
  NAND2_X1 U725 ( .A1(G87), .A2(n650), .ZN(n651) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(n651), .Z(n652) );
  NAND2_X1 U727 ( .A1(n653), .A2(n652), .ZN(G288) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(G288), .ZN(n654) );
  XNOR2_X1 U729 ( .A(n654), .B(n988), .ZN(n655) );
  XNOR2_X1 U730 ( .A(G305), .B(n655), .ZN(n670) );
  NAND2_X1 U731 ( .A1(G67), .A2(n656), .ZN(n659) );
  NAND2_X1 U732 ( .A1(G93), .A2(n657), .ZN(n658) );
  NAND2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n665) );
  NAND2_X1 U734 ( .A1(G80), .A2(n660), .ZN(n663) );
  NAND2_X1 U735 ( .A1(G55), .A2(n661), .ZN(n662) );
  NAND2_X1 U736 ( .A1(n663), .A2(n662), .ZN(n664) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  XOR2_X1 U738 ( .A(KEYINPUT82), .B(n666), .Z(n851) );
  XNOR2_X1 U739 ( .A(n973), .B(n851), .ZN(n668) );
  XNOR2_X1 U740 ( .A(G290), .B(G166), .ZN(n667) );
  XNOR2_X1 U741 ( .A(n668), .B(n667), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n670), .B(n669), .ZN(n914) );
  NAND2_X1 U743 ( .A1(n972), .A2(G559), .ZN(n848) );
  XOR2_X1 U744 ( .A(n914), .B(n848), .Z(n671) );
  NAND2_X1 U745 ( .A1(G868), .A2(n671), .ZN(n674) );
  NAND2_X1 U746 ( .A1(n851), .A2(n672), .ZN(n673) );
  NAND2_X1 U747 ( .A1(n674), .A2(n673), .ZN(G295) );
  NAND2_X1 U748 ( .A1(G2078), .A2(G2084), .ZN(n675) );
  XOR2_X1 U749 ( .A(KEYINPUT20), .B(n675), .Z(n676) );
  NAND2_X1 U750 ( .A1(G2090), .A2(n676), .ZN(n677) );
  XNOR2_X1 U751 ( .A(KEYINPUT21), .B(n677), .ZN(n678) );
  NAND2_X1 U752 ( .A1(n678), .A2(G2072), .ZN(G158) );
  XOR2_X1 U753 ( .A(KEYINPUT70), .B(G57), .Z(G237) );
  XNOR2_X1 U754 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U755 ( .A1(G120), .A2(G69), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT89), .B(n679), .Z(n680) );
  NOR2_X1 U757 ( .A1(G237), .A2(n680), .ZN(n681) );
  XNOR2_X1 U758 ( .A(KEYINPUT90), .B(n681), .ZN(n682) );
  NAND2_X1 U759 ( .A1(n682), .A2(G108), .ZN(n853) );
  NAND2_X1 U760 ( .A1(G567), .A2(n853), .ZN(n683) );
  XNOR2_X1 U761 ( .A(n683), .B(KEYINPUT91), .ZN(n689) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n684) );
  XNOR2_X1 U763 ( .A(KEYINPUT22), .B(n684), .ZN(n685) );
  NAND2_X1 U764 ( .A1(n685), .A2(G96), .ZN(n686) );
  NOR2_X1 U765 ( .A1(n686), .A2(G218), .ZN(n687) );
  XOR2_X1 U766 ( .A(n687), .B(KEYINPUT88), .Z(n852) );
  AND2_X1 U767 ( .A1(n852), .A2(G2106), .ZN(n688) );
  NOR2_X1 U768 ( .A1(n689), .A2(n688), .ZN(G319) );
  INV_X1 U769 ( .A(G319), .ZN(n692) );
  NAND2_X1 U770 ( .A1(G661), .A2(G483), .ZN(n690) );
  XNOR2_X1 U771 ( .A(KEYINPUT92), .B(n690), .ZN(n691) );
  NOR2_X1 U772 ( .A1(n692), .A2(n691), .ZN(n846) );
  NAND2_X1 U773 ( .A1(n846), .A2(G36), .ZN(G176) );
  NAND2_X1 U774 ( .A1(G114), .A2(n901), .ZN(n693) );
  XNOR2_X1 U775 ( .A(n693), .B(KEYINPUT94), .ZN(n696) );
  NAND2_X1 U776 ( .A1(G126), .A2(n902), .ZN(n694) );
  XOR2_X1 U777 ( .A(KEYINPUT93), .B(n694), .Z(n695) );
  NAND2_X1 U778 ( .A1(n696), .A2(n695), .ZN(n700) );
  NAND2_X1 U779 ( .A1(n898), .A2(G138), .ZN(n698) );
  NAND2_X1 U780 ( .A1(n897), .A2(G102), .ZN(n697) );
  NAND2_X1 U781 ( .A1(n698), .A2(n697), .ZN(n699) );
  NOR2_X1 U782 ( .A1(n700), .A2(n699), .ZN(G164) );
  INV_X1 U783 ( .A(G166), .ZN(G303) );
  XNOR2_X1 U784 ( .A(KEYINPUT29), .B(KEYINPUT105), .ZN(n726) );
  NAND2_X1 U785 ( .A1(G40), .A2(n701), .ZN(n806) );
  INV_X1 U786 ( .A(n806), .ZN(n702) );
  NOR2_X1 U787 ( .A1(G164), .A2(G1384), .ZN(n807) );
  NAND2_X1 U788 ( .A1(G1996), .A2(n728), .ZN(n703) );
  XNOR2_X1 U789 ( .A(n703), .B(KEYINPUT26), .ZN(n705) );
  NAND2_X1 U790 ( .A1(G1341), .A2(n744), .ZN(n704) );
  NAND2_X1 U791 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U792 ( .A(KEYINPUT104), .B(n706), .ZN(n707) );
  NAND2_X1 U793 ( .A1(n972), .A2(n712), .ZN(n711) );
  NOR2_X1 U794 ( .A1(n728), .A2(G1348), .ZN(n709) );
  NOR2_X1 U795 ( .A1(G2067), .A2(n744), .ZN(n708) );
  NOR2_X1 U796 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U797 ( .A1(n711), .A2(n710), .ZN(n714) );
  OR2_X1 U798 ( .A1(n972), .A2(n712), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n719) );
  NAND2_X1 U800 ( .A1(n728), .A2(G2072), .ZN(n715) );
  XNOR2_X1 U801 ( .A(n715), .B(KEYINPUT27), .ZN(n717) );
  INV_X1 U802 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U803 ( .A1(n999), .A2(n728), .ZN(n716) );
  NOR2_X1 U804 ( .A1(n717), .A2(n716), .ZN(n720) );
  NAND2_X1 U805 ( .A1(n973), .A2(n720), .ZN(n718) );
  NAND2_X1 U806 ( .A1(n719), .A2(n718), .ZN(n724) );
  NOR2_X1 U807 ( .A1(n973), .A2(n720), .ZN(n722) );
  XNOR2_X1 U808 ( .A(KEYINPUT103), .B(KEYINPUT28), .ZN(n721) );
  XNOR2_X1 U809 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U810 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U811 ( .A(n726), .B(n725), .ZN(n733) );
  XOR2_X1 U812 ( .A(G2078), .B(KEYINPUT25), .Z(n957) );
  NOR2_X1 U813 ( .A1(n957), .A2(n744), .ZN(n727) );
  XOR2_X1 U814 ( .A(KEYINPUT102), .B(n727), .Z(n731) );
  NOR2_X1 U815 ( .A1(n728), .A2(G1961), .ZN(n729) );
  XNOR2_X1 U816 ( .A(KEYINPUT101), .B(n729), .ZN(n730) );
  NAND2_X1 U817 ( .A1(n731), .A2(n730), .ZN(n738) );
  NAND2_X1 U818 ( .A1(n738), .A2(G171), .ZN(n732) );
  NAND2_X1 U819 ( .A1(n733), .A2(n732), .ZN(n743) );
  NAND2_X1 U820 ( .A1(G8), .A2(n744), .ZN(n770) );
  NOR2_X1 U821 ( .A1(G1966), .A2(n770), .ZN(n758) );
  NOR2_X1 U822 ( .A1(G2084), .A2(n744), .ZN(n754) );
  NOR2_X1 U823 ( .A1(n758), .A2(n754), .ZN(n734) );
  NAND2_X1 U824 ( .A1(G8), .A2(n734), .ZN(n735) );
  XNOR2_X1 U825 ( .A(KEYINPUT30), .B(n735), .ZN(n736) );
  NOR2_X1 U826 ( .A1(G168), .A2(n736), .ZN(n737) );
  XNOR2_X1 U827 ( .A(n737), .B(KEYINPUT106), .ZN(n740) );
  NOR2_X1 U828 ( .A1(G171), .A2(n738), .ZN(n739) );
  NOR2_X1 U829 ( .A1(n740), .A2(n739), .ZN(n741) );
  XOR2_X1 U830 ( .A(KEYINPUT31), .B(n741), .Z(n742) );
  NAND2_X1 U831 ( .A1(n743), .A2(n742), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n756), .A2(G286), .ZN(n752) );
  INV_X1 U833 ( .A(G8), .ZN(n750) );
  NOR2_X1 U834 ( .A1(G1971), .A2(n770), .ZN(n746) );
  NOR2_X1 U835 ( .A1(G2090), .A2(n744), .ZN(n745) );
  NOR2_X1 U836 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U837 ( .A1(n747), .A2(G303), .ZN(n748) );
  XOR2_X1 U838 ( .A(KEYINPUT107), .B(n748), .Z(n749) );
  OR2_X1 U839 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U840 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U841 ( .A(KEYINPUT32), .B(n753), .ZN(n774) );
  NAND2_X1 U842 ( .A1(G8), .A2(n754), .ZN(n755) );
  NAND2_X1 U843 ( .A1(n756), .A2(n755), .ZN(n757) );
  NOR2_X1 U844 ( .A1(n758), .A2(n757), .ZN(n772) );
  NOR2_X1 U845 ( .A1(G2090), .A2(G303), .ZN(n759) );
  NAND2_X1 U846 ( .A1(G8), .A2(n759), .ZN(n760) );
  NAND2_X1 U847 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U848 ( .A1(n762), .A2(n770), .ZN(n764) );
  INV_X1 U849 ( .A(KEYINPUT109), .ZN(n763) );
  XNOR2_X1 U850 ( .A(n764), .B(n763), .ZN(n790) );
  NOR2_X1 U851 ( .A1(G305), .A2(G1981), .ZN(n765) );
  XOR2_X1 U852 ( .A(n765), .B(KEYINPUT24), .Z(n766) );
  NOR2_X1 U853 ( .A1(n770), .A2(n766), .ZN(n767) );
  XNOR2_X1 U854 ( .A(n767), .B(KEYINPUT100), .ZN(n788) );
  XNOR2_X1 U855 ( .A(G305), .B(G1981), .ZN(n990) );
  NAND2_X1 U856 ( .A1(G1976), .A2(G288), .ZN(n975) );
  INV_X1 U857 ( .A(KEYINPUT33), .ZN(n780) );
  OR2_X1 U858 ( .A1(G1976), .A2(G288), .ZN(n776) );
  OR2_X1 U859 ( .A1(n770), .A2(n776), .ZN(n768) );
  NOR2_X1 U860 ( .A1(n780), .A2(n768), .ZN(n769) );
  XOR2_X1 U861 ( .A(n769), .B(KEYINPUT108), .Z(n779) );
  NAND2_X1 U862 ( .A1(n975), .A2(n779), .ZN(n771) );
  OR2_X1 U863 ( .A1(n771), .A2(n770), .ZN(n775) );
  OR2_X1 U864 ( .A1(n772), .A2(n775), .ZN(n773) );
  NOR2_X1 U865 ( .A1(n774), .A2(n773), .ZN(n785) );
  INV_X1 U866 ( .A(n775), .ZN(n778) );
  INV_X1 U867 ( .A(G1971), .ZN(n1010) );
  NAND2_X1 U868 ( .A1(G166), .A2(n1010), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n777), .A2(n776), .ZN(n981) );
  AND2_X1 U870 ( .A1(n778), .A2(n981), .ZN(n783) );
  INV_X1 U871 ( .A(n779), .ZN(n781) );
  NOR2_X1 U872 ( .A1(n781), .A2(n780), .ZN(n782) );
  OR2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n784) );
  NOR2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n786) );
  NOR2_X1 U875 ( .A1(n990), .A2(n786), .ZN(n787) );
  NOR2_X1 U876 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U877 ( .A1(n790), .A2(n789), .ZN(n810) );
  NAND2_X1 U878 ( .A1(G95), .A2(n897), .ZN(n792) );
  NAND2_X1 U879 ( .A1(G131), .A2(n898), .ZN(n791) );
  NAND2_X1 U880 ( .A1(n792), .A2(n791), .ZN(n796) );
  NAND2_X1 U881 ( .A1(G107), .A2(n901), .ZN(n794) );
  NAND2_X1 U882 ( .A1(G119), .A2(n902), .ZN(n793) );
  NAND2_X1 U883 ( .A1(n794), .A2(n793), .ZN(n795) );
  NOR2_X1 U884 ( .A1(n796), .A2(n795), .ZN(n881) );
  INV_X1 U885 ( .A(G1991), .ZN(n962) );
  NOR2_X1 U886 ( .A1(n881), .A2(n962), .ZN(n805) );
  NAND2_X1 U887 ( .A1(G117), .A2(n901), .ZN(n798) );
  NAND2_X1 U888 ( .A1(G141), .A2(n898), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n801) );
  NAND2_X1 U890 ( .A1(n897), .A2(G105), .ZN(n799) );
  XOR2_X1 U891 ( .A(KEYINPUT38), .B(n799), .Z(n800) );
  NOR2_X1 U892 ( .A1(n801), .A2(n800), .ZN(n803) );
  NAND2_X1 U893 ( .A1(n902), .A2(G129), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n893) );
  AND2_X1 U895 ( .A1(G1996), .A2(n893), .ZN(n804) );
  NOR2_X1 U896 ( .A1(n805), .A2(n804), .ZN(n934) );
  NOR2_X1 U897 ( .A1(n807), .A2(n806), .ZN(n838) );
  INV_X1 U898 ( .A(n838), .ZN(n808) );
  NOR2_X1 U899 ( .A1(n934), .A2(n808), .ZN(n830) );
  INV_X1 U900 ( .A(n830), .ZN(n809) );
  NAND2_X1 U901 ( .A1(n810), .A2(n809), .ZN(n813) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n977) );
  NAND2_X1 U903 ( .A1(n838), .A2(n977), .ZN(n811) );
  XNOR2_X1 U904 ( .A(KEYINPUT95), .B(n811), .ZN(n812) );
  NOR2_X1 U905 ( .A1(n813), .A2(n812), .ZN(n827) );
  XNOR2_X1 U906 ( .A(KEYINPUT36), .B(KEYINPUT98), .ZN(n814) );
  XNOR2_X1 U907 ( .A(n814), .B(KEYINPUT97), .ZN(n825) );
  NAND2_X1 U908 ( .A1(n898), .A2(G140), .ZN(n815) );
  XNOR2_X1 U909 ( .A(n815), .B(KEYINPUT96), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G104), .A2(n897), .ZN(n816) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  XNOR2_X1 U912 ( .A(KEYINPUT34), .B(n818), .ZN(n823) );
  NAND2_X1 U913 ( .A1(G116), .A2(n901), .ZN(n820) );
  NAND2_X1 U914 ( .A1(G128), .A2(n902), .ZN(n819) );
  NAND2_X1 U915 ( .A1(n820), .A2(n819), .ZN(n821) );
  XOR2_X1 U916 ( .A(n821), .B(KEYINPUT35), .Z(n822) );
  NOR2_X1 U917 ( .A1(n823), .A2(n822), .ZN(n824) );
  XOR2_X1 U918 ( .A(n825), .B(n824), .Z(n910) );
  XNOR2_X1 U919 ( .A(G2067), .B(KEYINPUT37), .ZN(n835) );
  NOR2_X1 U920 ( .A1(n910), .A2(n835), .ZN(n940) );
  NAND2_X1 U921 ( .A1(n940), .A2(n838), .ZN(n826) );
  XOR2_X1 U922 ( .A(KEYINPUT99), .B(n826), .Z(n833) );
  NAND2_X1 U923 ( .A1(n827), .A2(n833), .ZN(n840) );
  NOR2_X1 U924 ( .A1(G1996), .A2(n893), .ZN(n931) );
  NOR2_X1 U925 ( .A1(G1986), .A2(G290), .ZN(n828) );
  AND2_X1 U926 ( .A1(n962), .A2(n881), .ZN(n936) );
  NOR2_X1 U927 ( .A1(n828), .A2(n936), .ZN(n829) );
  NOR2_X1 U928 ( .A1(n830), .A2(n829), .ZN(n831) );
  NOR2_X1 U929 ( .A1(n931), .A2(n831), .ZN(n832) );
  XNOR2_X1 U930 ( .A(KEYINPUT39), .B(n832), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n834), .A2(n833), .ZN(n836) );
  NAND2_X1 U932 ( .A1(n910), .A2(n835), .ZN(n928) );
  NAND2_X1 U933 ( .A1(n836), .A2(n928), .ZN(n837) );
  NAND2_X1 U934 ( .A1(n838), .A2(n837), .ZN(n839) );
  NAND2_X1 U935 ( .A1(n840), .A2(n839), .ZN(n842) );
  XNOR2_X1 U936 ( .A(KEYINPUT40), .B(KEYINPUT110), .ZN(n841) );
  XNOR2_X1 U937 ( .A(n842), .B(n841), .ZN(G329) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n843), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n844) );
  NAND2_X1 U940 ( .A1(G661), .A2(n844), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n845) );
  NAND2_X1 U942 ( .A1(n846), .A2(n845), .ZN(G188) );
  XOR2_X1 U943 ( .A(G69), .B(KEYINPUT112), .Z(G235) );
  XOR2_X1 U945 ( .A(KEYINPUT81), .B(n988), .Z(n847) );
  XNOR2_X1 U946 ( .A(n848), .B(n847), .ZN(n849) );
  NOR2_X1 U947 ( .A1(G860), .A2(n849), .ZN(n850) );
  XOR2_X1 U948 ( .A(n851), .B(n850), .Z(G145) );
  INV_X1 U949 ( .A(G120), .ZN(G236) );
  INV_X1 U950 ( .A(G108), .ZN(G238) );
  INV_X1 U951 ( .A(G96), .ZN(G221) );
  NOR2_X1 U952 ( .A1(n853), .A2(n852), .ZN(G325) );
  INV_X1 U953 ( .A(G325), .ZN(G261) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2084), .Z(n855) );
  XNOR2_X1 U955 ( .A(G2072), .B(G2078), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n856), .B(G2100), .Z(n858) );
  XNOR2_X1 U958 ( .A(G2067), .B(G2090), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U960 ( .A(G2096), .B(KEYINPUT43), .Z(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT113), .B(G2678), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(n862), .B(n861), .Z(G227) );
  XOR2_X1 U964 ( .A(G1961), .B(G1956), .Z(n864) );
  XNOR2_X1 U965 ( .A(G1986), .B(G1966), .ZN(n863) );
  XNOR2_X1 U966 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U967 ( .A(n865), .B(G2474), .Z(n867) );
  XNOR2_X1 U968 ( .A(G1976), .B(G1971), .ZN(n866) );
  XNOR2_X1 U969 ( .A(n867), .B(n866), .ZN(n871) );
  XOR2_X1 U970 ( .A(KEYINPUT41), .B(G1981), .Z(n869) );
  XNOR2_X1 U971 ( .A(G1996), .B(G1991), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n869), .B(n868), .ZN(n870) );
  XNOR2_X1 U973 ( .A(n871), .B(n870), .ZN(G229) );
  NAND2_X1 U974 ( .A1(G136), .A2(n898), .ZN(n872) );
  XNOR2_X1 U975 ( .A(n872), .B(KEYINPUT114), .ZN(n875) );
  NAND2_X1 U976 ( .A1(G124), .A2(n902), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n873), .B(KEYINPUT44), .ZN(n874) );
  NAND2_X1 U978 ( .A1(n875), .A2(n874), .ZN(n880) );
  NAND2_X1 U979 ( .A1(G112), .A2(n901), .ZN(n877) );
  NAND2_X1 U980 ( .A1(G100), .A2(n897), .ZN(n876) );
  NAND2_X1 U981 ( .A1(n877), .A2(n876), .ZN(n878) );
  XOR2_X1 U982 ( .A(KEYINPUT115), .B(n878), .Z(n879) );
  NOR2_X1 U983 ( .A1(n880), .A2(n879), .ZN(G162) );
  XOR2_X1 U984 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n883) );
  XNOR2_X1 U985 ( .A(n881), .B(KEYINPUT116), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n892) );
  NAND2_X1 U987 ( .A1(G118), .A2(n901), .ZN(n885) );
  NAND2_X1 U988 ( .A1(G130), .A2(n902), .ZN(n884) );
  NAND2_X1 U989 ( .A1(n885), .A2(n884), .ZN(n890) );
  NAND2_X1 U990 ( .A1(G106), .A2(n897), .ZN(n887) );
  NAND2_X1 U991 ( .A1(G142), .A2(n898), .ZN(n886) );
  NAND2_X1 U992 ( .A1(n887), .A2(n886), .ZN(n888) );
  XOR2_X1 U993 ( .A(n888), .B(KEYINPUT45), .Z(n889) );
  NOR2_X1 U994 ( .A1(n890), .A2(n889), .ZN(n891) );
  XOR2_X1 U995 ( .A(n892), .B(n891), .Z(n896) );
  XNOR2_X1 U996 ( .A(G164), .B(G160), .ZN(n894) );
  XNOR2_X1 U997 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U998 ( .A(n896), .B(n895), .Z(n909) );
  NAND2_X1 U999 ( .A1(G103), .A2(n897), .ZN(n900) );
  NAND2_X1 U1000 ( .A1(G139), .A2(n898), .ZN(n899) );
  NAND2_X1 U1001 ( .A1(n900), .A2(n899), .ZN(n907) );
  NAND2_X1 U1002 ( .A1(G115), .A2(n901), .ZN(n904) );
  NAND2_X1 U1003 ( .A1(G127), .A2(n902), .ZN(n903) );
  NAND2_X1 U1004 ( .A1(n904), .A2(n903), .ZN(n905) );
  XOR2_X1 U1005 ( .A(KEYINPUT47), .B(n905), .Z(n906) );
  NOR2_X1 U1006 ( .A1(n907), .A2(n906), .ZN(n923) );
  XNOR2_X1 U1007 ( .A(n923), .B(G162), .ZN(n908) );
  XNOR2_X1 U1008 ( .A(n909), .B(n908), .ZN(n912) );
  XOR2_X1 U1009 ( .A(n933), .B(n910), .Z(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  NOR2_X1 U1011 ( .A1(G37), .A2(n913), .ZN(G395) );
  XOR2_X1 U1012 ( .A(n914), .B(G286), .Z(n916) );
  XNOR2_X1 U1013 ( .A(n972), .B(G301), .ZN(n915) );
  XNOR2_X1 U1014 ( .A(n916), .B(n915), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G37), .A2(n917), .ZN(G397) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n918) );
  XNOR2_X1 U1017 ( .A(KEYINPUT49), .B(n918), .ZN(n919) );
  NOR2_X1 U1018 ( .A1(G401), .A2(n919), .ZN(n920) );
  AND2_X1 U1019 ( .A1(G319), .A2(n920), .ZN(n922) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n921) );
  NAND2_X1 U1021 ( .A1(n922), .A2(n921), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  XOR2_X1 U1023 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(KEYINPUT50), .B(n926), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n927), .B(KEYINPUT118), .ZN(n929) );
  NAND2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n945) );
  XOR2_X1 U1029 ( .A(G2090), .B(G162), .Z(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XOR2_X1 U1031 ( .A(KEYINPUT51), .B(n932), .Z(n942) );
  XNOR2_X1 U1032 ( .A(G2084), .B(G160), .ZN(n938) );
  NAND2_X1 U1033 ( .A1(n934), .A2(n933), .ZN(n935) );
  NOR2_X1 U1034 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1035 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  NAND2_X1 U1037 ( .A1(n942), .A2(n941), .ZN(n943) );
  XOR2_X1 U1038 ( .A(n943), .B(KEYINPUT117), .Z(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1040 ( .A(KEYINPUT119), .B(n946), .Z(n947) );
  XNOR2_X1 U1041 ( .A(KEYINPUT52), .B(n947), .ZN(n948) );
  INV_X1 U1042 ( .A(KEYINPUT55), .ZN(n1027) );
  NAND2_X1 U1043 ( .A1(n948), .A2(n1027), .ZN(n949) );
  NAND2_X1 U1044 ( .A1(n949), .A2(G29), .ZN(n1033) );
  XNOR2_X1 U1045 ( .A(G2090), .B(G35), .ZN(n954) );
  XOR2_X1 U1046 ( .A(G34), .B(KEYINPUT122), .Z(n951) );
  XNOR2_X1 U1047 ( .A(G2084), .B(KEYINPUT54), .ZN(n950) );
  XNOR2_X1 U1048 ( .A(n951), .B(n950), .ZN(n952) );
  XNOR2_X1 U1049 ( .A(n952), .B(KEYINPUT121), .ZN(n953) );
  NOR2_X1 U1050 ( .A1(n954), .A2(n953), .ZN(n969) );
  XNOR2_X1 U1051 ( .A(G2067), .B(G26), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(G33), .B(G2072), .ZN(n955) );
  NOR2_X1 U1053 ( .A1(n956), .A2(n955), .ZN(n961) );
  XNOR2_X1 U1054 ( .A(G1996), .B(G32), .ZN(n959) );
  XNOR2_X1 U1055 ( .A(G27), .B(n957), .ZN(n958) );
  NOR2_X1 U1056 ( .A1(n959), .A2(n958), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n965) );
  XNOR2_X1 U1058 ( .A(G25), .B(n962), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n963), .A2(G28), .ZN(n964) );
  NOR2_X1 U1060 ( .A1(n965), .A2(n964), .ZN(n967) );
  XOR2_X1 U1061 ( .A(KEYINPUT120), .B(KEYINPUT53), .Z(n966) );
  XNOR2_X1 U1062 ( .A(n967), .B(n966), .ZN(n968) );
  NAND2_X1 U1063 ( .A1(n969), .A2(n968), .ZN(n1026) );
  NOR2_X1 U1064 ( .A1(G29), .A2(KEYINPUT55), .ZN(n970) );
  NAND2_X1 U1065 ( .A1(n1026), .A2(n970), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(G11), .A2(n971), .ZN(n1031) );
  XNOR2_X1 U1067 ( .A(G16), .B(KEYINPUT56), .ZN(n998) );
  XNOR2_X1 U1068 ( .A(G1348), .B(n972), .ZN(n986) );
  XNOR2_X1 U1069 ( .A(n973), .B(G1956), .ZN(n979) );
  NAND2_X1 U1070 ( .A1(G1971), .A2(G303), .ZN(n974) );
  NAND2_X1 U1071 ( .A1(n975), .A2(n974), .ZN(n976) );
  NOR2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  NAND2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NOR2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  XOR2_X1 U1075 ( .A(KEYINPUT124), .B(n982), .Z(n984) );
  XNOR2_X1 U1076 ( .A(G301), .B(G1961), .ZN(n983) );
  NOR2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  NAND2_X1 U1078 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n987), .ZN(n996) );
  XNOR2_X1 U1080 ( .A(n988), .B(G1341), .ZN(n994) );
  XOR2_X1 U1081 ( .A(G1966), .B(G168), .Z(n989) );
  NOR2_X1 U1082 ( .A1(n990), .A2(n989), .ZN(n991) );
  XOR2_X1 U1083 ( .A(KEYINPUT57), .B(n991), .Z(n992) );
  XNOR2_X1 U1084 ( .A(KEYINPUT123), .B(n992), .ZN(n993) );
  NOR2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1086 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1087 ( .A1(n998), .A2(n997), .ZN(n1024) );
  XOR2_X1 U1088 ( .A(G16), .B(KEYINPUT126), .Z(n1022) );
  XOR2_X1 U1089 ( .A(G1966), .B(G21), .Z(n1009) );
  XNOR2_X1 U1090 ( .A(G20), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G19), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .Z(n1004) );
  XNOR2_X1 U1096 ( .A(G4), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1007), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1019) );
  XOR2_X1 U1100 ( .A(G1961), .B(G5), .Z(n1017) );
  XOR2_X1 U1101 ( .A(G1976), .B(G23), .Z(n1012) );
  XNOR2_X1 U1102 ( .A(n1010), .B(G22), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1014) );
  XNOR2_X1 U1104 ( .A(G24), .B(G1986), .ZN(n1013) );
  NOR2_X1 U1105 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1106 ( .A(n1015), .B(KEYINPUT58), .ZN(n1016) );
  NAND2_X1 U1107 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1108 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(n1020), .B(KEYINPUT61), .ZN(n1021) );
  NAND2_X1 U1110 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1111 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1112 ( .A(KEYINPUT127), .B(n1025), .ZN(n1029) );
  OR2_X1 U1113 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NOR2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XOR2_X1 U1117 ( .A(KEYINPUT62), .B(n1034), .Z(G311) );
  INV_X1 U1118 ( .A(G311), .ZN(G150) );
endmodule

