//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 0 0 1 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:23 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n679, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n702, new_n703, new_n704, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n911, new_n912,
    new_n913, new_n915, new_n916, new_n917, new_n918, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973;
  INV_X1    g000(.A(KEYINPUT77), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT28), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT11), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT67), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(G134), .B(G137), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT67), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n192), .B1(new_n193), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G137), .ZN(new_n197));
  AOI21_X1  g011(.A(new_n191), .B1(G134), .B2(new_n197), .ZN(new_n198));
  OAI21_X1  g012(.A(G131), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n198), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(G134), .ZN(new_n201));
  INV_X1    g015(.A(G134), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G137), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n195), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(new_n191), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT68), .B(G131), .Z(new_n206));
  NAND3_X1  g020(.A1(new_n200), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n199), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT64), .B(G146), .ZN(new_n210));
  INV_X1    g024(.A(G143), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(G146), .ZN(new_n214));
  INV_X1    g028(.A(G146), .ZN(new_n215));
  NOR2_X1   g029(.A1(new_n215), .A2(KEYINPUT64), .ZN(new_n216));
  OAI211_X1 g030(.A(KEYINPUT65), .B(G143), .C1(new_n214), .C2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n215), .A2(G143), .ZN(new_n219));
  XNOR2_X1  g033(.A(new_n219), .B(KEYINPUT66), .ZN(new_n220));
  NAND4_X1  g034(.A1(new_n218), .A2(KEYINPUT0), .A3(G128), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n215), .A2(G143), .ZN(new_n222));
  INV_X1    g036(.A(new_n210), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n223), .B2(G143), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT0), .B(G128), .Z(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n208), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT71), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT69), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n230), .B(KEYINPUT1), .C1(new_n210), .C2(new_n211), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(G143), .B1(new_n214), .B2(new_n216), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n230), .B1(new_n233), .B2(KEYINPUT1), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n224), .B1(new_n232), .B2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n218), .A2(new_n236), .A3(G128), .A4(new_n220), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n193), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(G131), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n207), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n208), .A2(new_n221), .A3(KEYINPUT71), .A4(new_n226), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n229), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G119), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G116), .ZN(new_n247));
  INV_X1    g061(.A(G116), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G119), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT2), .B(G113), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n252), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n229), .A2(new_n243), .A3(new_n254), .A4(new_n244), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n189), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n243), .A2(new_n254), .A3(new_n227), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(new_n189), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  XNOR2_X1  g073(.A(KEYINPUT72), .B(G237), .ZN(new_n260));
  INV_X1    g074(.A(G953), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n260), .A2(G210), .A3(new_n261), .ZN(new_n262));
  XNOR2_X1  g076(.A(KEYINPUT26), .B(G101), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n262), .B(new_n263), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT73), .B(KEYINPUT27), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT29), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n256), .A2(new_n259), .A3(new_n267), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n188), .B1(new_n268), .B2(KEYINPUT76), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT76), .ZN(new_n270));
  NOR4_X1   g084(.A1(new_n256), .A2(new_n270), .A3(new_n259), .A4(new_n267), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n187), .B1(new_n269), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n253), .A2(new_n255), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(KEYINPUT28), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(new_n258), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n270), .B1(new_n275), .B2(new_n267), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n268), .A2(KEYINPUT76), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n276), .A2(KEYINPUT77), .A3(new_n277), .A4(new_n188), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT30), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n241), .B1(new_n235), .B2(new_n237), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT70), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n227), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI211_X1 g096(.A(KEYINPUT70), .B(new_n241), .C1(new_n235), .C2(new_n237), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND4_X1  g098(.A1(new_n229), .A2(new_n243), .A3(KEYINPUT30), .A4(new_n244), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n284), .A2(new_n252), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n255), .ZN(new_n287));
  INV_X1    g101(.A(new_n266), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT29), .ZN(new_n290));
  NOR2_X1   g104(.A1(new_n282), .A2(new_n283), .ZN(new_n291));
  OAI21_X1  g105(.A(new_n255), .B1(new_n291), .B2(new_n254), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n292), .A2(KEYINPUT28), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n258), .ZN(new_n294));
  OAI211_X1 g108(.A(new_n289), .B(new_n290), .C1(new_n294), .C2(new_n288), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n272), .A2(new_n278), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G472), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n286), .A2(new_n255), .A3(new_n266), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT74), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n286), .A2(KEYINPUT74), .A3(new_n255), .A4(new_n266), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n300), .A2(KEYINPUT31), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n298), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n266), .B1(new_n293), .B2(new_n258), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G472), .ZN(new_n309));
  NAND4_X1  g123(.A1(new_n308), .A2(KEYINPUT32), .A3(new_n309), .A4(new_n188), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n306), .B1(new_n302), .B2(new_n304), .ZN(new_n311));
  NOR3_X1   g125(.A1(new_n311), .A2(G472), .A3(G902), .ZN(new_n312));
  XNOR2_X1  g126(.A(KEYINPUT75), .B(KEYINPUT32), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n297), .B(new_n310), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G217), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n315), .B1(G234), .B2(new_n188), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n261), .A2(G221), .A3(G234), .ZN(new_n317));
  XNOR2_X1  g131(.A(new_n317), .B(KEYINPUT79), .ZN(new_n318));
  XNOR2_X1  g132(.A(KEYINPUT22), .B(G137), .ZN(new_n319));
  XNOR2_X1  g133(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  OR2_X1    g135(.A1(KEYINPUT24), .A2(G110), .ZN(new_n322));
  INV_X1    g136(.A(G128), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G119), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n246), .A2(G128), .ZN(new_n325));
  NAND2_X1  g139(.A1(KEYINPUT24), .A2(G110), .ZN(new_n326));
  NAND4_X1  g140(.A1(new_n322), .A2(new_n324), .A3(new_n325), .A4(new_n326), .ZN(new_n327));
  OAI21_X1  g141(.A(KEYINPUT23), .B1(new_n246), .B2(G128), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT23), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(new_n323), .A3(G119), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n328), .A2(new_n330), .B1(new_n246), .B2(G128), .ZN(new_n331));
  INV_X1    g145(.A(G110), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n327), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(G140), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(G125), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(G140), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n337), .A3(KEYINPUT16), .ZN(new_n338));
  OR3_X1    g152(.A1(new_n336), .A2(KEYINPUT16), .A3(G140), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n215), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n338), .A2(new_n339), .A3(G146), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n333), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n324), .A2(new_n325), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n322), .A2(new_n326), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n331), .A2(new_n332), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AND2_X1   g160(.A1(new_n335), .A2(new_n337), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n223), .A2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(new_n342), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n346), .A2(new_n349), .ZN(new_n350));
  NOR3_X1   g164(.A1(new_n321), .A2(new_n343), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT78), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n352), .B1(new_n343), .B2(new_n350), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n341), .A2(new_n342), .ZN(new_n354));
  OR2_X1    g168(.A1(new_n331), .A2(new_n332), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n354), .A2(new_n327), .A3(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n331), .A2(new_n332), .ZN(new_n357));
  AND2_X1   g171(.A1(new_n345), .A2(new_n344), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n342), .B(new_n348), .C1(new_n357), .C2(new_n358), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n359), .A3(KEYINPUT78), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n353), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n351), .B1(new_n361), .B2(new_n321), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT25), .B1(new_n362), .B2(new_n188), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n320), .B1(new_n353), .B2(new_n360), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  NOR4_X1   g179(.A1(new_n364), .A2(new_n351), .A3(new_n365), .A4(G902), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n316), .B1(new_n363), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(KEYINPUT80), .B(new_n316), .C1(new_n363), .C2(new_n366), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n316), .A2(G902), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n362), .A2(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(G104), .ZN(new_n376));
  OAI21_X1  g190(.A(new_n375), .B1(new_n376), .B2(G107), .ZN(new_n377));
  INV_X1    g191(.A(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n378), .A2(KEYINPUT3), .A3(G104), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n380), .B1(G104), .B2(new_n378), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n381), .A2(G101), .ZN(new_n382));
  INV_X1    g196(.A(G101), .ZN(new_n383));
  OAI211_X1 g197(.A(new_n380), .B(new_n383), .C1(G104), .C2(new_n378), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n382), .A2(KEYINPUT4), .A3(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT4), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n381), .A2(new_n386), .A3(G101), .ZN(new_n387));
  NAND4_X1  g201(.A1(new_n385), .A2(new_n221), .A3(new_n226), .A4(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n238), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n378), .A2(G104), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n376), .A2(G107), .ZN(new_n391));
  OAI21_X1  g205(.A(G101), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(KEYINPUT82), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT82), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n384), .A2(new_n395), .A3(new_n392), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(KEYINPUT10), .A3(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n388), .B1(new_n389), .B2(new_n397), .ZN(new_n398));
  AND2_X1   g212(.A1(new_n218), .A2(new_n220), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n323), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n400));
  OAI21_X1  g214(.A(new_n237), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(new_n393), .ZN(new_n402));
  AOI21_X1  g216(.A(KEYINPUT10), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NOR3_X1   g217(.A1(new_n398), .A2(new_n403), .A3(new_n208), .ZN(new_n404));
  XOR2_X1   g218(.A(G110), .B(G140), .Z(new_n405));
  XNOR2_X1  g219(.A(new_n405), .B(KEYINPUT81), .ZN(new_n406));
  INV_X1    g220(.A(G227), .ZN(new_n407));
  NOR2_X1   g221(.A1(new_n407), .A2(G953), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n406), .B(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n404), .A2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(KEYINPUT85), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n208), .B1(new_n398), .B2(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT85), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n414), .B1(new_n404), .B2(new_n410), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n401), .A2(new_n402), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n394), .A2(new_n396), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n418), .A2(new_n237), .A3(new_n235), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT12), .B1(new_n208), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n420), .A2(new_n208), .A3(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n389), .A2(new_n418), .B1(new_n401), .B2(new_n402), .ZN(new_n425));
  INV_X1    g239(.A(new_n208), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n422), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n404), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g242(.A(new_n410), .B1(new_n428), .B2(KEYINPUT84), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n424), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT10), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n417), .A2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n396), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n395), .B1(new_n384), .B2(new_n392), .ZN(new_n434));
  NOR3_X1   g248(.A1(new_n433), .A2(new_n434), .A3(new_n431), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n238), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n432), .A2(new_n426), .A3(new_n388), .A4(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n430), .A2(KEYINPUT84), .A3(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  OAI211_X1 g253(.A(new_n416), .B(G469), .C1(new_n429), .C2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G469), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(new_n188), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n437), .A2(new_n413), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n410), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n423), .B1(new_n420), .B2(new_n208), .ZN(new_n445));
  AOI211_X1 g259(.A(new_n422), .B(new_n426), .C1(new_n417), .C2(new_n419), .ZN(new_n446));
  OAI211_X1 g260(.A(new_n437), .B(new_n409), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n442), .B1(new_n448), .B2(new_n441), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n440), .A2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G221), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT9), .B(G234), .Z(new_n452));
  AOI21_X1  g266(.A(new_n451), .B1(new_n452), .B2(new_n188), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n450), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n260), .A2(G214), .A3(new_n261), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n456), .A2(KEYINPUT88), .A3(new_n211), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n211), .A2(KEYINPUT88), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n260), .A2(G214), .A3(new_n261), .A4(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n457), .A2(new_n206), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT92), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n457), .A2(new_n459), .ZN(new_n462));
  INV_X1    g276(.A(new_n206), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT92), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n457), .A2(new_n465), .A3(new_n206), .A4(new_n459), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n461), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(new_n347), .B(KEYINPUT19), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(new_n223), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n467), .A2(new_n342), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(KEYINPUT18), .A2(G131), .ZN(new_n471));
  XOR2_X1   g285(.A(new_n471), .B(KEYINPUT90), .Z(new_n472));
  NAND3_X1  g286(.A1(new_n457), .A2(new_n459), .A3(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT91), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n457), .A2(KEYINPUT91), .A3(new_n459), .A4(new_n472), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT89), .ZN(new_n478));
  OR3_X1    g292(.A1(new_n347), .A2(new_n478), .A3(new_n215), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n478), .B1(new_n347), .B2(new_n215), .ZN(new_n480));
  AND2_X1   g294(.A1(new_n480), .A2(new_n348), .ZN(new_n481));
  INV_X1    g295(.A(new_n471), .ZN(new_n482));
  AOI22_X1  g296(.A1(new_n479), .A2(new_n481), .B1(new_n462), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n477), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n470), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g299(.A(G113), .B(G122), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n486), .B(new_n376), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT17), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n461), .A2(new_n464), .A3(new_n490), .A4(new_n466), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n206), .B1(new_n457), .B2(new_n459), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n354), .B1(new_n492), .B2(KEYINPUT17), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(new_n484), .A3(new_n487), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n495), .A2(KEYINPUT93), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT93), .ZN(new_n497));
  AOI22_X1  g311(.A1(new_n491), .A2(new_n493), .B1(new_n477), .B2(new_n483), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n497), .B1(new_n498), .B2(new_n487), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n489), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT20), .ZN(new_n501));
  NOR2_X1   g315(.A1(G475), .A2(G902), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n495), .A2(KEYINPUT93), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n498), .A2(new_n497), .A3(new_n487), .ZN(new_n505));
  AOI22_X1  g319(.A1(new_n504), .A2(new_n505), .B1(new_n488), .B2(new_n485), .ZN(new_n506));
  INV_X1    g320(.A(new_n502), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT20), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR2_X1   g322(.A1(new_n496), .A2(new_n499), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n498), .A2(new_n487), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n188), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI22_X1  g325(.A1(new_n503), .A2(new_n508), .B1(new_n511), .B2(G475), .ZN(new_n512));
  AOI21_X1  g326(.A(KEYINPUT13), .B1(new_n323), .B2(G143), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n513), .A2(new_n202), .ZN(new_n514));
  XNOR2_X1  g328(.A(G128), .B(G143), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  INV_X1    g330(.A(G122), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(G116), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(G116), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n378), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n519), .A2(new_n378), .A3(new_n520), .ZN(new_n522));
  INV_X1    g336(.A(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n521), .B2(new_n523), .ZN(new_n524));
  OR2_X1    g338(.A1(new_n522), .A2(KEYINPUT94), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n515), .B(new_n202), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n522), .A2(KEYINPUT94), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT14), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n520), .B1(new_n518), .B2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT95), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n530), .A2(new_n531), .B1(new_n529), .B2(new_n518), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n378), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n524), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n452), .A2(G217), .A3(new_n261), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n535), .B(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(new_n188), .ZN(new_n538));
  INV_X1    g352(.A(G478), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n539), .A2(KEYINPUT15), .ZN(new_n540));
  XOR2_X1   g354(.A(new_n538), .B(new_n540), .Z(new_n541));
  NAND2_X1  g355(.A1(new_n512), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(G234), .A2(G237), .ZN(new_n543));
  AND3_X1   g357(.A1(new_n543), .A2(G952), .A3(new_n261), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n543), .A2(G902), .A3(G953), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT96), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT21), .B(G898), .Z(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n544), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n550), .B(KEYINPUT97), .ZN(new_n551));
  INV_X1    g365(.A(new_n551), .ZN(new_n552));
  OAI21_X1  g366(.A(G214), .B1(G237), .B2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  INV_X1    g369(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT87), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n247), .A2(new_n249), .A3(KEYINPUT5), .ZN(new_n558));
  OR3_X1    g372(.A1(new_n248), .A2(KEYINPUT5), .A3(G119), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n559), .A3(G113), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT86), .ZN(new_n561));
  OR2_X1    g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n250), .A2(new_n251), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n563), .B1(new_n560), .B2(new_n561), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n394), .A2(new_n562), .A3(new_n564), .A4(new_n396), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n385), .A2(new_n252), .A3(new_n387), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n557), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  AND2_X1   g381(.A1(new_n567), .A2(KEYINPUT6), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n555), .A3(new_n566), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n569), .B1(new_n567), .B2(KEYINPUT6), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n221), .A2(new_n226), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(G125), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n235), .A2(new_n336), .A3(new_n237), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(G224), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n575), .A2(G953), .ZN(new_n576));
  NOR2_X1   g390(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(new_n576), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n578), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  OAI22_X1  g393(.A1(new_n568), .A2(new_n570), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  XOR2_X1   g394(.A(new_n555), .B(KEYINPUT8), .Z(new_n581));
  INV_X1    g395(.A(new_n563), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n394), .A2(new_n582), .A3(new_n560), .A4(new_n396), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n562), .A2(new_n564), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(new_n393), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n583), .B2(new_n585), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n565), .A2(new_n566), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n555), .B2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT7), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n574), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n579), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n572), .A2(KEYINPUT7), .A3(new_n578), .A4(new_n573), .ZN(new_n592));
  NAND4_X1  g406(.A1(new_n588), .A2(new_n590), .A3(new_n591), .A4(new_n592), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n580), .A2(new_n593), .A3(new_n188), .ZN(new_n594));
  OAI21_X1  g408(.A(G210), .B1(G237), .B2(G902), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g411(.A1(new_n580), .A2(new_n593), .A3(new_n188), .A4(new_n595), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n554), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  NOR4_X1   g414(.A1(new_n455), .A2(new_n542), .A3(new_n552), .A4(new_n600), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n314), .A2(new_n374), .A3(new_n601), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(G101), .ZN(G3));
  NAND3_X1  g417(.A1(new_n308), .A2(new_n309), .A3(new_n188), .ZN(new_n604));
  AOI211_X1 g418(.A(new_n453), .B(new_n373), .C1(new_n440), .C2(new_n449), .ZN(new_n605));
  OAI21_X1  g419(.A(G472), .B1(new_n311), .B2(G902), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(KEYINPUT98), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT98), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n604), .A2(new_n605), .A3(new_n609), .A4(new_n606), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n510), .B1(new_n504), .B2(new_n505), .ZN(new_n611));
  OAI21_X1  g425(.A(G475), .B1(new_n611), .B2(G902), .ZN(new_n612));
  NOR3_X1   g426(.A1(new_n506), .A2(KEYINPUT20), .A3(new_n507), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n501), .B1(new_n500), .B2(new_n502), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT33), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n535), .A2(new_n536), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n616), .B1(new_n617), .B2(KEYINPUT99), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n537), .B(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n539), .A2(G902), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n619), .A2(new_n620), .B1(new_n539), .B2(new_n538), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n615), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n599), .A2(new_n551), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n608), .A2(new_n610), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT100), .ZN(new_n627));
  XNOR2_X1  g441(.A(KEYINPUT34), .B(G104), .ZN(new_n628));
  XNOR2_X1  g442(.A(new_n627), .B(new_n628), .ZN(G6));
  INV_X1    g443(.A(new_n541), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n512), .A2(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n631), .A2(new_n624), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n608), .A2(new_n610), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT35), .B(G107), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  AND2_X1   g449(.A1(new_n604), .A2(new_n606), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n321), .A2(KEYINPUT36), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n361), .B(new_n637), .ZN(new_n638));
  AND3_X1   g452(.A1(new_n638), .A2(KEYINPUT101), .A3(new_n371), .ZN(new_n639));
  AOI21_X1  g453(.A(KEYINPUT101), .B1(new_n638), .B2(new_n371), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n641), .A2(new_n369), .A3(new_n370), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n601), .A2(new_n636), .A3(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  INV_X1    g459(.A(G900), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n544), .B1(new_n547), .B2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(KEYINPUT102), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n631), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n453), .B1(new_n440), .B2(new_n449), .ZN(new_n650));
  NAND3_X1  g464(.A1(new_n650), .A2(new_n599), .A3(new_n642), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n314), .A2(new_n649), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT103), .B(G128), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G30));
  NAND2_X1  g469(.A1(new_n300), .A2(new_n301), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n273), .A2(new_n288), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n657), .A2(KEYINPUT104), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n656), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(G472), .B1(new_n660), .B2(G902), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n310), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n311), .A2(G902), .ZN(new_n663));
  AOI21_X1  g477(.A(new_n313), .B1(new_n663), .B2(new_n309), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(KEYINPUT105), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n648), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n650), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT40), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n597), .A2(new_n598), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(KEYINPUT38), .ZN(new_n671));
  INV_X1    g485(.A(new_n642), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(new_n553), .A3(new_n672), .ZN(new_n673));
  NOR4_X1   g487(.A1(new_n669), .A2(new_n541), .A3(new_n512), .A4(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G143), .ZN(G45));
  NOR3_X1   g490(.A1(new_n512), .A2(new_n621), .A3(new_n648), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n297), .A2(new_n310), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n652), .B(new_n677), .C1(new_n678), .C2(new_n664), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G146), .ZN(G48));
  AOI22_X1  g494(.A1(new_n411), .A2(new_n430), .B1(new_n443), .B2(new_n410), .ZN(new_n681));
  OAI21_X1  g495(.A(G469), .B1(new_n681), .B2(G902), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n448), .A2(new_n441), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n682), .A2(new_n683), .A3(new_n454), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT106), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n682), .A2(new_n683), .A3(KEYINPUT106), .A4(new_n454), .ZN(new_n687));
  AND2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n314), .A2(new_n374), .A3(new_n625), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(KEYINPUT41), .B(G113), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  AOI22_X1  g505(.A1(new_n312), .A2(KEYINPUT32), .B1(new_n296), .B2(G472), .ZN(new_n692));
  INV_X1    g506(.A(new_n313), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n604), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n373), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n632), .A4(new_n688), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n314), .A2(new_n374), .A3(new_n632), .A4(new_n688), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n698), .A2(KEYINPUT107), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(G116), .ZN(G18));
  AND3_X1   g515(.A1(new_n686), .A2(new_n599), .A3(new_n687), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n542), .A2(new_n552), .A3(new_n672), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n314), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G119), .ZN(G21));
  NAND3_X1  g519(.A1(new_n615), .A2(new_n599), .A3(new_n630), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT109), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n615), .A2(new_n599), .A3(KEYINPUT109), .A4(new_n630), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n552), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  NAND2_X1  g524(.A1(new_n275), .A2(new_n288), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n305), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g526(.A1(G472), .A2(G902), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  XOR2_X1   g528(.A(KEYINPUT108), .B(G472), .Z(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n311), .B2(G902), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n710), .A2(new_n717), .A3(new_n374), .A4(new_n688), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G122), .ZN(G24));
  NAND4_X1  g533(.A1(new_n714), .A2(new_n716), .A3(new_n642), .A4(new_n677), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n686), .A2(new_n599), .A3(new_n687), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(new_n336), .ZN(G27));
  NOR2_X1   g537(.A1(new_n512), .A2(new_n621), .ZN(new_n724));
  INV_X1    g538(.A(new_n648), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n597), .A2(new_n553), .A3(new_n598), .ZN(new_n727));
  NOR3_X1   g541(.A1(new_n726), .A2(new_n455), .A3(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n312), .A2(KEYINPUT32), .ZN(new_n729));
  OAI211_X1 g543(.A(new_n728), .B(new_n374), .C1(new_n678), .C2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n730), .A2(KEYINPUT42), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n455), .A2(new_n727), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n726), .A2(KEYINPUT42), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n314), .A2(new_n374), .A3(new_n732), .A4(new_n733), .ZN(new_n734));
  AND2_X1   g548(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G131), .ZN(G33));
  NAND4_X1  g550(.A1(new_n314), .A2(new_n374), .A3(new_n649), .A4(new_n732), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G134), .ZN(G36));
  OAI21_X1  g552(.A(new_n416), .B1(new_n429), .B2(new_n439), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT45), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n739), .A2(new_n740), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT46), .ZN(new_n745));
  OR3_X1    g559(.A1(new_n744), .A2(new_n745), .A3(new_n442), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n745), .B1(new_n744), .B2(new_n442), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n746), .A2(new_n683), .A3(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n454), .A3(new_n667), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(KEYINPUT110), .ZN(new_n750));
  INV_X1    g564(.A(new_n727), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n512), .A2(new_n622), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n752), .A2(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n753), .A2(KEYINPUT43), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n752), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n642), .B1(new_n755), .B2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n636), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n751), .B1(new_n759), .B2(KEYINPUT44), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(KEYINPUT44), .B2(new_n759), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n750), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(G137), .ZN(G39));
  NAND2_X1  g577(.A1(new_n748), .A2(new_n454), .ZN(new_n764));
  INV_X1    g578(.A(KEYINPUT47), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NOR4_X1   g580(.A1(new_n314), .A2(new_n374), .A3(new_n726), .A4(new_n727), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G140), .ZN(G42));
  INV_X1    g583(.A(KEYINPUT113), .ZN(new_n770));
  INV_X1    g584(.A(new_n624), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n770), .B1(new_n771), .B2(new_n724), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n623), .A2(new_n624), .A3(KEYINPUT113), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n608), .A2(new_n610), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n775), .A2(new_n776), .A3(new_n602), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n633), .A2(new_n643), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n689), .A2(new_n704), .A3(new_n718), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n697), .B2(new_n699), .ZN(new_n781));
  INV_X1    g595(.A(new_n720), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n650), .A2(new_n642), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n597), .A2(new_n553), .A3(new_n598), .A4(new_n725), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n784), .B1(new_n542), .B2(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(new_n785), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT115), .A3(new_n541), .A4(new_n512), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n783), .B1(new_n786), .B2(new_n788), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n782), .A2(new_n732), .B1(new_n314), .B2(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n731), .A2(new_n790), .A3(new_n734), .A4(new_n737), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n776), .B1(new_n775), .B2(new_n602), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n779), .A2(new_n781), .A3(new_n791), .A4(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT116), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NOR3_X1   g610(.A1(new_n777), .A2(new_n792), .A3(new_n778), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n797), .A2(KEYINPUT116), .A3(new_n781), .A4(new_n791), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n796), .A2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n651), .B1(new_n692), .B2(new_n694), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n722), .B1(new_n801), .B2(new_n649), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT117), .ZN(new_n803));
  AND4_X1   g617(.A1(new_n369), .A2(new_n641), .A3(new_n370), .A4(new_n725), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n450), .A2(new_n804), .A3(new_n454), .ZN(new_n805));
  AOI21_X1  g619(.A(new_n805), .B1(new_n708), .B2(new_n709), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n806), .B1(new_n662), .B2(new_n664), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n802), .A2(new_n803), .A3(new_n679), .A4(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n717), .A2(new_n642), .A3(new_n702), .A4(new_n677), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n653), .A2(new_n679), .A3(new_n810), .A4(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT117), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(KEYINPUT52), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n815), .A2(KEYINPUT53), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n808), .A2(new_n809), .A3(new_n812), .ZN(new_n817));
  AOI21_X1  g631(.A(new_n809), .B1(new_n808), .B2(new_n812), .ZN(new_n818));
  OAI21_X1  g632(.A(KEYINPUT118), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n811), .A2(KEYINPUT117), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n811), .A2(KEYINPUT117), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT52), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT118), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n822), .A2(new_n823), .A3(new_n813), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n819), .A2(new_n796), .A3(new_n824), .A4(new_n798), .ZN(new_n825));
  AOI22_X1  g639(.A1(new_n800), .A2(new_n816), .B1(new_n825), .B2(KEYINPUT53), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n826), .A2(KEYINPUT54), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n825), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT119), .ZN(new_n830));
  INV_X1    g644(.A(new_n700), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n830), .B1(new_n831), .B2(new_n780), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n781), .A2(KEYINPUT119), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n731), .A2(KEYINPUT53), .A3(new_n734), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n790), .A2(new_n737), .ZN(new_n835));
  NOR2_X1   g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n833), .A3(new_n797), .A4(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(new_n815), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n829), .A2(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n827), .B1(KEYINPUT54), .B2(new_n840), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n544), .B1(new_n755), .B2(new_n757), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n843), .A2(new_n374), .A3(new_n717), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n682), .A2(new_n683), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(KEYINPUT112), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n846), .A2(new_n454), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n751), .B(new_n844), .C1(new_n766), .C2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n717), .A2(new_n374), .A3(new_n688), .ZN(new_n849));
  NOR4_X1   g663(.A1(new_n849), .A2(new_n842), .A3(new_n553), .A4(new_n671), .ZN(new_n850));
  INV_X1    g664(.A(new_n850), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n851), .A2(KEYINPUT50), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n851), .A2(KEYINPUT50), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n688), .A2(new_n751), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT120), .ZN(new_n855));
  AND4_X1   g669(.A1(new_n642), .A2(new_n855), .A3(new_n717), .A4(new_n843), .ZN(new_n856));
  NOR3_X1   g670(.A1(new_n852), .A2(new_n853), .A3(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(new_n666), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n858), .A2(new_n374), .A3(new_n544), .A4(new_n855), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n512), .A2(new_n621), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n848), .B(new_n857), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT51), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n861), .A2(new_n862), .ZN(new_n864));
  INV_X1    g678(.A(G952), .ZN(new_n865));
  AOI211_X1 g679(.A(new_n865), .B(G953), .C1(new_n844), .C2(new_n702), .ZN(new_n866));
  OAI21_X1  g680(.A(new_n374), .B1(new_n678), .B2(new_n729), .ZN(new_n867));
  INV_X1    g681(.A(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n855), .A2(new_n868), .A3(new_n843), .ZN(new_n869));
  INV_X1    g683(.A(new_n869), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n866), .B1(new_n870), .B2(KEYINPUT48), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n859), .A2(new_n623), .ZN(new_n872));
  AOI211_X1 g686(.A(new_n871), .B(new_n872), .C1(KEYINPUT48), .C2(new_n870), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n863), .A2(new_n864), .A3(new_n873), .ZN(new_n874));
  OAI22_X1  g688(.A1(new_n841), .A2(new_n874), .B1(G952), .B2(G953), .ZN(new_n875));
  XOR2_X1   g689(.A(new_n846), .B(KEYINPUT49), .Z(new_n876));
  INV_X1    g690(.A(new_n752), .ZN(new_n877));
  NOR4_X1   g691(.A1(new_n671), .A2(new_n373), .A3(new_n554), .A4(new_n453), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n875), .B1(new_n666), .B2(new_n879), .ZN(G75));
  AOI21_X1  g694(.A(new_n838), .B1(new_n825), .B2(new_n828), .ZN(new_n881));
  INV_X1    g695(.A(G210), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n882), .A3(new_n188), .ZN(new_n883));
  INV_X1    g697(.A(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT56), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n568), .A2(new_n570), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n886), .B(KEYINPUT121), .ZN(new_n887));
  XNOR2_X1  g701(.A(new_n887), .B(KEYINPUT55), .ZN(new_n888));
  OR2_X1    g702(.A1(new_n577), .A2(new_n579), .ZN(new_n889));
  XOR2_X1   g703(.A(new_n888), .B(new_n889), .Z(new_n890));
  INV_X1    g704(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n884), .A2(new_n885), .A3(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n883), .B2(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n865), .A2(G953), .ZN(new_n894));
  XOR2_X1   g708(.A(new_n894), .B(KEYINPUT122), .Z(new_n895));
  NAND3_X1  g709(.A1(new_n892), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT123), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n892), .A2(new_n893), .A3(KEYINPUT123), .A4(new_n895), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(G51));
  INV_X1    g714(.A(new_n895), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n881), .A2(new_n188), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n902), .A2(new_n744), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT124), .Z(new_n904));
  XNOR2_X1  g718(.A(new_n840), .B(KEYINPUT54), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n442), .B(KEYINPUT57), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n681), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n901), .B1(new_n904), .B2(new_n909), .ZN(G54));
  AND3_X1   g724(.A1(new_n902), .A2(KEYINPUT58), .A3(G475), .ZN(new_n911));
  OR2_X1    g725(.A1(new_n911), .A2(new_n506), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n506), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n901), .B1(new_n912), .B2(new_n913), .ZN(G60));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT59), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n905), .A2(new_n619), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n619), .B1(new_n841), .B2(new_n916), .ZN(new_n918));
  NOR3_X1   g732(.A1(new_n917), .A2(new_n901), .A3(new_n918), .ZN(G63));
  NAND2_X1  g733(.A1(G217), .A2(G902), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n920), .B(KEYINPUT60), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n840), .A2(new_n638), .A3(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(new_n362), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n881), .B2(new_n921), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n895), .A3(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(KEYINPUT126), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT125), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT61), .B1(new_n923), .B2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT126), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n923), .A2(new_n925), .A3(new_n930), .A4(new_n895), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n929), .B1(new_n927), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n932), .A2(new_n933), .ZN(G66));
  NAND2_X1  g748(.A1(new_n797), .A2(new_n781), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n261), .ZN(new_n936));
  OAI21_X1  g750(.A(G953), .B1(new_n549), .B2(new_n575), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g752(.A(new_n887), .B1(G898), .B2(new_n261), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(G69));
  AND2_X1   g754(.A1(new_n762), .A2(new_n768), .ZN(new_n941));
  AND2_X1   g755(.A1(new_n802), .A2(new_n679), .ZN(new_n942));
  INV_X1    g756(.A(new_n737), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n708), .A2(new_n709), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n868), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n943), .B1(new_n750), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n941), .A2(new_n735), .A3(new_n942), .A4(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n284), .A2(new_n285), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(new_n468), .Z(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g766(.A(G953), .B1(new_n949), .B2(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n942), .A2(new_n675), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT62), .Z(new_n955));
  NAND2_X1  g769(.A1(new_n631), .A2(new_n623), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n668), .A2(new_n727), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n695), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n941), .A2(new_n955), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n951), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n952), .A2(G227), .ZN(new_n961));
  AOI211_X1 g775(.A(new_n646), .B(new_n261), .C1(new_n951), .C2(new_n407), .ZN(new_n962));
  AOI22_X1  g776(.A1(new_n953), .A2(new_n960), .B1(new_n961), .B2(new_n962), .ZN(G72));
  NAND2_X1  g777(.A1(G472), .A2(G902), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT63), .Z(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n948), .B2(new_n935), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n966), .A2(new_n255), .A3(new_n288), .A4(new_n286), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n965), .B1(new_n959), .B2(new_n935), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n968), .A2(new_n266), .A3(new_n287), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n967), .A2(new_n895), .A3(new_n969), .ZN(new_n970));
  INV_X1    g784(.A(new_n965), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n971), .B1(new_n656), .B2(new_n289), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT127), .Z(new_n973));
  AOI21_X1  g787(.A(new_n970), .B1(new_n826), .B2(new_n973), .ZN(G57));
endmodule


