

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n464, n465, n466, n467, n468, n469, n470, n471,
         n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
         n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493,
         n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504,
         n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515,
         n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772;

  XNOR2_X1 U371 ( .A(n436), .B(n362), .ZN(n556) );
  XNOR2_X1 U372 ( .A(n461), .B(n460), .ZN(n506) );
  XNOR2_X1 U373 ( .A(n468), .B(n522), .ZN(n748) );
  XNOR2_X1 U374 ( .A(n483), .B(n482), .ZN(n371) );
  INV_X4 U375 ( .A(G953), .ZN(n743) );
  XNOR2_X1 U376 ( .A(n481), .B(n480), .ZN(n483) );
  NAND2_X1 U377 ( .A1(n648), .A2(n365), .ZN(n650) );
  XNOR2_X2 U378 ( .A(n585), .B(KEYINPUT45), .ZN(n365) );
  XNOR2_X2 U379 ( .A(n350), .B(KEYINPUT85), .ZN(n458) );
  NAND2_X2 U380 ( .A1(n572), .A2(n571), .ZN(n350) );
  AND2_X2 U381 ( .A1(n451), .A2(G469), .ZN(n360) );
  INV_X1 U382 ( .A(n556), .ZN(n563) );
  INV_X1 U383 ( .A(n573), .ZN(n701) );
  XNOR2_X1 U384 ( .A(n575), .B(KEYINPUT106), .ZN(n770) );
  XOR2_X1 U385 ( .A(n471), .B(n470), .Z(n351) );
  XOR2_X1 U386 ( .A(n600), .B(KEYINPUT30), .Z(n352) );
  NAND2_X1 U387 ( .A1(n453), .A2(KEYINPUT84), .ZN(n452) );
  NOR2_X1 U388 ( .A1(n411), .A2(n618), .ZN(n620) );
  NAND2_X1 U389 ( .A1(n770), .A2(n768), .ZN(n581) );
  XNOR2_X1 U390 ( .A(n542), .B(KEYINPUT22), .ZN(n409) );
  XOR2_X1 U391 ( .A(n701), .B(KEYINPUT105), .Z(n606) );
  XNOR2_X1 U392 ( .A(n501), .B(n500), .ZN(n565) );
  XNOR2_X1 U393 ( .A(n528), .B(n429), .ZN(n505) );
  XOR2_X1 U394 ( .A(n353), .B(KEYINPUT95), .Z(n706) );
  NAND2_X1 U395 ( .A1(n697), .A2(n449), .ZN(n353) );
  BUF_X1 U396 ( .A(n400), .Z(n354) );
  BUF_X1 U397 ( .A(n768), .Z(n355) );
  XNOR2_X1 U398 ( .A(n578), .B(KEYINPUT32), .ZN(n768) );
  NAND2_X1 U399 ( .A1(n553), .A2(n555), .ZN(n356) );
  NAND2_X1 U400 ( .A1(n553), .A2(n555), .ZN(n656) );
  XNOR2_X2 U401 ( .A(n633), .B(n428), .ZN(n427) );
  AND2_X1 U402 ( .A1(n446), .A2(n357), .ZN(n445) );
  AND2_X2 U403 ( .A1(n455), .A2(n584), .ZN(n359) );
  AND2_X2 U404 ( .A1(n451), .A2(n730), .ZN(n738) );
  XOR2_X1 U405 ( .A(KEYINPUT67), .B(G131), .Z(n496) );
  XNOR2_X1 U406 ( .A(n469), .B(G140), .ZN(n754) );
  XNOR2_X1 U407 ( .A(n529), .B(KEYINPUT10), .ZN(n469) );
  INV_X1 U408 ( .A(KEYINPUT48), .ZN(n428) );
  INV_X1 U409 ( .A(KEYINPUT8), .ZN(n460) );
  NAND2_X1 U410 ( .A1(n743), .A2(G234), .ZN(n461) );
  XOR2_X1 U411 ( .A(G137), .B(KEYINPUT68), .Z(n547) );
  XNOR2_X1 U412 ( .A(n488), .B(G472), .ZN(n573) );
  XNOR2_X1 U413 ( .A(n476), .B(KEYINPUT25), .ZN(n477) );
  XNOR2_X1 U414 ( .A(n505), .B(n479), .ZN(n549) );
  NOR2_X1 U415 ( .A1(n676), .A2(n605), .ZN(n613) );
  XNOR2_X1 U416 ( .A(G104), .B(G122), .ZN(n492) );
  XNOR2_X1 U417 ( .A(G113), .B(G143), .ZN(n497) );
  NAND2_X1 U418 ( .A1(n607), .A2(n606), .ZN(n383) );
  INV_X1 U419 ( .A(KEYINPUT28), .ZN(n382) );
  NAND2_X1 U420 ( .A1(n537), .A2(G214), .ZN(n684) );
  XOR2_X1 U421 ( .A(KEYINPUT90), .B(n534), .Z(n535) );
  NOR2_X1 U422 ( .A1(n680), .A2(n385), .ZN(n384) );
  INV_X1 U423 ( .A(n679), .ZN(n385) );
  XOR2_X1 U424 ( .A(KEYINPUT74), .B(KEYINPUT16), .Z(n523) );
  XNOR2_X1 U425 ( .A(n464), .B(n754), .ZN(n651) );
  XNOR2_X1 U426 ( .A(n465), .B(n472), .ZN(n464) );
  XNOR2_X1 U427 ( .A(n351), .B(n466), .ZN(n465) );
  INV_X1 U428 ( .A(G134), .ZN(n429) );
  XNOR2_X1 U429 ( .A(G107), .B(G116), .ZN(n502) );
  XOR2_X1 U430 ( .A(KEYINPUT9), .B(G122), .Z(n503) );
  XNOR2_X1 U431 ( .A(n628), .B(n430), .ZN(n638) );
  INV_X1 U432 ( .A(KEYINPUT39), .ZN(n430) );
  NOR2_X1 U433 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U434 ( .A(G478), .B(n512), .Z(n566) );
  INV_X1 U435 ( .A(KEYINPUT99), .ZN(n395) );
  INV_X1 U436 ( .A(KEYINPUT22), .ZN(n402) );
  NAND2_X1 U437 ( .A1(n407), .A2(G472), .ZN(n424) );
  NAND2_X1 U438 ( .A1(n738), .A2(G217), .ZN(n393) );
  INV_X1 U439 ( .A(n651), .ZN(n392) );
  INV_X1 U440 ( .A(n671), .ZN(n668) );
  AND2_X1 U441 ( .A1(n698), .A2(n701), .ZN(n449) );
  XNOR2_X1 U442 ( .A(n547), .B(n473), .ZN(n466) );
  INV_X1 U443 ( .A(KEYINPUT73), .ZN(n397) );
  XNOR2_X1 U444 ( .A(G902), .B(KEYINPUT15), .ZN(n645) );
  XOR2_X1 U445 ( .A(G125), .B(G146), .Z(n529) );
  XOR2_X1 U446 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n526) );
  NAND2_X1 U447 ( .A1(G237), .A2(G234), .ZN(n516) );
  INV_X1 U448 ( .A(KEYINPUT31), .ZN(n439) );
  XNOR2_X1 U449 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n538) );
  XNOR2_X1 U450 ( .A(n377), .B(n376), .ZN(n375) );
  XNOR2_X1 U451 ( .A(KEYINPUT5), .B(KEYINPUT94), .ZN(n377) );
  XNOR2_X1 U452 ( .A(G146), .B(G137), .ZN(n376) );
  XNOR2_X1 U453 ( .A(n414), .B(n499), .ZN(n654) );
  XNOR2_X1 U454 ( .A(n754), .B(n498), .ZN(n414) );
  XOR2_X1 U455 ( .A(G146), .B(G140), .Z(n544) );
  XNOR2_X1 U456 ( .A(n549), .B(n548), .ZN(n755) );
  INV_X1 U457 ( .A(KEYINPUT33), .ZN(n404) );
  NOR2_X1 U458 ( .A1(n757), .A2(n647), .ZN(n648) );
  XNOR2_X1 U459 ( .A(n380), .B(n379), .ZN(n624) );
  INV_X1 U460 ( .A(KEYINPUT109), .ZN(n379) );
  XNOR2_X1 U461 ( .A(n383), .B(n382), .ZN(n381) );
  NAND2_X1 U462 ( .A1(n369), .A2(n425), .ZN(n437) );
  NOR2_X1 U463 ( .A1(n563), .A2(n439), .ZN(n369) );
  NAND2_X1 U464 ( .A1(n352), .A2(n431), .ZN(n627) );
  NOR2_X1 U465 ( .A1(n601), .A2(n432), .ZN(n431) );
  INV_X1 U466 ( .A(n602), .ZN(n432) );
  NAND2_X1 U467 ( .A1(n372), .A2(n373), .ZN(n400) );
  NAND2_X1 U468 ( .A1(n374), .A2(n403), .ZN(n373) );
  XOR2_X1 U469 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n508) );
  NAND2_X1 U470 ( .A1(n407), .A2(G475), .ZN(n388) );
  XNOR2_X1 U471 ( .A(n629), .B(KEYINPUT40), .ZN(n771) );
  AND2_X1 U472 ( .A1(n638), .A2(n668), .ZN(n629) );
  NOR2_X1 U473 ( .A1(n622), .A2(n634), .ZN(n597) );
  AND2_X1 U474 ( .A1(n574), .A2(n417), .ZN(n416) );
  NAND2_X1 U475 ( .A1(n415), .A2(n565), .ZN(n671) );
  NAND2_X1 U476 ( .A1(n367), .A2(n366), .ZN(n658) );
  NOR2_X1 U477 ( .A1(n601), .A2(n701), .ZN(n366) );
  AND2_X1 U478 ( .A1(n443), .A2(n358), .ZN(n419) );
  XNOR2_X1 U479 ( .A(n424), .B(n363), .ZN(n420) );
  INV_X1 U480 ( .A(KEYINPUT124), .ZN(n389) );
  INV_X1 U481 ( .A(KEYINPUT56), .ZN(n421) );
  OR2_X1 U482 ( .A1(n448), .A2(KEYINPUT83), .ZN(n357) );
  XNOR2_X1 U483 ( .A(KEYINPUT102), .B(n594), .ZN(n358) );
  INV_X1 U484 ( .A(n680), .ZN(n426) );
  INV_X1 U485 ( .A(n706), .ZN(n425) );
  XOR2_X1 U486 ( .A(KEYINPUT65), .B(KEYINPUT1), .Z(n361) );
  INV_X1 U487 ( .A(n467), .ZN(n448) );
  INV_X1 U488 ( .A(KEYINPUT83), .ZN(n447) );
  XNOR2_X1 U489 ( .A(KEYINPUT0), .B(KEYINPUT86), .ZN(n362) );
  XOR2_X1 U490 ( .A(n652), .B(KEYINPUT62), .Z(n363) );
  XOR2_X1 U491 ( .A(n654), .B(n653), .Z(n364) );
  INV_X1 U492 ( .A(KEYINPUT84), .ZN(n462) );
  NOR2_X1 U493 ( .A1(G952), .A2(n743), .ZN(n742) );
  NAND2_X1 U494 ( .A1(n644), .A2(n365), .ZN(n681) );
  NAND2_X1 U495 ( .A1(n365), .A2(n743), .ZN(n747) );
  NAND2_X1 U496 ( .A1(n368), .A2(n658), .ZN(n440) );
  INV_X1 U497 ( .A(n563), .ZN(n367) );
  NAND2_X1 U498 ( .A1(n438), .A2(n437), .ZN(n368) );
  NAND2_X1 U499 ( .A1(n370), .A2(n439), .ZN(n438) );
  NAND2_X1 U500 ( .A1(n367), .A2(n425), .ZN(n370) );
  INV_X1 U501 ( .A(n371), .ZN(n374) );
  NAND2_X1 U502 ( .A1(n371), .A2(n524), .ZN(n372) );
  XNOR2_X1 U503 ( .A(n371), .B(n549), .ZN(n487) );
  XNOR2_X1 U504 ( .A(n521), .B(n375), .ZN(n485) );
  XNOR2_X2 U505 ( .A(n378), .B(KEYINPUT4), .ZN(n521) );
  XNOR2_X2 U506 ( .A(G101), .B(KEYINPUT66), .ZN(n378) );
  NAND2_X1 U507 ( .A1(n381), .A2(n608), .ZN(n380) );
  NAND2_X1 U508 ( .A1(n427), .A2(n426), .ZN(n643) );
  NAND2_X1 U509 ( .A1(n427), .A2(n384), .ZN(n757) );
  XNOR2_X1 U510 ( .A(n400), .B(n546), .ZN(n441) );
  XNOR2_X1 U511 ( .A(n386), .B(n655), .ZN(G60) );
  NAND2_X1 U512 ( .A1(n387), .A2(n729), .ZN(n386) );
  XNOR2_X1 U513 ( .A(n388), .B(n364), .ZN(n387) );
  XNOR2_X1 U514 ( .A(n390), .B(n389), .ZN(G66) );
  NAND2_X1 U515 ( .A1(n391), .A2(n729), .ZN(n390) );
  XNOR2_X1 U516 ( .A(n393), .B(n392), .ZN(n391) );
  BUF_X1 U517 ( .A(n718), .Z(n394) );
  XNOR2_X1 U518 ( .A(n405), .B(n404), .ZN(n718) );
  XNOR2_X1 U519 ( .A(n511), .B(n395), .ZN(n512) );
  NAND2_X1 U520 ( .A1(n521), .A2(KEYINPUT73), .ZN(n398) );
  NAND2_X1 U521 ( .A1(n396), .A2(n397), .ZN(n399) );
  NAND2_X1 U522 ( .A1(n398), .A2(n399), .ZN(n442) );
  INV_X1 U523 ( .A(n521), .ZN(n396) );
  XNOR2_X1 U524 ( .A(n542), .B(n402), .ZN(n401) );
  INV_X1 U525 ( .A(n524), .ZN(n403) );
  XNOR2_X1 U526 ( .A(n523), .B(G122), .ZN(n524) );
  NAND2_X1 U527 ( .A1(n562), .A2(n467), .ZN(n405) );
  BUF_X1 U528 ( .A(n438), .Z(n406) );
  AND2_X2 U529 ( .A1(n730), .A2(n451), .ZN(n407) );
  INV_X1 U530 ( .A(n606), .ZN(n417) );
  BUF_X1 U531 ( .A(n586), .Z(n637) );
  XNOR2_X1 U532 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U533 ( .A(n550), .B(n755), .ZN(n734) );
  XNOR2_X1 U534 ( .A(n546), .B(n545), .ZN(n550) );
  BUF_X1 U535 ( .A(n697), .Z(n435) );
  BUF_X1 U536 ( .A(n724), .Z(n408) );
  XNOR2_X1 U537 ( .A(n441), .B(n532), .ZN(n724) );
  NAND2_X1 U538 ( .A1(n406), .A2(n437), .ZN(n410) );
  NAND2_X1 U539 ( .A1(n617), .A2(n616), .ZN(n411) );
  XNOR2_X1 U540 ( .A(n354), .B(n749), .ZN(n750) );
  XNOR2_X2 U541 ( .A(n442), .B(n748), .ZN(n546) );
  XNOR2_X1 U542 ( .A(n412), .B(KEYINPUT122), .ZN(G54) );
  NOR2_X2 U543 ( .A1(n737), .A2(n742), .ZN(n412) );
  NAND2_X1 U544 ( .A1(n582), .A2(KEYINPUT44), .ZN(n571) );
  XNOR2_X2 U545 ( .A(n570), .B(KEYINPUT35), .ZN(n582) );
  INV_X1 U546 ( .A(n435), .ZN(n555) );
  NAND2_X1 U547 ( .A1(n697), .A2(n698), .ZN(n450) );
  XNOR2_X2 U548 ( .A(n557), .B(n361), .ZN(n697) );
  XNOR2_X1 U549 ( .A(n413), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U550 ( .A1(n420), .A2(n729), .ZN(n413) );
  NAND2_X1 U551 ( .A1(n569), .A2(n568), .ZN(n570) );
  XNOR2_X1 U552 ( .A(n539), .B(n538), .ZN(n609) );
  INV_X1 U553 ( .A(n566), .ZN(n415) );
  NAND2_X1 U554 ( .A1(n581), .A2(KEYINPUT44), .ZN(n579) );
  NAND2_X1 U555 ( .A1(n418), .A2(n416), .ZN(n575) );
  INV_X1 U556 ( .A(n409), .ZN(n418) );
  NOR2_X1 U557 ( .A1(n467), .A2(n447), .ZN(n444) );
  NOR2_X2 U558 ( .A1(n609), .A2(n540), .ZN(n436) );
  AND2_X2 U559 ( .A1(n445), .A2(n419), .ZN(n553) );
  NAND2_X1 U560 ( .A1(n556), .A2(n541), .ZN(n542) );
  XNOR2_X1 U561 ( .A(n422), .B(n421), .ZN(G51) );
  NAND2_X1 U562 ( .A1(n434), .A2(n729), .ZN(n422) );
  NOR2_X2 U563 ( .A1(G902), .A2(n734), .ZN(n552) );
  NAND2_X1 U564 ( .A1(n423), .A2(n656), .ZN(n561) );
  XNOR2_X1 U565 ( .A(n459), .B(KEYINPUT100), .ZN(n423) );
  XNOR2_X2 U566 ( .A(G128), .B(G143), .ZN(n528) );
  NAND2_X1 U567 ( .A1(n418), .A2(n433), .ZN(n578) );
  AND2_X1 U568 ( .A1(n577), .A2(n448), .ZN(n433) );
  XNOR2_X1 U569 ( .A(n727), .B(n728), .ZN(n434) );
  OR2_X2 U570 ( .A1(n580), .A2(n462), .ZN(n455) );
  XNOR2_X1 U571 ( .A(n579), .B(KEYINPUT64), .ZN(n580) );
  NAND2_X1 U572 ( .A1(n440), .A2(n560), .ZN(n459) );
  NAND2_X1 U573 ( .A1(n401), .A2(n444), .ZN(n443) );
  NAND2_X1 U574 ( .A1(n409), .A2(n447), .ZN(n446) );
  XNOR2_X1 U575 ( .A(n450), .B(KEYINPUT107), .ZN(n562) );
  XNOR2_X1 U576 ( .A(n487), .B(n486), .ZN(n652) );
  AND2_X2 U577 ( .A1(n681), .A2(n646), .ZN(n730) );
  NAND2_X2 U578 ( .A1(n650), .A2(n649), .ZN(n451) );
  NAND2_X1 U579 ( .A1(n682), .A2(n451), .ZN(n717) );
  NAND2_X2 U580 ( .A1(n454), .A2(n452), .ZN(n585) );
  INV_X1 U581 ( .A(n458), .ZN(n453) );
  AND2_X2 U582 ( .A1(n456), .A2(n359), .ZN(n454) );
  NAND2_X1 U583 ( .A1(n458), .A2(n457), .ZN(n456) );
  AND2_X1 U584 ( .A1(n580), .A2(n462), .ZN(n457) );
  XNOR2_X1 U585 ( .A(n736), .B(n735), .ZN(n737) );
  XNOR2_X2 U586 ( .A(G119), .B(G116), .ZN(n481) );
  AND2_X2 U587 ( .A1(n594), .A2(n554), .ZN(n698) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n573), .ZN(n467) );
  XOR2_X1 U589 ( .A(G104), .B(G107), .Z(n468) );
  INV_X1 U590 ( .A(KEYINPUT69), .ZN(n619) );
  XNOR2_X1 U591 ( .A(n630), .B(KEYINPUT46), .ZN(n631) );
  INV_X1 U592 ( .A(n496), .ZN(n479) );
  XNOR2_X1 U593 ( .A(n529), .B(n528), .ZN(n530) );
  INV_X1 U594 ( .A(n547), .ZN(n548) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(n532) );
  INV_X1 U596 ( .A(G469), .ZN(n551) );
  OR2_X1 U597 ( .A1(n624), .A2(n609), .ZN(n614) );
  NAND2_X1 U598 ( .A1(G221), .A2(n506), .ZN(n472) );
  XOR2_X1 U599 ( .A(G128), .B(G119), .Z(n471) );
  XNOR2_X1 U600 ( .A(KEYINPUT82), .B(G110), .ZN(n470) );
  XNOR2_X1 U601 ( .A(KEYINPUT23), .B(KEYINPUT24), .ZN(n473) );
  NOR2_X1 U602 ( .A1(G902), .A2(n651), .ZN(n478) );
  NAND2_X1 U603 ( .A1(n645), .A2(G234), .ZN(n475) );
  XNOR2_X1 U604 ( .A(KEYINPUT92), .B(KEYINPUT20), .ZN(n474) );
  XNOR2_X1 U605 ( .A(n475), .B(n474), .ZN(n513) );
  NAND2_X1 U606 ( .A1(G217), .A2(n513), .ZN(n476) );
  XNOR2_X2 U607 ( .A(n478), .B(n477), .ZN(n594) );
  INV_X1 U608 ( .A(KEYINPUT3), .ZN(n480) );
  XOR2_X1 U609 ( .A(KEYINPUT72), .B(G113), .Z(n482) );
  NOR2_X1 U610 ( .A1(G953), .A2(G237), .ZN(n489) );
  NAND2_X1 U611 ( .A1(n489), .A2(G210), .ZN(n484) );
  XNOR2_X1 U612 ( .A(n485), .B(n484), .ZN(n486) );
  NOR2_X1 U613 ( .A1(n652), .A2(G902), .ZN(n488) );
  XNOR2_X1 U614 ( .A(KEYINPUT13), .B(G475), .ZN(n501) );
  XOR2_X1 U615 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n491) );
  NAND2_X1 U616 ( .A1(n489), .A2(G214), .ZN(n490) );
  XNOR2_X1 U617 ( .A(n491), .B(n490), .ZN(n495) );
  XOR2_X1 U618 ( .A(KEYINPUT96), .B(KEYINPUT11), .Z(n493) );
  XNOR2_X1 U619 ( .A(n493), .B(n492), .ZN(n494) );
  XOR2_X1 U620 ( .A(n495), .B(n494), .Z(n499) );
  XNOR2_X1 U621 ( .A(n497), .B(n496), .ZN(n498) );
  NOR2_X1 U622 ( .A1(G902), .A2(n654), .ZN(n500) );
  XNOR2_X1 U623 ( .A(n503), .B(n502), .ZN(n504) );
  XOR2_X1 U624 ( .A(n505), .B(n504), .Z(n510) );
  NAND2_X1 U625 ( .A1(G217), .A2(n506), .ZN(n507) );
  XNOR2_X1 U626 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U627 ( .A(n510), .B(n509), .ZN(n740) );
  NOR2_X1 U628 ( .A1(G902), .A2(n740), .ZN(n511) );
  NOR2_X1 U629 ( .A1(n565), .A2(n566), .ZN(n621) );
  NAND2_X1 U630 ( .A1(n513), .A2(G221), .ZN(n514) );
  XOR2_X1 U631 ( .A(KEYINPUT21), .B(n514), .Z(n695) );
  XOR2_X1 U632 ( .A(KEYINPUT93), .B(n695), .Z(n554) );
  NAND2_X1 U633 ( .A1(n621), .A2(n554), .ZN(n515) );
  XNOR2_X1 U634 ( .A(KEYINPUT101), .B(n515), .ZN(n541) );
  XNOR2_X1 U635 ( .A(n516), .B(KEYINPUT14), .ZN(n518) );
  NAND2_X1 U636 ( .A1(n518), .A2(G952), .ZN(n517) );
  XNOR2_X1 U637 ( .A(n517), .B(KEYINPUT91), .ZN(n714) );
  NAND2_X1 U638 ( .A1(n714), .A2(n743), .ZN(n591) );
  NAND2_X1 U639 ( .A1(G902), .A2(n518), .ZN(n588) );
  INV_X1 U640 ( .A(n588), .ZN(n519) );
  NOR2_X1 U641 ( .A1(G898), .A2(n743), .ZN(n751) );
  NAND2_X1 U642 ( .A1(n519), .A2(n751), .ZN(n520) );
  AND2_X1 U643 ( .A1(n591), .A2(n520), .ZN(n540) );
  XNOR2_X1 U644 ( .A(G110), .B(KEYINPUT88), .ZN(n522) );
  NAND2_X1 U645 ( .A1(G224), .A2(n743), .ZN(n525) );
  XNOR2_X1 U646 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U647 ( .A(n527), .B(KEYINPUT89), .Z(n531) );
  NAND2_X1 U648 ( .A1(n724), .A2(n645), .ZN(n536) );
  NOR2_X1 U649 ( .A1(G902), .A2(G237), .ZN(n533) );
  XOR2_X1 U650 ( .A(KEYINPUT76), .B(n533), .Z(n537) );
  NAND2_X1 U651 ( .A1(n537), .A2(G210), .ZN(n534) );
  XNOR2_X2 U652 ( .A(n536), .B(n535), .ZN(n586) );
  NAND2_X1 U653 ( .A1(n586), .A2(n684), .ZN(n539) );
  NAND2_X1 U654 ( .A1(G227), .A2(n743), .ZN(n543) );
  XNOR2_X1 U655 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X2 U656 ( .A(n552), .B(n551), .ZN(n557) );
  INV_X1 U657 ( .A(n557), .ZN(n558) );
  INV_X1 U658 ( .A(n558), .ZN(n608) );
  NAND2_X1 U659 ( .A1(n608), .A2(n698), .ZN(n601) );
  INV_X1 U660 ( .A(n565), .ZN(n559) );
  NAND2_X1 U661 ( .A1(n559), .A2(n566), .ZN(n673) );
  INV_X1 U662 ( .A(n673), .ZN(n664) );
  NOR2_X1 U663 ( .A1(n668), .A2(n664), .ZN(n688) );
  INV_X1 U664 ( .A(n688), .ZN(n560) );
  XNOR2_X1 U665 ( .A(n561), .B(KEYINPUT103), .ZN(n572) );
  NOR2_X1 U666 ( .A1(n563), .A2(n718), .ZN(n564) );
  XNOR2_X1 U667 ( .A(n564), .B(KEYINPUT34), .ZN(n569) );
  NAND2_X1 U668 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U669 ( .A(n567), .B(KEYINPUT108), .ZN(n603) );
  INV_X1 U670 ( .A(n603), .ZN(n568) );
  NOR2_X1 U671 ( .A1(n435), .A2(n594), .ZN(n574) );
  XNOR2_X1 U672 ( .A(KEYINPUT87), .B(n697), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n599), .A2(n358), .ZN(n576) );
  XNOR2_X1 U674 ( .A(KEYINPUT104), .B(n576), .ZN(n577) );
  NOR2_X1 U675 ( .A1(n581), .A2(KEYINPUT44), .ZN(n583) );
  INV_X1 U676 ( .A(n582), .ZN(n767) );
  NAND2_X1 U677 ( .A1(n583), .A2(n767), .ZN(n584) );
  INV_X1 U678 ( .A(n637), .ZN(n622) );
  NAND2_X1 U679 ( .A1(n467), .A2(n684), .ZN(n587) );
  NOR2_X1 U680 ( .A1(n671), .A2(n587), .ZN(n596) );
  NOR2_X1 U681 ( .A1(G900), .A2(n588), .ZN(n589) );
  NAND2_X1 U682 ( .A1(G953), .A2(n589), .ZN(n590) );
  NAND2_X1 U683 ( .A1(n591), .A2(n590), .ZN(n602) );
  NAND2_X1 U684 ( .A1(n695), .A2(n602), .ZN(n592) );
  XOR2_X1 U685 ( .A(KEYINPUT71), .B(n592), .Z(n593) );
  NOR2_X1 U686 ( .A1(n594), .A2(n593), .ZN(n595) );
  XNOR2_X1 U687 ( .A(KEYINPUT70), .B(n595), .ZN(n607) );
  NAND2_X1 U688 ( .A1(n596), .A2(n607), .ZN(n634) );
  XOR2_X1 U689 ( .A(KEYINPUT36), .B(n597), .Z(n598) );
  NOR2_X1 U690 ( .A1(n599), .A2(n598), .ZN(n676) );
  NAND2_X1 U691 ( .A1(n606), .A2(n684), .ZN(n600) );
  NOR2_X1 U692 ( .A1(n603), .A2(n627), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n604), .A2(n637), .ZN(n667) );
  XNOR2_X1 U694 ( .A(KEYINPUT81), .B(n667), .ZN(n605) );
  INV_X1 U695 ( .A(n614), .ZN(n669) );
  NOR2_X1 U696 ( .A1(KEYINPUT47), .A2(n688), .ZN(n610) );
  XOR2_X1 U697 ( .A(KEYINPUT75), .B(n610), .Z(n611) );
  NAND2_X1 U698 ( .A1(n669), .A2(n611), .ZN(n612) );
  NAND2_X1 U699 ( .A1(n613), .A2(n612), .ZN(n618) );
  NAND2_X1 U700 ( .A1(n614), .A2(KEYINPUT47), .ZN(n615) );
  XNOR2_X1 U701 ( .A(n615), .B(KEYINPUT80), .ZN(n617) );
  NAND2_X1 U702 ( .A1(n688), .A2(KEYINPUT47), .ZN(n616) );
  XNOR2_X1 U703 ( .A(n620), .B(n619), .ZN(n632) );
  INV_X1 U704 ( .A(n621), .ZN(n686) );
  XOR2_X1 U705 ( .A(n622), .B(KEYINPUT38), .Z(n626) );
  INV_X1 U706 ( .A(n626), .ZN(n683) );
  NAND2_X1 U707 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U708 ( .A1(n686), .A2(n689), .ZN(n623) );
  XNOR2_X1 U709 ( .A(n623), .B(KEYINPUT41), .ZN(n719) );
  NOR2_X1 U710 ( .A1(n719), .A2(n624), .ZN(n625) );
  XNOR2_X1 U711 ( .A(n625), .B(KEYINPUT42), .ZN(n772) );
  NOR2_X1 U712 ( .A1(n772), .A2(n771), .ZN(n630) );
  NAND2_X1 U713 ( .A1(n632), .A2(n631), .ZN(n633) );
  NOR2_X1 U714 ( .A1(n435), .A2(n634), .ZN(n635) );
  XNOR2_X1 U715 ( .A(n635), .B(KEYINPUT43), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n680) );
  INV_X1 U717 ( .A(KEYINPUT78), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n638), .A2(n664), .ZN(n679) );
  NAND2_X1 U719 ( .A1(n647), .A2(n679), .ZN(n641) );
  NAND2_X1 U720 ( .A1(n679), .A2(KEYINPUT2), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n639), .A2(KEYINPUT78), .ZN(n640) );
  NAND2_X1 U722 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U723 ( .A1(n643), .A2(n642), .ZN(n644) );
  INV_X1 U724 ( .A(n645), .ZN(n646) );
  INV_X1 U725 ( .A(KEYINPUT2), .ZN(n649) );
  INV_X1 U726 ( .A(KEYINPUT60), .ZN(n655) );
  XNOR2_X1 U727 ( .A(KEYINPUT59), .B(KEYINPUT123), .ZN(n653) );
  INV_X1 U728 ( .A(n742), .ZN(n729) );
  XNOR2_X1 U729 ( .A(n356), .B(G101), .ZN(G3) );
  NOR2_X1 U730 ( .A1(n671), .A2(n658), .ZN(n657) );
  XOR2_X1 U731 ( .A(G104), .B(n657), .Z(G6) );
  NOR2_X1 U732 ( .A1(n673), .A2(n658), .ZN(n663) );
  XOR2_X1 U733 ( .A(KEYINPUT110), .B(KEYINPUT111), .Z(n660) );
  XNOR2_X1 U734 ( .A(G107), .B(KEYINPUT26), .ZN(n659) );
  XNOR2_X1 U735 ( .A(n660), .B(n659), .ZN(n661) );
  XNOR2_X1 U736 ( .A(KEYINPUT27), .B(n661), .ZN(n662) );
  XNOR2_X1 U737 ( .A(n663), .B(n662), .ZN(G9) );
  XOR2_X1 U738 ( .A(G128), .B(KEYINPUT29), .Z(n666) );
  NAND2_X1 U739 ( .A1(n664), .A2(n669), .ZN(n665) );
  XNOR2_X1 U740 ( .A(n666), .B(n665), .ZN(G30) );
  XNOR2_X1 U741 ( .A(G143), .B(n667), .ZN(G45) );
  NAND2_X1 U742 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U743 ( .A(n670), .B(G146), .ZN(G48) );
  NOR2_X1 U744 ( .A1(n671), .A2(n410), .ZN(n672) );
  XOR2_X1 U745 ( .A(G113), .B(n672), .Z(G15) );
  NOR2_X1 U746 ( .A1(n673), .A2(n410), .ZN(n674) );
  XOR2_X1 U747 ( .A(KEYINPUT112), .B(n674), .Z(n675) );
  XNOR2_X1 U748 ( .A(G116), .B(n675), .ZN(G18) );
  XNOR2_X1 U749 ( .A(G125), .B(n676), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n677), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U751 ( .A(G134), .B(KEYINPUT113), .Z(n678) );
  XNOR2_X1 U752 ( .A(n679), .B(n678), .ZN(G36) );
  XOR2_X1 U753 ( .A(G140), .B(n680), .Z(G42) );
  BUF_X1 U754 ( .A(n681), .Z(n682) );
  NOR2_X1 U755 ( .A1(n684), .A2(n683), .ZN(n685) );
  NOR2_X1 U756 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U757 ( .A(n687), .B(KEYINPUT116), .ZN(n691) );
  NOR2_X1 U758 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U759 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U760 ( .A(KEYINPUT117), .B(n692), .Z(n693) );
  NOR2_X1 U761 ( .A1(n394), .A2(n693), .ZN(n694) );
  XNOR2_X1 U762 ( .A(n694), .B(KEYINPUT118), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n358), .A2(n695), .ZN(n696) );
  XNOR2_X1 U764 ( .A(KEYINPUT49), .B(n696), .ZN(n704) );
  NOR2_X1 U765 ( .A1(n698), .A2(n435), .ZN(n700) );
  XNOR2_X1 U766 ( .A(KEYINPUT50), .B(KEYINPUT114), .ZN(n699) );
  XNOR2_X1 U767 ( .A(n700), .B(n699), .ZN(n702) );
  NOR2_X1 U768 ( .A1(n702), .A2(n701), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n704), .A2(n703), .ZN(n705) );
  NAND2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n708) );
  XOR2_X1 U771 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n707) );
  XNOR2_X1 U772 ( .A(n708), .B(n707), .ZN(n709) );
  NOR2_X1 U773 ( .A1(n719), .A2(n709), .ZN(n710) );
  NOR2_X1 U774 ( .A1(n711), .A2(n710), .ZN(n712) );
  XNOR2_X1 U775 ( .A(n712), .B(KEYINPUT119), .ZN(n713) );
  XNOR2_X1 U776 ( .A(n713), .B(KEYINPUT52), .ZN(n715) );
  NAND2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n716) );
  NAND2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n721) );
  NOR2_X1 U779 ( .A1(n719), .A2(n394), .ZN(n720) );
  NOR2_X1 U780 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X1 U781 ( .A1(n743), .A2(n722), .ZN(n723) );
  XOR2_X1 U782 ( .A(KEYINPUT53), .B(n723), .Z(G75) );
  XNOR2_X1 U783 ( .A(KEYINPUT55), .B(KEYINPUT79), .ZN(n726) );
  XNOR2_X1 U784 ( .A(n408), .B(KEYINPUT54), .ZN(n725) );
  XNOR2_X1 U785 ( .A(n726), .B(n725), .ZN(n728) );
  NAND2_X1 U786 ( .A1(n407), .A2(G210), .ZN(n727) );
  NAND2_X1 U787 ( .A1(n360), .A2(n730), .ZN(n736) );
  XOR2_X1 U788 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n732) );
  XNOR2_X1 U789 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n731) );
  XOR2_X1 U790 ( .A(n732), .B(n731), .Z(n733) );
  NAND2_X1 U791 ( .A1(G478), .A2(n738), .ZN(n739) );
  XNOR2_X1 U792 ( .A(n740), .B(n739), .ZN(n741) );
  NOR2_X1 U793 ( .A1(n742), .A2(n741), .ZN(G63) );
  NAND2_X1 U794 ( .A1(G953), .A2(G224), .ZN(n744) );
  XNOR2_X1 U795 ( .A(KEYINPUT61), .B(n744), .ZN(n745) );
  NAND2_X1 U796 ( .A1(n745), .A2(G898), .ZN(n746) );
  NAND2_X1 U797 ( .A1(n747), .A2(n746), .ZN(n753) );
  XNOR2_X1 U798 ( .A(G101), .B(n748), .ZN(n749) );
  NOR2_X1 U799 ( .A1(n751), .A2(n750), .ZN(n752) );
  XNOR2_X1 U800 ( .A(n753), .B(n752), .ZN(G69) );
  XNOR2_X1 U801 ( .A(n754), .B(KEYINPUT4), .ZN(n756) );
  XNOR2_X1 U802 ( .A(n756), .B(n755), .ZN(n761) );
  INV_X1 U803 ( .A(n761), .ZN(n758) );
  XNOR2_X1 U804 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U805 ( .A1(G953), .A2(n759), .ZN(n760) );
  XNOR2_X1 U806 ( .A(KEYINPUT125), .B(n760), .ZN(n766) );
  XNOR2_X1 U807 ( .A(G227), .B(n761), .ZN(n762) );
  NAND2_X1 U808 ( .A1(n762), .A2(G900), .ZN(n763) );
  XNOR2_X1 U809 ( .A(KEYINPUT126), .B(n763), .ZN(n764) );
  NAND2_X1 U810 ( .A1(n764), .A2(G953), .ZN(n765) );
  NAND2_X1 U811 ( .A1(n766), .A2(n765), .ZN(G72) );
  XNOR2_X1 U812 ( .A(G122), .B(n767), .ZN(G24) );
  XOR2_X1 U813 ( .A(G119), .B(n355), .Z(n769) );
  XNOR2_X1 U814 ( .A(KEYINPUT127), .B(n769), .ZN(G21) );
  XNOR2_X1 U815 ( .A(G110), .B(n770), .ZN(G12) );
  XOR2_X1 U816 ( .A(G131), .B(n771), .Z(G33) );
  XOR2_X1 U817 ( .A(G137), .B(n772), .Z(G39) );
endmodule

