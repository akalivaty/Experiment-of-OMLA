//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 0 0 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:07 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n533, new_n534, new_n535,
    new_n536, new_n537, new_n538, new_n540, new_n541, new_n543, new_n544,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n565, new_n566, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n599, new_n600, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n936, new_n937, new_n938,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT64), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  AOI22_X1  g033(.A1(new_n454), .A2(G2106), .B1(G567), .B2(new_n456), .ZN(G319));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2105), .ZN(new_n464));
  NAND4_X1  g039(.A1(new_n461), .A2(new_n463), .A3(G137), .A4(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT65), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n468), .A2(KEYINPUT65), .A3(G137), .A4(new_n464), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n460), .A2(G2105), .ZN(new_n470));
  AOI22_X1  g045(.A1(new_n467), .A2(new_n469), .B1(G101), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g046(.A1(G113), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n461), .A2(new_n463), .ZN(new_n473));
  INV_X1    g048(.A(G125), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n472), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n473), .A2(new_n464), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n473), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  NOR2_X1   g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI21_X1  g058(.A(G2104), .B1(new_n464), .B2(G112), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n480), .B(new_n482), .C1(new_n483), .C2(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND4_X1  g061(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n464), .ZN(new_n487));
  XOR2_X1   g062(.A(KEYINPUT66), .B(KEYINPUT4), .Z(new_n488));
  AND2_X1   g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AND3_X1   g064(.A1(KEYINPUT66), .A2(KEYINPUT4), .A3(G138), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n490), .A2(new_n461), .A3(new_n463), .ZN(new_n491));
  NAND2_X1  g066(.A1(G102), .A2(G2104), .ZN(new_n492));
  AOI21_X1  g067(.A(G2105), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n461), .A2(new_n463), .A3(G126), .ZN(new_n494));
  NAND2_X1  g069(.A1(G114), .A2(G2104), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n464), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NOR3_X1   g071(.A1(new_n489), .A2(new_n493), .A3(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT5), .ZN(new_n498));
  NOR2_X1   g073(.A1(new_n498), .A2(G543), .ZN(new_n499));
  INV_X1    g074(.A(G543), .ZN(new_n500));
  OAI21_X1  g075(.A(KEYINPUT67), .B1(new_n500), .B2(KEYINPUT5), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT67), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(new_n498), .A3(G543), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n499), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OR2_X1    g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  XNOR2_X1  g082(.A(KEYINPUT6), .B(G651), .ZN(new_n508));
  AND2_X1   g083(.A1(new_n504), .A2(new_n508), .ZN(new_n509));
  AND2_X1   g084(.A1(new_n508), .A2(G543), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n509), .A2(G88), .B1(G50), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(G303));
  INV_X1    g087(.A(G303), .ZN(G166));
  NAND2_X1  g088(.A1(new_n509), .A2(G89), .ZN(new_n514));
  AND2_X1   g089(.A1(G63), .A2(G651), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n510), .A2(G51), .B1(new_n504), .B2(new_n515), .ZN(new_n516));
  XOR2_X1   g091(.A(KEYINPUT68), .B(KEYINPUT7), .Z(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n514), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(KEYINPUT69), .ZN(new_n521));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n514), .A2(new_n522), .A3(new_n516), .A4(new_n519), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n521), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n504), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n506), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n504), .A2(new_n508), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  INV_X1    g103(.A(G52), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(G543), .ZN(new_n530));
  OAI22_X1  g105(.A1(new_n527), .A2(new_n528), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n526), .A2(new_n531), .ZN(G171));
  AOI22_X1  g107(.A1(new_n504), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n533), .A2(new_n506), .ZN(new_n534));
  XNOR2_X1  g109(.A(KEYINPUT70), .B(G81), .ZN(new_n535));
  INV_X1    g110(.A(G43), .ZN(new_n536));
  OAI22_X1  g111(.A1(new_n527), .A2(new_n535), .B1(new_n536), .B2(new_n530), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  AND3_X1   g114(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G36), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT71), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n540), .A2(new_n544), .ZN(G188));
  INV_X1    g120(.A(KEYINPUT9), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(KEYINPUT72), .ZN(new_n547));
  AOI21_X1  g122(.A(new_n547), .B1(new_n510), .B2(G53), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n504), .A2(G65), .ZN(new_n549));
  NAND2_X1  g124(.A1(G78), .A2(G543), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g126(.A(new_n548), .B1(G651), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n509), .A2(G91), .ZN(new_n553));
  OR2_X1    g128(.A1(new_n546), .A2(KEYINPUT72), .ZN(new_n554));
  NAND4_X1  g129(.A1(new_n510), .A2(G53), .A3(new_n547), .A4(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n552), .A2(new_n553), .A3(new_n555), .ZN(G299));
  INV_X1    g131(.A(G171), .ZN(G301));
  AND2_X1   g132(.A1(new_n521), .A2(new_n523), .ZN(G286));
  NAND2_X1  g133(.A1(new_n510), .A2(G49), .ZN(new_n559));
  OAI21_X1  g134(.A(G651), .B1(new_n504), .B2(G74), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n504), .A2(G87), .A3(new_n508), .ZN(new_n561));
  NAND3_X1  g136(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n562));
  INV_X1    g137(.A(KEYINPUT73), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n562), .B(new_n563), .ZN(G288));
  AND2_X1   g139(.A1(new_n504), .A2(G61), .ZN(new_n565));
  AND2_X1   g140(.A1(G73), .A2(G543), .ZN(new_n566));
  OAI211_X1 g141(.A(KEYINPUT74), .B(G651), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n568));
  AOI21_X1  g143(.A(new_n566), .B1(new_n504), .B2(G61), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n569), .B2(new_n506), .ZN(new_n570));
  AND2_X1   g145(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(G86), .ZN(new_n572));
  INV_X1    g147(.A(G48), .ZN(new_n573));
  OAI22_X1  g148(.A1(new_n527), .A2(new_n572), .B1(new_n573), .B2(new_n530), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  AND2_X1   g150(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  INV_X1    g151(.A(new_n576), .ZN(G305));
  AOI22_X1  g152(.A1(new_n509), .A2(G85), .B1(G47), .B2(new_n510), .ZN(new_n578));
  INV_X1    g153(.A(KEYINPUT75), .ZN(new_n579));
  XNOR2_X1  g154(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n504), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n581));
  OR2_X1    g156(.A1(new_n581), .A2(new_n506), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n580), .A2(new_n582), .ZN(G290));
  NAND2_X1  g158(.A1(G301), .A2(G868), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT10), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n509), .A2(new_n585), .A3(G92), .ZN(new_n586));
  INV_X1    g161(.A(G92), .ZN(new_n587));
  OAI21_X1  g162(.A(KEYINPUT10), .B1(new_n527), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n510), .A2(G54), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n504), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n506), .ZN(new_n592));
  OR2_X1    g167(.A1(new_n589), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n593), .A2(KEYINPUT76), .ZN(new_n594));
  OR3_X1    g169(.A1(new_n589), .A2(KEYINPUT76), .A3(new_n592), .ZN(new_n595));
  AND2_X1   g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n584), .B1(new_n596), .B2(G868), .ZN(G284));
  OAI21_X1  g172(.A(new_n584), .B1(new_n596), .B2(G868), .ZN(G321));
  INV_X1    g173(.A(G868), .ZN(new_n599));
  NAND2_X1  g174(.A1(G299), .A2(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G297));
  OAI21_X1  g176(.A(new_n600), .B1(G168), .B2(new_n599), .ZN(G280));
  INV_X1    g177(.A(G559), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n596), .B1(new_n603), .B2(G860), .ZN(new_n604));
  XNOR2_X1  g179(.A(new_n604), .B(KEYINPUT77), .ZN(G148));
  NAND3_X1  g180(.A1(new_n594), .A2(new_n603), .A3(new_n595), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(G868), .ZN(new_n607));
  OAI211_X1 g182(.A(new_n607), .B(KEYINPUT78), .C1(G868), .C2(new_n538), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n608), .B1(KEYINPUT78), .B2(new_n607), .ZN(new_n609));
  XNOR2_X1  g184(.A(new_n609), .B(KEYINPUT79), .ZN(G323));
  XNOR2_X1  g185(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g186(.A1(new_n468), .A2(new_n470), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT12), .ZN(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT13), .ZN(new_n614));
  XNOR2_X1  g189(.A(KEYINPUT80), .B(G2100), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  NOR2_X1   g191(.A1(new_n464), .A2(G111), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(KEYINPUT81), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n618), .B(G2104), .C1(G99), .C2(G2105), .ZN(new_n619));
  AOI22_X1  g194(.A1(G123), .A2(new_n479), .B1(new_n481), .B2(G135), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n616), .A2(new_n622), .ZN(G156));
  XNOR2_X1  g198(.A(KEYINPUT15), .B(G2435), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2438), .ZN(new_n625));
  XOR2_X1   g200(.A(G2427), .B(G2430), .Z(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n628));
  NAND2_X1  g203(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT82), .B(KEYINPUT16), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XOR2_X1   g206(.A(G2443), .B(G2446), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT83), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2451), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n631), .B(new_n635), .ZN(new_n636));
  XOR2_X1   g211(.A(G1341), .B(G1348), .Z(new_n637));
  NOR2_X1   g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(KEYINPUT85), .ZN(new_n639));
  INV_X1    g214(.A(G14), .ZN(new_n640));
  AOI21_X1  g215(.A(new_n640), .B1(new_n636), .B2(new_n637), .ZN(new_n641));
  AND2_X1   g216(.A1(new_n639), .A2(new_n641), .ZN(G401));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT86), .ZN(new_n644));
  XOR2_X1   g219(.A(G2072), .B(G2078), .Z(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g222(.A1(new_n644), .A2(new_n645), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT18), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n644), .A2(new_n645), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(KEYINPUT17), .ZN(new_n651));
  OAI211_X1 g226(.A(new_n650), .B(new_n647), .C1(new_n644), .C2(new_n651), .ZN(new_n652));
  NAND3_X1  g227(.A1(new_n644), .A2(new_n651), .A3(new_n646), .ZN(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT87), .B(G2096), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n654), .B(new_n656), .ZN(G227));
  XNOR2_X1  g232(.A(G1971), .B(G1976), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT19), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XOR2_X1   g235(.A(G1956), .B(G2474), .Z(new_n661));
  XOR2_X1   g236(.A(G1961), .B(G1966), .Z(new_n662));
  NOR2_X1   g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n660), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g239(.A(new_n664), .B(KEYINPUT88), .Z(new_n665));
  NAND2_X1  g240(.A1(new_n661), .A2(new_n662), .ZN(new_n666));
  INV_X1    g241(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n660), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT20), .ZN(new_n669));
  OR3_X1    g244(.A1(new_n660), .A2(new_n663), .A3(new_n667), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n665), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  XOR2_X1   g246(.A(KEYINPUT89), .B(G1986), .Z(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT90), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n671), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(G1996), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1991), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n674), .B(new_n678), .ZN(G229));
  NOR2_X1   g254(.A1(G29), .A2(G32), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n481), .A2(G141), .ZN(new_n681));
  XOR2_X1   g256(.A(new_n681), .B(KEYINPUT95), .Z(new_n682));
  AND2_X1   g257(.A1(new_n470), .A2(G105), .ZN(new_n683));
  NAND3_X1  g258(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT26), .ZN(new_n685));
  AOI211_X1 g260(.A(new_n683), .B(new_n685), .C1(G129), .C2(new_n479), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  INV_X1    g262(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n680), .B1(new_n688), .B2(G29), .ZN(new_n689));
  XOR2_X1   g264(.A(KEYINPUT27), .B(G1996), .Z(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(G34), .ZN(new_n693));
  INV_X1    g268(.A(G29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(new_n477), .B2(new_n694), .ZN(new_n696));
  INV_X1    g271(.A(G2084), .ZN(new_n697));
  NAND2_X1  g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n694), .A2(G35), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n699), .B1(G162), .B2(new_n694), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(KEYINPUT29), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n698), .B1(new_n701), .B2(G2090), .ZN(new_n702));
  NAND2_X1  g277(.A1(G164), .A2(G29), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n703), .B1(G27), .B2(G29), .ZN(new_n704));
  INV_X1    g279(.A(G2078), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT30), .B(G28), .Z(new_n707));
  NAND2_X1  g282(.A1(G171), .A2(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n708), .B1(G5), .B2(G16), .ZN(new_n709));
  INV_X1    g284(.A(G1961), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n706), .B1(G29), .B2(new_n707), .C1(new_n709), .C2(new_n710), .ZN(new_n711));
  NOR3_X1   g286(.A1(new_n691), .A2(new_n702), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g287(.A1(new_n619), .A2(new_n620), .A3(G29), .ZN(new_n713));
  INV_X1    g288(.A(G16), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n714), .A2(KEYINPUT23), .A3(G20), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT23), .ZN(new_n716));
  INV_X1    g291(.A(G20), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n716), .B1(new_n717), .B2(G16), .ZN(new_n718));
  INV_X1    g293(.A(G53), .ZN(new_n719));
  OAI211_X1 g294(.A(KEYINPUT72), .B(new_n546), .C1(new_n530), .C2(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(G91), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n504), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n722));
  OAI221_X1 g297(.A(new_n720), .B1(new_n527), .B2(new_n721), .C1(new_n722), .C2(new_n506), .ZN(new_n723));
  INV_X1    g298(.A(new_n555), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n715), .B(new_n718), .C1(new_n725), .C2(new_n714), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT98), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT97), .B(G1956), .Z(new_n728));
  OR2_X1    g303(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n727), .A2(new_n728), .ZN(new_n730));
  NAND4_X1  g305(.A1(new_n712), .A2(new_n713), .A3(new_n729), .A4(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G26), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n479), .A2(G128), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n481), .A2(G140), .ZN(new_n735));
  NOR2_X1   g310(.A1(G104), .A2(G2105), .ZN(new_n736));
  OAI21_X1  g311(.A(G2104), .B1(new_n464), .B2(G116), .ZN(new_n737));
  OAI211_X1 g312(.A(new_n734), .B(new_n735), .C1(new_n736), .C2(new_n737), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n733), .B1(new_n738), .B2(G29), .ZN(new_n739));
  MUX2_X1   g314(.A(new_n733), .B(new_n739), .S(KEYINPUT28), .Z(new_n740));
  XOR2_X1   g315(.A(KEYINPUT91), .B(G2067), .Z(new_n741));
  XOR2_X1   g316(.A(new_n740), .B(new_n741), .Z(new_n742));
  AND2_X1   g317(.A1(new_n709), .A2(new_n710), .ZN(new_n743));
  NOR2_X1   g318(.A1(new_n696), .A2(new_n697), .ZN(new_n744));
  NOR2_X1   g319(.A1(G16), .A2(G19), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(new_n538), .B2(G16), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n744), .B1(G1341), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G1341), .B2(new_n746), .ZN(new_n748));
  OR3_X1    g323(.A1(new_n742), .A2(new_n743), .A3(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n714), .A2(G4), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n596), .B2(new_n714), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n751), .A2(G1348), .ZN(new_n752));
  NOR2_X1   g327(.A1(G16), .A2(G21), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(G168), .B2(G16), .ZN(new_n754));
  INV_X1    g329(.A(G1966), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT92), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G29), .B2(G33), .ZN(new_n759));
  OR3_X1    g334(.A1(new_n758), .A2(G29), .A3(G33), .ZN(new_n760));
  NAND2_X1  g335(.A1(G115), .A2(G2104), .ZN(new_n761));
  INV_X1    g336(.A(G127), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n761), .B1(new_n473), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n763), .A2(G2105), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(KEYINPUT93), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n481), .A2(G139), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n470), .A2(G103), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n759), .B(new_n760), .C1(new_n769), .C2(new_n694), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(G2072), .ZN(new_n771));
  XNOR2_X1  g346(.A(KEYINPUT31), .B(G11), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NOR4_X1   g348(.A1(new_n731), .A2(new_n749), .A3(new_n757), .A4(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n701), .A2(G2090), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT96), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n714), .A2(G6), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n576), .B2(new_n714), .ZN(new_n778));
  XOR2_X1   g353(.A(KEYINPUT32), .B(G1981), .Z(new_n779));
  XNOR2_X1  g354(.A(new_n778), .B(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n714), .A2(G22), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G166), .B2(new_n714), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1971), .ZN(new_n783));
  NOR2_X1   g358(.A1(G16), .A2(G23), .ZN(new_n784));
  AND3_X1   g359(.A1(new_n559), .A2(new_n560), .A3(new_n561), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n784), .B1(new_n785), .B2(G16), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT33), .B(G1976), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n783), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n780), .A2(new_n789), .ZN(new_n790));
  INV_X1    g365(.A(KEYINPUT34), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n780), .A2(new_n789), .A3(KEYINPUT34), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT36), .ZN(new_n795));
  AND2_X1   g370(.A1(new_n714), .A2(G24), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G290), .B2(G16), .ZN(new_n797));
  INV_X1    g372(.A(G1986), .ZN(new_n798));
  AND2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g374(.A1(new_n797), .A2(new_n798), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n694), .A2(G25), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n479), .A2(G119), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n481), .A2(G131), .ZN(new_n803));
  OR2_X1    g378(.A1(G95), .A2(G2105), .ZN(new_n804));
  OAI211_X1 g379(.A(new_n804), .B(G2104), .C1(G107), .C2(new_n464), .ZN(new_n805));
  AND3_X1   g380(.A1(new_n802), .A2(new_n803), .A3(new_n805), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n801), .B1(new_n806), .B2(new_n694), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT35), .B(G1991), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n807), .B(new_n808), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n799), .A2(new_n800), .A3(new_n809), .ZN(new_n810));
  AND3_X1   g385(.A1(new_n794), .A2(new_n795), .A3(new_n810), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n795), .B1(new_n794), .B2(new_n810), .ZN(new_n812));
  OAI211_X1 g387(.A(new_n774), .B(new_n776), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n704), .A2(new_n705), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n751), .A2(G1348), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(G311));
  INV_X1    g391(.A(G311), .ZN(G150));
  AOI22_X1  g392(.A1(new_n504), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n506), .ZN(new_n819));
  XOR2_X1   g394(.A(KEYINPUT99), .B(G93), .Z(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n527), .A2(new_n820), .B1(new_n821), .B2(new_n530), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n824), .A2(G860), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(KEYINPUT37), .Z(new_n826));
  NAND2_X1  g401(.A1(new_n596), .A2(G559), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n538), .B1(new_n819), .B2(new_n822), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n823), .B1(new_n534), .B2(new_n537), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n827), .B(new_n832), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n826), .B1(new_n833), .B2(G860), .ZN(G145));
  XNOR2_X1  g409(.A(new_n621), .B(new_n477), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(G162), .ZN(new_n836));
  INV_X1    g411(.A(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(G164), .B(new_n738), .ZN(new_n838));
  XOR2_X1   g413(.A(new_n838), .B(new_n769), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(new_n687), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT101), .ZN(new_n841));
  INV_X1    g416(.A(new_n806), .ZN(new_n842));
  INV_X1    g417(.A(new_n613), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT100), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n481), .A2(new_n844), .A3(G142), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n468), .A2(new_n464), .ZN(new_n846));
  INV_X1    g421(.A(G142), .ZN(new_n847));
  OAI21_X1  g422(.A(KEYINPUT100), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n479), .A2(G130), .ZN(new_n849));
  OR2_X1    g424(.A1(G106), .A2(G2105), .ZN(new_n850));
  OAI211_X1 g425(.A(new_n850), .B(G2104), .C1(G118), .C2(new_n464), .ZN(new_n851));
  NAND4_X1  g426(.A1(new_n845), .A2(new_n848), .A3(new_n849), .A4(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n843), .A2(new_n852), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n842), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR3_X1   g431(.A1(new_n853), .A2(new_n854), .A3(new_n842), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n841), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n852), .B(new_n613), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(new_n806), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n860), .A2(KEYINPUT101), .A3(new_n855), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n838), .B(new_n769), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(new_n688), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n840), .A2(new_n862), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n862), .B1(new_n840), .B2(new_n864), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n837), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n840), .A2(new_n864), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n856), .A2(new_n857), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n840), .A2(new_n862), .A3(new_n864), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(new_n871), .A3(new_n836), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n867), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(KEYINPUT102), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g451(.A1(new_n867), .A2(new_n872), .A3(KEYINPUT102), .A4(new_n873), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g454(.A(KEYINPUT106), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT42), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(G303), .B(new_n562), .ZN(new_n883));
  AND2_X1   g458(.A1(new_n883), .A2(G290), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n883), .A2(G290), .ZN(new_n885));
  OAI21_X1  g460(.A(G305), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n883), .A2(G290), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n883), .A2(G290), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n576), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n886), .A2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n880), .A2(new_n881), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n882), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n882), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n893), .B1(new_n886), .B2(new_n889), .ZN(new_n894));
  OAI21_X1  g469(.A(KEYINPUT107), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n830), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n606), .B(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT103), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n723), .B2(new_n724), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n552), .A2(KEYINPUT103), .A3(new_n553), .A4(new_n555), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n593), .A2(new_n899), .A3(new_n900), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n589), .A2(new_n592), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n725), .A2(new_n902), .A3(KEYINPUT103), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT104), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n903), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n897), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(KEYINPUT105), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT41), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n901), .A2(new_n910), .A3(new_n903), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n910), .B1(new_n901), .B2(new_n903), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n909), .B1(new_n914), .B2(new_n897), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n890), .A2(new_n882), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT107), .ZN(new_n917));
  AOI22_X1  g492(.A1(new_n886), .A2(new_n889), .B1(new_n880), .B2(new_n881), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n916), .B(new_n917), .C1(new_n918), .C2(new_n882), .ZN(new_n919));
  NOR2_X1   g494(.A1(new_n897), .A2(new_n914), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(KEYINPUT105), .ZN(new_n921));
  NAND4_X1  g496(.A1(new_n895), .A2(new_n915), .A3(new_n919), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n916), .B1(new_n918), .B2(new_n882), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n920), .B1(KEYINPUT105), .B2(new_n908), .ZN(new_n924));
  INV_X1    g499(.A(new_n921), .ZN(new_n925));
  OAI211_X1 g500(.A(KEYINPUT107), .B(new_n923), .C1(new_n924), .C2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n922), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(G868), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT108), .ZN(new_n929));
  NOR2_X1   g504(.A1(new_n824), .A2(G868), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g506(.A1(new_n928), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n599), .B1(new_n922), .B2(new_n926), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT108), .B1(new_n933), .B2(new_n930), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n932), .A2(new_n934), .ZN(G295));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n928), .A2(new_n936), .A3(new_n931), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT109), .B1(new_n933), .B2(new_n930), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n937), .A2(new_n938), .ZN(G331));
  NAND2_X1  g514(.A1(new_n830), .A2(G286), .ZN(new_n940));
  NAND3_X1  g515(.A1(G168), .A2(new_n828), .A3(new_n829), .ZN(new_n941));
  AND3_X1   g516(.A1(new_n940), .A2(G171), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(G171), .B1(new_n940), .B2(new_n941), .ZN(new_n943));
  INV_X1    g518(.A(new_n906), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n942), .A2(new_n943), .B1(new_n944), .B2(new_n904), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT111), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(new_n913), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT110), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n948), .A2(new_n949), .A3(new_n911), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n940), .A2(G171), .A3(new_n941), .ZN(new_n951));
  INV_X1    g526(.A(new_n941), .ZN(new_n952));
  AOI21_X1  g527(.A(G168), .B1(new_n828), .B2(new_n829), .ZN(new_n953));
  OAI21_X1  g528(.A(G301), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n913), .A2(KEYINPUT110), .ZN(new_n955));
  NAND4_X1  g530(.A1(new_n950), .A2(new_n951), .A3(new_n954), .A4(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n907), .B(KEYINPUT111), .C1(new_n942), .C2(new_n943), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n947), .A2(new_n956), .A3(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n890), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n903), .B(new_n901), .C1(new_n942), .C2(new_n943), .ZN(new_n961));
  OAI211_X1 g536(.A(new_n954), .B(new_n951), .C1(new_n912), .C2(new_n913), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n961), .A2(new_n890), .A3(new_n962), .ZN(new_n963));
  AND2_X1   g538(.A1(new_n963), .A2(new_n873), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT43), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n960), .A2(new_n964), .A3(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT112), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n961), .A2(new_n962), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(new_n959), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n873), .A3(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT112), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n960), .A2(new_n964), .A3(new_n972), .A4(new_n965), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n967), .A2(new_n971), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT44), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n960), .A2(new_n964), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n975), .B1(new_n977), .B2(KEYINPUT43), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT113), .ZN(new_n979));
  OR3_X1    g554(.A1(new_n970), .A2(new_n979), .A3(KEYINPUT43), .ZN(new_n980));
  OAI21_X1  g555(.A(new_n979), .B1(new_n970), .B2(KEYINPUT43), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n976), .A2(new_n982), .ZN(G397));
  NOR2_X1   g558(.A1(new_n738), .A2(G2067), .ZN(new_n984));
  INV_X1    g559(.A(G1996), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n688), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(G2067), .ZN(new_n987));
  XNOR2_X1  g562(.A(new_n738), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n687), .A2(G1996), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n986), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(new_n990), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n842), .A2(new_n808), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n984), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G40), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n475), .B2(G2105), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n471), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT114), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n471), .A2(new_n995), .A3(KEYINPUT114), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1001), .B1(G164), .B2(G1384), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g578(.A(new_n1003), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n993), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n1004), .B1(new_n688), .B2(new_n988), .ZN(new_n1006));
  AND3_X1   g581(.A1(new_n1003), .A2(KEYINPUT46), .A3(new_n985), .ZN(new_n1007));
  AOI21_X1  g582(.A(KEYINPUT46), .B1(new_n1003), .B2(new_n985), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n1009), .B(KEYINPUT47), .ZN(new_n1010));
  INV_X1    g585(.A(new_n808), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n991), .B1(new_n1011), .B2(new_n806), .ZN(new_n1012));
  OAI21_X1  g587(.A(new_n1003), .B1(new_n1012), .B2(new_n992), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n580), .A2(new_n798), .A3(new_n582), .ZN(new_n1014));
  NOR2_X1   g589(.A1(new_n1004), .A2(new_n1014), .ZN(new_n1015));
  XOR2_X1   g590(.A(new_n1015), .B(KEYINPUT48), .Z(new_n1016));
  AOI211_X1 g591(.A(new_n1005), .B(new_n1010), .C1(new_n1013), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G8), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n491), .A2(new_n492), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(new_n464), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n494), .A2(new_n495), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n1021), .A2(G2105), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n487), .A2(new_n488), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1022), .A3(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(G1384), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1024), .A2(KEYINPUT45), .A3(new_n1025), .ZN(new_n1026));
  NAND4_X1  g601(.A1(new_n1002), .A2(new_n998), .A3(new_n999), .A4(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(G1971), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1030), .B1(G164), .B2(G1384), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1024), .A2(KEYINPUT50), .A3(new_n1025), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n471), .A2(KEYINPUT114), .A3(new_n995), .ZN(new_n1034));
  AOI21_X1  g609(.A(KEYINPUT114), .B1(new_n471), .B2(new_n995), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g611(.A(G2090), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n1033), .A2(new_n1036), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1018), .B1(new_n1029), .B2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(new_n1018), .B1(new_n507), .B2(new_n511), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT115), .ZN(new_n1041));
  NOR2_X1   g616(.A1(new_n1041), .A2(KEYINPUT55), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT115), .B(KEYINPUT55), .Z(new_n1044));
  OAI21_X1  g619(.A(new_n1043), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  XNOR2_X1  g621(.A(new_n1039), .B(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT52), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n493), .A2(new_n496), .ZN(new_n1049));
  AOI21_X1  g624(.A(G1384), .B1(new_n1049), .B2(new_n1023), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n998), .A2(new_n999), .A3(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  INV_X1    g627(.A(G1976), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1052), .B1(new_n562), .B2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n785), .A2(KEYINPUT116), .A3(G1976), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1051), .A2(new_n1054), .A3(G8), .A4(new_n1055), .ZN(new_n1056));
  NAND2_X1  g631(.A1(G288), .A2(new_n1053), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1048), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1018), .B1(new_n1036), .B2(new_n1050), .ZN(new_n1059));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1059), .A2(new_n1060), .A3(new_n1054), .A4(new_n1055), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1058), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1981), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n575), .A2(new_n567), .A3(new_n1063), .A4(new_n570), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n569), .A2(new_n506), .ZN(new_n1065));
  OAI21_X1  g640(.A(G1981), .B1(new_n1065), .B2(new_n574), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1067), .A2(KEYINPUT118), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT49), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1070), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1069), .A2(new_n1059), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g647(.A(new_n1056), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n1073), .A2(new_n1060), .A3(new_n1048), .A4(new_n1057), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n1062), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT127), .B1(new_n1047), .B2(new_n1075), .ZN(new_n1076));
  AND3_X1   g651(.A1(new_n1062), .A2(new_n1072), .A3(new_n1074), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT127), .ZN(new_n1078));
  XNOR2_X1  g653(.A(new_n1039), .B(new_n1045), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1077), .A2(new_n1078), .A3(new_n1079), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1076), .A2(new_n1080), .ZN(new_n1081));
  AND3_X1   g656(.A1(new_n1024), .A2(KEYINPUT50), .A3(new_n1025), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT50), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1083));
  NOR2_X1   g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  OAI21_X1  g659(.A(KEYINPUT122), .B1(new_n1084), .B2(new_n1000), .ZN(new_n1085));
  INV_X1    g660(.A(KEYINPUT122), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1033), .A2(new_n1036), .A3(new_n1086), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n1085), .A2(new_n710), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT53), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1027), .B2(G2078), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1027), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1091), .A2(KEYINPUT53), .A3(new_n705), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1088), .A2(new_n1090), .A3(new_n1092), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1093), .A2(G171), .ZN(new_n1094));
  NOR2_X1   g669(.A1(G168), .A2(new_n1018), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT126), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT51), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1027), .A2(new_n755), .ZN(new_n1098));
  XNOR2_X1  g673(.A(KEYINPUT119), .B(G2084), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1033), .A2(new_n1036), .A3(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1018), .B1(new_n1098), .B2(new_n1100), .ZN(new_n1101));
  OR3_X1    g676(.A1(new_n1097), .A2(new_n1101), .A3(new_n1095), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(G286), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1097), .B1(new_n1101), .B2(new_n1095), .ZN(new_n1104));
  NAND3_X1  g679(.A1(new_n1102), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(KEYINPUT62), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT62), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1102), .A2(new_n1107), .A3(new_n1103), .A4(new_n1104), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1081), .A2(new_n1094), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(new_n1059), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1111));
  NOR2_X1   g686(.A1(G288), .A2(G1976), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g688(.A(new_n1110), .B1(new_n1113), .B2(new_n1064), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1039), .A2(new_n1046), .ZN(new_n1115));
  OAI211_X1 g690(.A(G168), .B(new_n1101), .C1(new_n1039), .C2(new_n1046), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(KEYINPUT63), .ZN(new_n1117));
  AOI21_X1  g692(.A(new_n1114), .B1(new_n1117), .B2(new_n1077), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT120), .ZN(new_n1119));
  OAI21_X1  g694(.A(KEYINPUT63), .B1(new_n1075), .B2(new_n1116), .ZN(new_n1120));
  AND3_X1   g695(.A1(new_n1118), .A2(new_n1119), .A3(new_n1120), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1119), .B1(new_n1118), .B2(new_n1120), .ZN(new_n1122));
  OAI21_X1  g697(.A(new_n1109), .B1(new_n1121), .B2(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(G1348), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1085), .A2(new_n1124), .A3(new_n1087), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT121), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1036), .A2(new_n1126), .A3(new_n1050), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1051), .A2(KEYINPUT121), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1127), .A2(new_n1128), .A3(new_n987), .ZN(new_n1129));
  AOI21_X1  g704(.A(KEYINPUT123), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1125), .A2(KEYINPUT123), .A3(new_n1129), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1131), .A2(new_n596), .A3(new_n1132), .ZN(new_n1133));
  AND3_X1   g708(.A1(new_n1125), .A2(KEYINPUT123), .A3(new_n1129), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT60), .ZN(new_n1135));
  NOR3_X1   g710(.A1(new_n1134), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  OAI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(new_n596), .ZN(new_n1137));
  XOR2_X1   g712(.A(KEYINPUT125), .B(KEYINPUT60), .Z(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1137), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(new_n725), .B(KEYINPUT57), .ZN(new_n1141));
  XNOR2_X1  g716(.A(KEYINPUT56), .B(G2072), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1091), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1956), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1084), .B2(new_n1000), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1143), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT124), .ZN(new_n1147));
  INV_X1    g722(.A(KEYINPUT124), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1148), .A3(new_n1145), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1141), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n1151));
  AND3_X1   g726(.A1(new_n1143), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1152));
  NOR3_X1   g727(.A1(new_n1150), .A2(new_n1151), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1141), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1151), .B1(new_n1152), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT59), .ZN(new_n1156));
  XOR2_X1   g731(.A(KEYINPUT58), .B(G1341), .Z(new_n1157));
  INV_X1    g732(.A(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1158), .B1(new_n1127), .B2(new_n1128), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1027), .A2(G1996), .ZN(new_n1160));
  OR2_X1    g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1156), .B1(new_n1161), .B2(new_n538), .ZN(new_n1162));
  OAI211_X1 g737(.A(new_n1156), .B(new_n538), .C1(new_n1159), .C2(new_n1160), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1155), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  NOR2_X1   g740(.A1(new_n1153), .A2(new_n1165), .ZN(new_n1166));
  OAI211_X1 g741(.A(new_n1133), .B(new_n1138), .C1(new_n1136), .C2(new_n596), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1140), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1133), .A2(new_n1152), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n1150), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1002), .A2(new_n1026), .ZN(new_n1172));
  OR4_X1    g747(.A1(new_n1089), .A2(new_n1172), .A3(G2078), .A4(new_n996), .ZN(new_n1173));
  XNOR2_X1  g748(.A(G171), .B(KEYINPUT54), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1173), .A2(new_n1088), .A3(new_n1174), .A4(new_n1090), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1174), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1093), .A2(new_n1176), .ZN(new_n1177));
  AND4_X1   g752(.A1(new_n1081), .A2(new_n1175), .A3(new_n1177), .A4(new_n1105), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1123), .B1(new_n1171), .B2(new_n1178), .ZN(new_n1179));
  AOI211_X1 g754(.A(new_n992), .B(new_n1012), .C1(G1986), .C2(G290), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n1004), .B1(new_n1180), .B2(new_n1014), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1017), .B1(new_n1179), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g757(.A(G227), .B(G229), .C1(new_n876), .C2(new_n877), .ZN(new_n1184));
  INV_X1    g758(.A(G319), .ZN(new_n1185));
  NOR2_X1   g759(.A1(G401), .A2(new_n1185), .ZN(new_n1186));
  AND3_X1   g760(.A1(new_n1184), .A2(new_n974), .A3(new_n1186), .ZN(G308));
  NAND3_X1  g761(.A1(new_n1184), .A2(new_n974), .A3(new_n1186), .ZN(G225));
endmodule


