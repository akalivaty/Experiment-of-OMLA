//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:37 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n682,
    new_n683, new_n684, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n706,
    new_n707, new_n709, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n717, new_n718, new_n719, new_n720, new_n721, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  XOR2_X1   g000(.A(KEYINPUT9), .B(G234), .Z(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G221), .B1(new_n188), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G125), .ZN(new_n194));
  OR2_X1    g008(.A1(new_n194), .A2(KEYINPUT16), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n192), .A2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(G146), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(G146), .A3(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n198), .A2(new_n199), .ZN(new_n200));
  XOR2_X1   g014(.A(KEYINPUT24), .B(G110), .Z(new_n201));
  XNOR2_X1  g015(.A(G119), .B(G128), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(G119), .ZN(new_n206));
  MUX2_X1   g020(.A(KEYINPUT23), .B(new_n205), .S(new_n206), .Z(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G110), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n200), .A2(new_n203), .A3(new_n208), .ZN(new_n209));
  OAI22_X1  g023(.A1(new_n207), .A2(G110), .B1(new_n202), .B2(new_n201), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n191), .A2(new_n197), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n210), .A2(new_n199), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n212), .ZN(new_n213));
  INV_X1    g027(.A(G953), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(G221), .A3(G234), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT73), .ZN(new_n216));
  XNOR2_X1  g030(.A(KEYINPUT22), .B(G137), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(G902), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n209), .A2(new_n212), .A3(new_n218), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT74), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT25), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G217), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n227), .B1(G234), .B2(new_n221), .ZN(new_n228));
  AND2_X1   g042(.A1(new_n223), .A2(new_n225), .ZN(new_n229));
  OAI21_X1  g043(.A(KEYINPUT74), .B1(new_n223), .B2(new_n225), .ZN(new_n230));
  OAI211_X1 g044(.A(new_n226), .B(new_n228), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n220), .A2(new_n222), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n228), .A2(G902), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n231), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(G469), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT75), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT3), .ZN(new_n238));
  INV_X1    g052(.A(G107), .ZN(new_n239));
  NAND4_X1  g053(.A1(new_n237), .A2(new_n238), .A3(new_n239), .A4(G104), .ZN(new_n240));
  INV_X1    g054(.A(G104), .ZN(new_n241));
  AOI22_X1  g055(.A1(new_n241), .A2(G107), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n242));
  OAI22_X1  g056(.A1(new_n241), .A2(G107), .B1(KEYINPUT75), .B2(KEYINPUT3), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G101), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n240), .A2(new_n242), .A3(new_n243), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT76), .B(G101), .ZN(new_n247));
  AOI21_X1  g061(.A(KEYINPUT77), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  NAND4_X1  g062(.A1(new_n247), .A2(new_n240), .A3(new_n242), .A4(new_n243), .ZN(new_n249));
  INV_X1    g063(.A(KEYINPUT77), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  OAI211_X1 g065(.A(KEYINPUT4), .B(new_n245), .C1(new_n248), .C2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G143), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(G146), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n197), .A2(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  OR3_X1    g070(.A1(KEYINPUT65), .A2(KEYINPUT0), .A3(G128), .ZN(new_n257));
  NAND2_X1  g071(.A1(KEYINPUT0), .A2(G128), .ZN(new_n258));
  OAI21_X1  g072(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n256), .A2(new_n257), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n255), .A3(KEYINPUT0), .A4(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  OR2_X1    g077(.A1(new_n245), .A2(KEYINPUT4), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n252), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n241), .A2(G107), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n239), .A2(G104), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n268), .A2(G101), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n254), .A3(new_n255), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n204), .A2(new_n197), .A3(G143), .ZN(new_n273));
  OAI211_X1 g087(.A(new_n253), .B(G146), .C1(new_n204), .C2(KEYINPUT1), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n270), .B(new_n275), .C1(new_n248), .C2(new_n251), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT10), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT11), .ZN(new_n279));
  INV_X1    g093(.A(G134), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n279), .B1(new_n280), .B2(G137), .ZN(new_n281));
  INV_X1    g095(.A(G137), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT11), .A3(G134), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(G131), .ZN(new_n286));
  INV_X1    g100(.A(G131), .ZN(new_n287));
  NAND4_X1  g101(.A1(new_n281), .A2(new_n283), .A3(new_n287), .A4(new_n284), .ZN(new_n288));
  AND2_X1   g102(.A1(new_n286), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n246), .A2(KEYINPUT77), .A3(new_n247), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n249), .A2(new_n250), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n269), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n275), .A2(KEYINPUT69), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT69), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n272), .A2(new_n294), .A3(new_n273), .A4(new_n274), .ZN(new_n295));
  AOI21_X1  g109(.A(new_n277), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n292), .A2(new_n296), .ZN(new_n297));
  NAND4_X1  g111(.A1(new_n265), .A2(new_n278), .A3(new_n289), .A4(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(G110), .B(G140), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n214), .A2(G227), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n299), .B(new_n300), .Z(new_n301));
  NAND2_X1  g115(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT12), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n270), .B1(new_n248), .B2(new_n251), .ZN(new_n304));
  INV_X1    g118(.A(new_n275), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AOI211_X1 g120(.A(new_n303), .B(new_n289), .C1(new_n306), .C2(new_n276), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n276), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n286), .A2(new_n288), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n303), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n302), .B1(new_n308), .B2(new_n312), .ZN(new_n313));
  AOI22_X1  g127(.A1(new_n276), .A2(new_n277), .B1(new_n292), .B2(new_n296), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(new_n265), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n310), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n301), .B1(new_n316), .B2(new_n298), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n236), .B(new_n221), .C1(new_n313), .C2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(KEYINPUT78), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT12), .B1(new_n309), .B2(new_n310), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n298), .B(new_n301), .C1(new_n320), .C2(new_n307), .ZN(new_n321));
  INV_X1    g135(.A(new_n301), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n314), .A2(new_n289), .A3(new_n265), .ZN(new_n323));
  AOI21_X1  g137(.A(new_n289), .B1(new_n314), .B2(new_n265), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  AOI21_X1  g139(.A(G902), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT78), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n326), .A2(new_n327), .A3(new_n236), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n319), .A2(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n302), .A2(new_n324), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n298), .B1(new_n320), .B2(new_n307), .ZN(new_n331));
  AOI21_X1  g145(.A(new_n330), .B1(new_n322), .B2(new_n331), .ZN(new_n332));
  OAI21_X1  g146(.A(G469), .B1(new_n332), .B2(G902), .ZN(new_n333));
  AOI211_X1 g147(.A(new_n190), .B(new_n235), .C1(new_n329), .C2(new_n333), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT89), .A2(G952), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  NAND2_X1  g150(.A1(KEYINPUT89), .A2(G952), .ZN(new_n337));
  AOI21_X1  g151(.A(G953), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G234), .ZN(new_n339));
  INV_X1    g153(.A(G237), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n338), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  XOR2_X1   g155(.A(KEYINPUT21), .B(G898), .Z(new_n342));
  AOI211_X1 g156(.A(new_n221), .B(new_n214), .C1(G234), .C2(G237), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n341), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(new_n345), .ZN(new_n346));
  OAI21_X1  g160(.A(G214), .B1(G237), .B2(G902), .ZN(new_n347));
  INV_X1    g161(.A(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G116), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n349), .A2(G119), .ZN(new_n350));
  AND2_X1   g164(.A1(new_n349), .A2(G119), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT68), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G116), .B(G119), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT67), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT2), .ZN(new_n358));
  INV_X1    g172(.A(G113), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n357), .B1(new_n358), .B2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(KEYINPUT67), .A2(KEYINPUT2), .A3(G113), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OR2_X1    g176(.A1(KEYINPUT2), .A2(G113), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n356), .A2(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n362), .A2(new_n363), .A3(new_n353), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n252), .A2(new_n264), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n366), .ZN(new_n369));
  XOR2_X1   g183(.A(KEYINPUT79), .B(KEYINPUT5), .Z(new_n370));
  NAND3_X1  g184(.A1(new_n352), .A2(new_n355), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n370), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n359), .B1(new_n372), .B2(new_n350), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n369), .B1(new_n371), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n292), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n368), .A2(new_n375), .ZN(new_n376));
  XOR2_X1   g190(.A(G110), .B(G122), .Z(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n377), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n368), .A2(new_n379), .A3(new_n375), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n378), .A2(KEYINPUT6), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n263), .A2(G125), .ZN(new_n382));
  INV_X1    g196(.A(G125), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n275), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n214), .A2(G224), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n385), .B(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n376), .A2(new_n388), .A3(new_n377), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n381), .A2(new_n387), .A3(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n353), .A2(KEYINPUT5), .ZN(new_n391));
  AND2_X1   g205(.A1(new_n373), .A2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n292), .B1(new_n392), .B2(new_n369), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n304), .A2(new_n374), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n377), .A2(KEYINPUT8), .ZN(new_n395));
  OR2_X1    g209(.A1(new_n377), .A2(KEYINPUT8), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n393), .A2(new_n394), .A3(new_n395), .A4(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n386), .A2(KEYINPUT7), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n382), .A2(new_n398), .A3(new_n384), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n386), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n380), .A2(new_n397), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n390), .A2(new_n221), .A3(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(G210), .B1(G237), .B2(G902), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n390), .A2(new_n221), .A3(new_n403), .A4(new_n401), .ZN(new_n406));
  AOI211_X1 g220(.A(new_n346), .B(new_n348), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G475), .ZN(new_n408));
  XNOR2_X1  g222(.A(G113), .B(G122), .ZN(new_n409));
  XNOR2_X1  g223(.A(new_n409), .B(new_n241), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n410), .A2(KEYINPUT84), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n383), .A2(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n194), .A2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G146), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT80), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n414), .A2(new_n211), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(G237), .A2(G953), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(G143), .A3(G214), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(G143), .B1(new_n417), .B2(G214), .ZN(new_n420));
  OAI211_X1 g234(.A(KEYINPUT18), .B(G131), .C1(new_n419), .C2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n413), .A2(KEYINPUT80), .A3(G146), .ZN(new_n422));
  AND3_X1   g236(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n340), .A2(new_n214), .A3(G214), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n253), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT18), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT81), .B1(new_n426), .B2(new_n287), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(KEYINPUT18), .A3(G131), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n425), .A2(new_n418), .A3(new_n427), .A4(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT82), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n427), .A2(new_n429), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n433), .A2(KEYINPUT82), .A3(new_n425), .A4(new_n418), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n423), .A2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n419), .B2(new_n420), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n425), .A2(new_n287), .A3(new_n418), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  NAND4_X1  g255(.A1(new_n439), .A2(new_n199), .A3(new_n198), .A4(new_n441), .ZN(new_n442));
  AOI21_X1  g256(.A(new_n411), .B1(new_n436), .B2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G902), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n436), .A2(new_n411), .A3(new_n442), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n408), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(KEYINPUT83), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n383), .A2(G140), .ZN(new_n448));
  NOR2_X1   g262(.A1(new_n193), .A2(G125), .ZN(new_n449));
  OAI21_X1  g263(.A(KEYINPUT19), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT19), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n194), .A2(new_n412), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n450), .A2(new_n197), .A3(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n199), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n437), .A2(new_n440), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n423), .A2(new_n435), .B1(new_n454), .B2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(new_n447), .B1(new_n456), .B2(new_n410), .ZN(new_n457));
  INV_X1    g271(.A(new_n410), .ZN(new_n458));
  NAND3_X1  g272(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(new_n432), .B2(new_n434), .ZN(new_n460));
  AND3_X1   g274(.A1(new_n455), .A2(new_n199), .A3(new_n453), .ZN(new_n461));
  OAI211_X1 g275(.A(KEYINPUT83), .B(new_n458), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n442), .A2(new_n436), .A3(new_n410), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n457), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n464), .A2(new_n408), .A3(new_n221), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(KEYINPUT20), .ZN(new_n466));
  INV_X1    g280(.A(KEYINPUT20), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n464), .A2(new_n467), .A3(new_n408), .A4(new_n221), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n446), .B1(new_n466), .B2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT86), .ZN(new_n470));
  AOI21_X1  g284(.A(KEYINPUT13), .B1(new_n253), .B2(G128), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT85), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n204), .A2(G143), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n253), .A2(G128), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT13), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  AOI211_X1 g291(.A(KEYINPUT85), .B(KEYINPUT13), .C1(new_n253), .C2(G128), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n473), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n470), .B1(new_n479), .B2(new_n280), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n471), .B(new_n472), .ZN(new_n481));
  OAI211_X1 g295(.A(KEYINPUT86), .B(G134), .C1(new_n481), .C2(new_n477), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n475), .A2(new_n474), .A3(new_n483), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n483), .B1(new_n475), .B2(new_n474), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n280), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(G116), .B(G122), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(new_n239), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n480), .A2(new_n482), .A3(new_n486), .A4(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n349), .A2(G122), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n239), .B1(new_n490), .B2(KEYINPUT14), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT14), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n487), .A2(new_n492), .ZN(new_n493));
  AOI22_X1  g307(.A1(new_n491), .A2(new_n493), .B1(new_n239), .B2(new_n487), .ZN(new_n494));
  INV_X1    g308(.A(new_n486), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n484), .A2(new_n485), .A3(new_n280), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n494), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n188), .A2(new_n227), .A3(G953), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n489), .A2(new_n497), .A3(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n498), .B1(new_n489), .B2(new_n497), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n221), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT88), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n503), .A2(KEYINPUT15), .ZN(new_n506));
  OAI21_X1  g320(.A(G478), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n502), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n501), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(new_n499), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n511), .A2(new_n221), .A3(new_n507), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n469), .A2(new_n509), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n293), .A2(new_n295), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT66), .ZN(new_n515));
  XNOR2_X1  g329(.A(G134), .B(G137), .ZN(new_n516));
  OAI21_X1  g330(.A(new_n515), .B1(new_n516), .B2(new_n287), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n280), .A2(G137), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n282), .A2(G134), .ZN(new_n519));
  OAI211_X1 g333(.A(KEYINPUT66), .B(G131), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n288), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI22_X1  g336(.A1(new_n514), .A2(new_n522), .B1(new_n263), .B2(new_n310), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n367), .B1(new_n523), .B2(KEYINPUT70), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT70), .ZN(new_n525));
  AOI21_X1  g339(.A(new_n521), .B1(new_n293), .B2(new_n295), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n289), .A2(new_n262), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(KEYINPUT28), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT72), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n526), .A2(new_n527), .A3(new_n367), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n369), .B1(new_n356), .B2(new_n364), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n514), .A2(new_n522), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n263), .A2(new_n310), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT28), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(KEYINPUT72), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n531), .B1(new_n538), .B2(new_n529), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n417), .A2(G210), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(G101), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n541), .B(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n539), .A2(KEYINPUT29), .A3(new_n543), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n534), .A2(KEYINPUT30), .A3(new_n535), .ZN(new_n545));
  NAND4_X1  g359(.A1(new_n275), .A2(new_n517), .A3(new_n288), .A4(new_n520), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n546), .B1(new_n289), .B2(new_n262), .ZN(new_n547));
  XOR2_X1   g361(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n549), .A3(new_n367), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n523), .A2(new_n533), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n543), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT29), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT28), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n547), .A2(new_n367), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n557), .B1(new_n551), .B2(new_n558), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n529), .A2(new_n559), .A3(new_n553), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT71), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n534), .A2(KEYINPUT70), .A3(new_n535), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n562), .A2(new_n533), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n523), .A2(KEYINPUT70), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n557), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n551), .A2(new_n558), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(KEYINPUT28), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(new_n567), .A3(new_n543), .ZN(new_n568));
  AOI21_X1  g382(.A(KEYINPUT29), .B1(new_n552), .B2(new_n553), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT71), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n544), .A2(new_n561), .A3(new_n221), .A4(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(G472), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n550), .A2(new_n551), .A3(new_n543), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT31), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n550), .A2(KEYINPUT31), .A3(new_n551), .A4(new_n543), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n553), .B1(new_n529), .B2(new_n559), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(G472), .A2(G902), .ZN(new_n581));
  AOI21_X1  g395(.A(KEYINPUT32), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(KEYINPUT32), .ZN(new_n583));
  INV_X1    g397(.A(new_n581), .ZN(new_n584));
  AOI211_X1 g398(.A(new_n583), .B(new_n584), .C1(new_n578), .C2(new_n579), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n513), .B1(new_n573), .B2(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n334), .A2(new_n407), .A3(new_n587), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(new_n247), .Z(G3));
  INV_X1    g403(.A(KEYINPUT33), .ZN(new_n590));
  INV_X1    g404(.A(new_n498), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n591), .B2(KEYINPUT90), .ZN(new_n592));
  INV_X1    g406(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n511), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n510), .A2(new_n499), .A3(new_n592), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n594), .A2(G478), .A3(new_n221), .A4(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT91), .B(G478), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n502), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n601), .A2(new_n469), .ZN(new_n602));
  AND2_X1   g416(.A1(new_n407), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n578), .B2(new_n579), .ZN(new_n604));
  INV_X1    g418(.A(G472), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n565), .A2(new_n567), .ZN(new_n606));
  AOI22_X1  g420(.A1(new_n576), .A2(new_n577), .B1(new_n606), .B2(new_n553), .ZN(new_n607));
  OAI22_X1  g421(.A1(new_n604), .A2(new_n605), .B1(new_n607), .B2(new_n584), .ZN(new_n608));
  INV_X1    g422(.A(new_n608), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n603), .A2(new_n334), .A3(new_n609), .ZN(new_n610));
  XOR2_X1   g424(.A(KEYINPUT34), .B(G104), .Z(new_n611));
  XNOR2_X1  g425(.A(new_n610), .B(new_n611), .ZN(G6));
  NAND2_X1  g426(.A1(new_n321), .A2(new_n325), .ZN(new_n613));
  AND4_X1   g427(.A1(new_n327), .A2(new_n613), .A3(new_n236), .A4(new_n221), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n327), .B1(new_n326), .B2(new_n236), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n333), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(new_n235), .ZN(new_n617));
  NAND4_X1  g431(.A1(new_n616), .A2(new_n609), .A3(new_n189), .A4(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n405), .A2(new_n406), .ZN(new_n619));
  AOI221_X4 g433(.A(new_n446), .B1(new_n509), .B2(new_n512), .C1(new_n466), .C2(new_n468), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n619), .A2(new_n620), .A3(new_n345), .A4(new_n347), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT92), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n348), .B1(new_n405), .B2(new_n406), .ZN(new_n624));
  NAND4_X1  g438(.A1(new_n624), .A2(KEYINPUT92), .A3(new_n345), .A4(new_n620), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n618), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(KEYINPUT35), .B(G107), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G9));
  AOI21_X1  g442(.A(new_n190), .B1(new_n329), .B2(new_n333), .ZN(new_n629));
  XNOR2_X1  g443(.A(new_n213), .B(KEYINPUT93), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n219), .A2(KEYINPUT36), .ZN(new_n631));
  AND2_X1   g445(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n233), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n231), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT94), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n231), .A2(new_n634), .A3(KEYINPUT94), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n513), .A2(new_n608), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n629), .A2(new_n407), .A3(new_n639), .A4(new_n640), .ZN(new_n641));
  XOR2_X1   g455(.A(KEYINPUT95), .B(KEYINPUT96), .Z(new_n642));
  XNOR2_X1  g456(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g457(.A(KEYINPUT37), .B(G110), .Z(new_n644));
  XNOR2_X1  g458(.A(new_n643), .B(new_n644), .ZN(G12));
  NAND2_X1  g459(.A1(new_n629), .A2(new_n639), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n573), .A2(new_n586), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(new_n624), .ZN(new_n648));
  NOR2_X1   g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n509), .A2(new_n512), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n469), .A2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n341), .ZN(new_n652));
  INV_X1    g466(.A(G900), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n652), .B1(new_n653), .B2(new_n343), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(KEYINPUT97), .B1(new_n649), .B2(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT97), .ZN(new_n657));
  INV_X1    g471(.A(new_n655), .ZN(new_n658));
  NOR4_X1   g472(.A1(new_n646), .A2(new_n648), .A3(new_n657), .A4(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(new_n204), .ZN(G30));
  OAI21_X1  g475(.A(new_n553), .B1(new_n532), .B2(new_n536), .ZN(new_n662));
  INV_X1    g476(.A(KEYINPUT99), .ZN(new_n663));
  OAI21_X1  g477(.A(new_n574), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n662), .A2(new_n663), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n221), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n666), .A2(G472), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n586), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(KEYINPUT100), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n669), .A2(new_n635), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n654), .B(KEYINPUT39), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n629), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n348), .B1(new_n673), .B2(KEYINPUT40), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n469), .B1(new_n509), .B2(new_n512), .ZN(new_n676));
  XNOR2_X1  g490(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n619), .B(new_n677), .ZN(new_n678));
  OAI211_X1 g492(.A(new_n676), .B(new_n678), .C1(new_n673), .C2(KEYINPUT40), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n675), .A2(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n680), .B(G143), .ZN(G45));
  INV_X1    g495(.A(new_n654), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n649), .A2(new_n602), .A3(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT101), .B(G146), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G48));
  AND3_X1   g499(.A1(new_n568), .A2(new_n569), .A3(new_n570), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n570), .B1(new_n568), .B2(new_n569), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n565), .A2(KEYINPUT72), .A3(new_n537), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n555), .B1(new_n689), .B2(new_n531), .ZN(new_n690));
  AOI21_X1  g504(.A(G902), .B1(new_n690), .B2(new_n543), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n605), .B1(new_n688), .B2(new_n691), .ZN(new_n692));
  OAI21_X1  g506(.A(new_n583), .B1(new_n607), .B2(new_n584), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n580), .A2(KEYINPUT32), .A3(new_n581), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n617), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  OR2_X1    g510(.A1(new_n326), .A2(new_n236), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n329), .A2(new_n189), .A3(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n603), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND2_X1  g516(.A1(new_n623), .A2(new_n625), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(new_n699), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(G116), .ZN(G18));
  INV_X1    g519(.A(new_n698), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n706), .A2(new_n587), .A3(new_n407), .A4(new_n639), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G119), .ZN(G21));
  INV_X1    g522(.A(new_n624), .ZN(new_n709));
  NOR2_X1   g523(.A1(new_n698), .A2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n604), .A2(new_n605), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n689), .A2(new_n553), .A3(new_n531), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n584), .B1(new_n712), .B2(new_n578), .ZN(new_n713));
  NOR4_X1   g527(.A1(new_n711), .A2(new_n235), .A3(new_n346), .A4(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n710), .A2(new_n676), .A3(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G122), .ZN(G24));
  NOR2_X1   g530(.A1(new_n711), .A2(new_n713), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n635), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n602), .A2(new_n682), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(new_n710), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G125), .ZN(G27));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT102), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n616), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n329), .A2(KEYINPUT102), .A3(new_n333), .ZN(new_n726));
  AND3_X1   g540(.A1(new_n725), .A2(new_n189), .A3(new_n726), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n235), .B1(new_n573), .B2(new_n586), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n619), .A2(new_n348), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n729), .A2(new_n602), .A3(new_n682), .ZN(new_n730));
  INV_X1    g544(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT42), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n723), .B1(new_n732), .B2(new_n733), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n728), .A2(new_n725), .A3(new_n189), .A4(new_n726), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n723), .B(new_n733), .C1(new_n735), .C2(new_n730), .ZN(new_n736));
  INV_X1    g550(.A(new_n736), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT104), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n725), .A2(new_n189), .A3(new_n726), .ZN(new_n739));
  NOR3_X1   g553(.A1(new_n739), .A2(new_n696), .A3(new_n730), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n738), .B1(new_n740), .B2(KEYINPUT42), .ZN(new_n741));
  NOR4_X1   g555(.A1(new_n735), .A2(KEYINPUT104), .A3(new_n733), .A4(new_n730), .ZN(new_n742));
  OAI22_X1  g556(.A1(new_n734), .A2(new_n737), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  INV_X1    g558(.A(new_n729), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n735), .A2(new_n658), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(new_n280), .ZN(G36));
  OR2_X1    g561(.A1(new_n332), .A2(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n332), .A2(KEYINPUT45), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n748), .A2(G469), .A3(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(G469), .A2(G902), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(KEYINPUT46), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n329), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT46), .B1(new_n750), .B2(new_n751), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n189), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  OR2_X1    g569(.A1(new_n755), .A2(new_n671), .ZN(new_n756));
  XOR2_X1   g570(.A(new_n756), .B(KEYINPUT105), .Z(new_n757));
  INV_X1    g571(.A(new_n469), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n601), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(KEYINPUT43), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n760), .A2(new_n608), .A3(new_n635), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR3_X1   g578(.A1(new_n763), .A2(new_n764), .A3(new_n745), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G137), .ZN(G39));
  INV_X1    g581(.A(KEYINPUT106), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT47), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n755), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n768), .A2(new_n769), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n770), .B1(new_n755), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n647), .A2(new_n617), .ZN(new_n774));
  INV_X1    g588(.A(new_n774), .ZN(new_n775));
  NOR4_X1   g589(.A1(new_n771), .A2(new_n773), .A3(new_n730), .A4(new_n775), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(new_n193), .ZN(G42));
  NAND2_X1  g591(.A1(new_n329), .A2(new_n697), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT107), .Z(new_n779));
  INV_X1    g593(.A(KEYINPUT49), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n779), .A2(new_n780), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n781), .A2(new_n782), .A3(new_n759), .ZN(new_n783));
  INV_X1    g597(.A(new_n669), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n784), .A2(new_n190), .A3(new_n678), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n783), .A2(new_n617), .A3(new_n347), .A4(new_n785), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT54), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n624), .A2(new_n676), .ZN(new_n788));
  INV_X1    g602(.A(new_n788), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n670), .A2(new_n682), .A3(new_n727), .A4(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n683), .B(new_n721), .C1(new_n656), .C2(new_n659), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT52), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n646), .A2(new_n648), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n794), .A2(new_n719), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n657), .B1(new_n794), .B2(new_n658), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n649), .A2(KEYINPUT97), .A3(new_n655), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n795), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n798), .A2(new_n799), .A3(new_n721), .A4(new_n790), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n793), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n725), .A2(new_n189), .A3(new_n726), .A4(new_n602), .ZN(new_n802));
  INV_X1    g616(.A(new_n587), .ZN(new_n803));
  OAI22_X1  g617(.A1(new_n802), .A2(new_n718), .B1(new_n803), .B2(new_n646), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n682), .A3(new_n729), .ZN(new_n805));
  INV_X1    g619(.A(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n727), .A2(KEYINPUT42), .A3(new_n728), .A4(new_n731), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(KEYINPUT104), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n740), .A2(new_n738), .A3(KEYINPUT42), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g624(.A(new_n733), .B1(new_n735), .B2(new_n730), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT103), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n736), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n806), .B1(new_n810), .B2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n513), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n647), .A2(new_n407), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n629), .A2(new_n617), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n641), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n651), .A2(KEYINPUT108), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n758), .A2(new_n600), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT108), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n469), .A2(new_n821), .A3(new_n650), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n819), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n823), .A2(new_n407), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n618), .ZN(new_n825));
  OAI21_X1  g639(.A(KEYINPUT109), .B1(new_n818), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n334), .A2(new_n407), .A3(new_n609), .A4(new_n823), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n827), .A2(new_n588), .A3(new_n828), .A4(new_n641), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(new_n746), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n704), .A2(new_n700), .A3(new_n707), .A4(new_n715), .ZN(new_n832));
  INV_X1    g646(.A(new_n832), .ZN(new_n833));
  AND3_X1   g647(.A1(new_n830), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n801), .A2(KEYINPUT53), .A3(new_n814), .A4(new_n834), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n793), .A2(new_n800), .ZN(new_n836));
  AOI21_X1  g650(.A(new_n832), .B1(new_n829), .B2(new_n826), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n743), .A2(new_n831), .A3(new_n805), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT110), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT110), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n834), .A2(new_n814), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n836), .B1(new_n839), .B2(new_n841), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT111), .B(KEYINPUT53), .ZN(new_n843));
  OAI211_X1 g657(.A(new_n787), .B(new_n835), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  AND3_X1   g660(.A1(new_n834), .A2(new_n814), .A3(new_n840), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n840), .B1(new_n834), .B2(new_n814), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n801), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  INV_X1    g663(.A(new_n843), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n851), .A2(KEYINPUT112), .A3(new_n787), .A4(new_n835), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n849), .A2(KEYINPUT53), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n842), .A2(new_n850), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n853), .A2(new_n854), .A3(KEYINPUT54), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n846), .A2(new_n852), .A3(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n706), .A2(new_n729), .ZN(new_n857));
  INV_X1    g671(.A(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n669), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n617), .A2(new_n652), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n859), .A2(new_n820), .A3(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n859), .A2(new_n758), .A3(new_n600), .A4(new_n860), .ZN(new_n862));
  AND4_X1   g676(.A1(new_n617), .A2(new_n760), .A3(new_n652), .A4(new_n717), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n863), .A2(new_n706), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n678), .A2(new_n347), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT113), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n866), .A2(KEYINPUT50), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(KEYINPUT50), .ZN(new_n868));
  AOI21_X1  g682(.A(new_n862), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n779), .A2(new_n190), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n870), .B1(new_n771), .B2(new_n773), .ZN(new_n871));
  AND2_X1   g685(.A1(new_n863), .A2(new_n729), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n858), .A2(new_n652), .A3(new_n760), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n874), .A2(new_n718), .ZN(new_n875));
  INV_X1    g689(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n869), .A2(new_n873), .A3(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT51), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n874), .A2(new_n696), .ZN(new_n880));
  XOR2_X1   g694(.A(new_n880), .B(KEYINPUT48), .Z(new_n881));
  INV_X1    g695(.A(KEYINPUT114), .ZN(new_n882));
  OR2_X1    g696(.A1(new_n871), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n871), .A2(new_n882), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n872), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n869), .A2(KEYINPUT51), .A3(new_n876), .A4(new_n885), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n879), .A2(new_n338), .A3(new_n881), .A4(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n864), .A2(new_n709), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n888), .B(KEYINPUT115), .ZN(new_n889));
  NOR4_X1   g703(.A1(new_n856), .A2(new_n861), .A3(new_n887), .A4(new_n889), .ZN(new_n890));
  NOR2_X1   g704(.A1(G952), .A2(G953), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT116), .Z(new_n892));
  OAI21_X1  g706(.A(new_n786), .B1(new_n890), .B2(new_n892), .ZN(G75));
  INV_X1    g707(.A(KEYINPUT53), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n836), .A2(new_n838), .A3(new_n894), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n849), .B2(new_n850), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n896), .A2(new_n221), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(G210), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT56), .ZN(new_n899));
  AND2_X1   g713(.A1(new_n381), .A2(new_n389), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n900), .B(new_n387), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n901), .B(KEYINPUT55), .Z(new_n902));
  AND3_X1   g716(.A1(new_n898), .A2(new_n899), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n898), .B2(new_n899), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n214), .A2(G952), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(G51));
  XOR2_X1   g720(.A(new_n751), .B(KEYINPUT57), .Z(new_n907));
  NOR2_X1   g721(.A1(new_n896), .A2(new_n787), .ZN(new_n908));
  INV_X1    g722(.A(new_n844), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(KEYINPUT117), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT117), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n912), .B(new_n907), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n911), .A2(new_n613), .A3(new_n913), .ZN(new_n914));
  OR3_X1    g728(.A1(new_n896), .A2(new_n221), .A3(new_n750), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n905), .B1(new_n914), .B2(new_n915), .ZN(G54));
  NAND3_X1  g730(.A1(new_n897), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  INV_X1    g731(.A(new_n464), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n917), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n905), .ZN(G60));
  XNOR2_X1  g735(.A(KEYINPUT118), .B(KEYINPUT59), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n922), .B(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n856), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n594), .A2(new_n595), .ZN(new_n926));
  AOI21_X1  g740(.A(KEYINPUT119), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  INV_X1    g741(.A(KEYINPUT119), .ZN(new_n928));
  INV_X1    g742(.A(new_n926), .ZN(new_n929));
  AOI211_X1 g743(.A(new_n928), .B(new_n929), .C1(new_n856), .C2(new_n924), .ZN(new_n930));
  INV_X1    g744(.A(new_n905), .ZN(new_n931));
  OAI21_X1  g745(.A(new_n924), .B1(new_n908), .B2(new_n909), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n926), .ZN(new_n933));
  NOR3_X1   g747(.A1(new_n927), .A2(new_n930), .A3(new_n933), .ZN(G63));
  NAND2_X1  g748(.A1(new_n851), .A2(new_n835), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n632), .A2(new_n633), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(KEYINPUT120), .B(KEYINPUT60), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n227), .A2(new_n221), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n938), .B(new_n939), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n935), .A2(new_n937), .A3(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n232), .ZN(new_n942));
  INV_X1    g756(.A(new_n940), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n896), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n941), .A2(new_n944), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT122), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n945), .A2(new_n946), .ZN(new_n948));
  OAI211_X1 g762(.A(new_n931), .B(new_n944), .C1(new_n941), .C2(KEYINPUT121), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n941), .A2(KEYINPUT121), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI22_X1  g765(.A1(new_n947), .A2(new_n948), .B1(new_n951), .B2(KEYINPUT61), .ZN(G66));
  AOI21_X1  g766(.A(new_n214), .B1(new_n342), .B2(G224), .ZN(new_n953));
  INV_X1    g767(.A(new_n837), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n953), .B1(new_n954), .B2(new_n214), .ZN(new_n955));
  INV_X1    g769(.A(G898), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n900), .B1(new_n956), .B2(G953), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n955), .B(new_n957), .ZN(G69));
  NAND2_X1  g772(.A1(new_n545), .A2(new_n549), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n450), .A2(new_n452), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n959), .B(new_n960), .Z(new_n961));
  INV_X1    g775(.A(new_n823), .ZN(new_n962));
  NOR4_X1   g776(.A1(new_n673), .A2(new_n962), .A3(new_n696), .A4(new_n745), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n757), .B2(new_n765), .ZN(new_n964));
  INV_X1    g778(.A(new_n792), .ZN(new_n965));
  NAND2_X1  g779(.A1(KEYINPUT123), .A2(KEYINPUT62), .ZN(new_n966));
  NAND3_X1  g780(.A1(new_n965), .A2(new_n680), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n965), .A2(new_n680), .ZN(new_n968));
  XNOR2_X1  g782(.A(KEYINPUT123), .B(KEYINPUT62), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n776), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g784(.A1(new_n964), .A2(new_n967), .A3(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(KEYINPUT124), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND4_X1  g787(.A1(new_n964), .A2(new_n970), .A3(KEYINPUT124), .A4(new_n967), .ZN(new_n974));
  AND2_X1   g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n961), .B1(new_n975), .B2(G953), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n653), .A2(new_n214), .ZN(new_n977));
  INV_X1    g791(.A(new_n961), .ZN(new_n978));
  NOR2_X1   g792(.A1(new_n696), .A2(new_n788), .ZN(new_n979));
  OR2_X1    g793(.A1(new_n765), .A2(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n746), .B1(new_n980), .B2(new_n757), .ZN(new_n981));
  INV_X1    g795(.A(new_n776), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n981), .A2(new_n743), .A3(new_n982), .A4(new_n965), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n978), .B1(new_n983), .B2(G953), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n976), .B1(new_n977), .B2(new_n984), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n214), .B1(G227), .B2(G900), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n985), .B(new_n986), .ZN(G72));
  XNOR2_X1  g801(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n605), .A2(new_n221), .ZN(new_n989));
  XOR2_X1   g803(.A(new_n988), .B(new_n989), .Z(new_n990));
  NAND2_X1  g804(.A1(new_n554), .A2(new_n574), .ZN(new_n991));
  AND4_X1   g805(.A1(new_n853), .A2(new_n854), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  XOR2_X1   g806(.A(new_n552), .B(KEYINPUT126), .Z(new_n993));
  NAND3_X1  g807(.A1(new_n973), .A2(new_n837), .A3(new_n974), .ZN(new_n994));
  AOI211_X1 g808(.A(new_n553), .B(new_n993), .C1(new_n994), .C2(new_n990), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n990), .B1(new_n983), .B2(new_n954), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n996), .A2(new_n553), .A3(new_n993), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n997), .A2(new_n931), .ZN(new_n998));
  OR2_X1    g812(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n998), .A2(KEYINPUT127), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n992), .B(new_n995), .C1(new_n999), .C2(new_n1000), .ZN(G57));
endmodule


