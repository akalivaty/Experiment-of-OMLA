//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:27 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n446, new_n450, new_n451, new_n453,
    new_n456, new_n457, new_n458, new_n459, new_n460, new_n461, new_n464,
    new_n465, new_n466, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n552, new_n554, new_n555, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n608, new_n611,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1172;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT64), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n446));
  XNOR2_X1  g021(.A(new_n446), .B(KEYINPUT65), .ZN(G259));
  BUF_X1    g022(.A(G452), .Z(G391));
  AND2_X1   g023(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g024(.A(KEYINPUT66), .B(KEYINPUT1), .ZN(new_n450));
  NAND2_X1  g025(.A1(G7), .A2(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(G223));
  INV_X1    g027(.A(new_n451), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n453), .A2(G567), .ZN(G234));
  NAND2_X1  g029(.A1(new_n453), .A2(G2106), .ZN(G217));
  NOR4_X1   g030(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT2), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR4_X1   g033(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n459));
  XNOR2_X1  g034(.A(new_n459), .B(KEYINPUT67), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(new_n461));
  NOR2_X1   g036(.A1(new_n458), .A2(new_n461), .ZN(G325));
  INV_X1    g037(.A(G325), .ZN(G261));
  NAND2_X1  g038(.A1(new_n458), .A2(G2106), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n461), .A2(G567), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(new_n466), .ZN(G319));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .A3(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .ZN(new_n471));
  AND2_X1   g046(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g047(.A(G2105), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT68), .ZN(new_n474));
  OAI21_X1  g049(.A(new_n474), .B1(new_n470), .B2(KEYINPUT3), .ZN(new_n475));
  AND3_X1   g050(.A1(new_n472), .A2(new_n473), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G137), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n468), .A2(G2104), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(new_n471), .ZN(new_n480));
  INV_X1    g055(.A(G125), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n482), .A2(G2105), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n473), .A2(G101), .A3(G2104), .ZN(new_n484));
  AND3_X1   g059(.A1(new_n477), .A2(new_n483), .A3(new_n484), .ZN(G160));
  NAND4_X1  g060(.A1(new_n475), .A2(new_n469), .A3(G2105), .A4(new_n471), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AND2_X1   g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(new_n490), .B1(G112), .B2(new_n473), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT69), .ZN(new_n492));
  AOI211_X1 g067(.A(new_n488), .B(new_n492), .C1(G136), .C2(new_n476), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT70), .ZN(G162));
  INV_X1    g069(.A(G126), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n473), .A2(G114), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  OAI22_X1  g072(.A1(new_n486), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n499), .A2(G2105), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n502), .A2(new_n480), .ZN(new_n503));
  NAND4_X1  g078(.A1(new_n475), .A2(new_n469), .A3(new_n500), .A4(new_n471), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT4), .ZN(new_n505));
  AOI21_X1  g080(.A(new_n503), .B1(new_n505), .B2(KEYINPUT71), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT71), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT4), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n498), .B1(new_n506), .B2(new_n508), .ZN(G164));
  XNOR2_X1  g084(.A(KEYINPUT72), .B(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT6), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT6), .A2(G651), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  XNOR2_X1  g089(.A(KEYINPUT5), .B(G543), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n515), .A2(G88), .B1(G50), .B2(G543), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n515), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(new_n510), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  INV_X1    g096(.A(new_n515), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G89), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n525), .A2(KEYINPUT7), .ZN(new_n527));
  AND2_X1   g102(.A1(G63), .A2(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n526), .A2(new_n527), .B1(new_n515), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n512), .A2(new_n513), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT73), .ZN(new_n531));
  OR3_X1    g106(.A1(new_n512), .A2(KEYINPUT73), .A3(new_n513), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n531), .A2(G543), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(G51), .ZN(new_n534));
  OAI211_X1 g109(.A(new_n524), .B(new_n529), .C1(new_n533), .C2(new_n534), .ZN(new_n535));
  XNOR2_X1  g110(.A(new_n535), .B(KEYINPUT74), .ZN(G168));
  INV_X1    g111(.A(new_n533), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n537), .A2(G52), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n539));
  OR2_X1    g114(.A1(new_n539), .A2(new_n510), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n523), .A2(G90), .ZN(new_n541));
  NAND3_X1  g116(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(G301));
  INV_X1    g117(.A(G301), .ZN(G171));
  NAND2_X1  g118(.A1(new_n537), .A2(G43), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n523), .A2(G81), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n515), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n546));
  AOI21_X1  g121(.A(new_n510), .B1(new_n546), .B2(KEYINPUT75), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n547), .B1(KEYINPUT75), .B2(new_n546), .ZN(new_n548));
  AND3_X1   g123(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n549), .A2(G860), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT76), .ZN(G153));
  NAND4_X1  g126(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n552));
  XOR2_X1   g127(.A(new_n552), .B(KEYINPUT77), .Z(G176));
  NAND2_X1  g128(.A1(G1), .A2(G3), .ZN(new_n554));
  XNOR2_X1  g129(.A(new_n554), .B(KEYINPUT8), .ZN(new_n555));
  NAND4_X1  g130(.A1(G319), .A2(G483), .A3(G661), .A4(new_n555), .ZN(G188));
  INV_X1    g131(.A(G53), .ZN(new_n557));
  OAI21_X1  g132(.A(KEYINPUT9), .B1(new_n533), .B2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n559), .B1(new_n530), .B2(KEYINPUT73), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n560), .A2(new_n561), .A3(G53), .A4(new_n532), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n558), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT78), .ZN(new_n564));
  OR2_X1    g139(.A1(new_n564), .A2(G65), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(G65), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n515), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(G78), .ZN(new_n568));
  OAI21_X1  g143(.A(new_n567), .B1(new_n568), .B2(new_n559), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n523), .A2(G91), .B1(G651), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(KEYINPUT79), .ZN(new_n572));
  XNOR2_X1  g147(.A(new_n571), .B(new_n572), .ZN(G299));
  INV_X1    g148(.A(G168), .ZN(G286));
  NAND2_X1  g149(.A1(new_n537), .A2(G49), .ZN(new_n575));
  OAI21_X1  g150(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n523), .A2(G87), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(G288));
  AOI22_X1  g153(.A1(new_n515), .A2(G86), .B1(G48), .B2(G543), .ZN(new_n579));
  NOR2_X1   g154(.A1(new_n514), .A2(new_n579), .ZN(new_n580));
  AOI22_X1  g155(.A1(new_n515), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n581));
  NOR2_X1   g156(.A1(new_n581), .A2(new_n510), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n580), .A2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(G305));
  XNOR2_X1  g159(.A(KEYINPUT81), .B(G85), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n523), .A2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G47), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n586), .B1(new_n533), .B2(new_n587), .ZN(new_n588));
  AND2_X1   g163(.A1(new_n588), .A2(KEYINPUT82), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n510), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT80), .ZN(new_n592));
  OAI21_X1  g167(.A(new_n592), .B1(new_n588), .B2(KEYINPUT82), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n589), .A2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n523), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT10), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n537), .A2(G54), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  XOR2_X1   g174(.A(KEYINPUT83), .B(G66), .Z(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n522), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n601), .A2(G651), .ZN(new_n602));
  AND3_X1   g177(.A1(new_n597), .A2(new_n598), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n595), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n595), .B1(new_n603), .B2(G868), .ZN(G321));
  INV_X1    g180(.A(G868), .ZN(new_n606));
  NOR2_X1   g181(.A1(G286), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n571), .B(KEYINPUT79), .ZN(new_n608));
  AOI21_X1  g183(.A(new_n607), .B1(new_n606), .B2(new_n608), .ZN(G297));
  XNOR2_X1  g184(.A(G297), .B(KEYINPUT84), .ZN(G280));
  INV_X1    g185(.A(G559), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n603), .B1(new_n611), .B2(G860), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT85), .ZN(G148));
  NAND2_X1  g188(.A1(new_n603), .A2(new_n611), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G868), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n549), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g192(.A(G123), .ZN(new_n618));
  OAI21_X1  g193(.A(KEYINPUT88), .B1(new_n473), .B2(G111), .ZN(new_n619));
  OR2_X1    g194(.A1(G99), .A2(G2105), .ZN(new_n620));
  NAND3_X1  g195(.A1(new_n619), .A2(G2104), .A3(new_n620), .ZN(new_n621));
  NOR3_X1   g196(.A1(new_n473), .A2(KEYINPUT88), .A3(G111), .ZN(new_n622));
  OAI22_X1  g197(.A1(new_n486), .A2(new_n618), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  AOI21_X1  g198(.A(KEYINPUT87), .B1(new_n476), .B2(G135), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n476), .A2(KEYINPUT87), .A3(G135), .ZN(new_n626));
  AOI21_X1  g201(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g202(.A(new_n627), .ZN(new_n628));
  OR2_X1    g203(.A1(new_n628), .A2(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(G2096), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n473), .A2(G2104), .ZN(new_n631));
  NOR2_X1   g206(.A1(new_n480), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XOR2_X1   g208(.A(KEYINPUT86), .B(G2100), .Z(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(KEYINPUT13), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n633), .B(new_n635), .ZN(new_n636));
  NAND3_X1  g211(.A1(new_n629), .A2(new_n630), .A3(new_n636), .ZN(G156));
  INV_X1    g212(.A(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2438), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G2430), .ZN(new_n640));
  XNOR2_X1  g215(.A(KEYINPUT15), .B(G2435), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n638), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  OAI21_X1  g217(.A(new_n642), .B1(new_n641), .B2(new_n640), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(G1341), .B(G1348), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n645), .B(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(new_n643), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  OR2_X1    g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n649), .ZN(new_n651));
  AND3_X1   g226(.A1(new_n650), .A2(G14), .A3(new_n651), .ZN(G401));
  XNOR2_X1  g227(.A(G2067), .B(G2678), .ZN(new_n653));
  NOR2_X1   g228(.A1(G2072), .A2(G2078), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n444), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g231(.A(new_n653), .B1(new_n656), .B2(KEYINPUT89), .ZN(new_n657));
  OAI21_X1  g232(.A(new_n657), .B1(KEYINPUT89), .B2(new_n656), .ZN(new_n658));
  XOR2_X1   g233(.A(G2084), .B(G2090), .Z(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n655), .B(KEYINPUT17), .ZN(new_n661));
  INV_X1    g236(.A(new_n653), .ZN(new_n662));
  OAI211_X1 g237(.A(new_n658), .B(new_n660), .C1(new_n661), .C2(new_n662), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n660), .A2(new_n655), .A3(new_n662), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT18), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n661), .A2(new_n662), .A3(new_n659), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g242(.A(G2096), .B(G2100), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(G227));
  XOR2_X1   g244(.A(G1971), .B(G1976), .Z(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT19), .ZN(new_n671));
  XNOR2_X1  g246(.A(G1956), .B(G2474), .ZN(new_n672));
  XNOR2_X1  g247(.A(G1961), .B(G1966), .ZN(new_n673));
  NOR2_X1   g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  AND2_X1   g249(.A1(new_n672), .A2(new_n673), .ZN(new_n675));
  NOR3_X1   g250(.A1(new_n671), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n671), .A2(new_n674), .ZN(new_n677));
  XOR2_X1   g252(.A(new_n677), .B(KEYINPUT20), .Z(new_n678));
  AOI211_X1 g253(.A(new_n676), .B(new_n678), .C1(new_n671), .C2(new_n675), .ZN(new_n679));
  XNOR2_X1  g254(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n680));
  XOR2_X1   g255(.A(new_n679), .B(new_n680), .Z(new_n681));
  XNOR2_X1  g256(.A(G1991), .B(G1996), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(KEYINPUT90), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n681), .B(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(G1981), .B(G1986), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(G229));
  INV_X1    g261(.A(G288), .ZN(new_n687));
  INV_X1    g262(.A(G16), .ZN(new_n688));
  NOR2_X1   g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n688), .B2(G23), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g266(.A(KEYINPUT33), .B(G1976), .Z(new_n692));
  OR2_X1    g267(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n691), .A2(new_n692), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n688), .A2(G22), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G166), .B2(new_n688), .ZN(new_n696));
  INV_X1    g271(.A(G1971), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g273(.A1(G6), .A2(G16), .ZN(new_n699));
  AOI21_X1  g274(.A(new_n699), .B1(new_n583), .B2(G16), .ZN(new_n700));
  XOR2_X1   g275(.A(KEYINPUT32), .B(G1981), .Z(new_n701));
  XNOR2_X1  g276(.A(new_n700), .B(new_n701), .ZN(new_n702));
  NAND4_X1  g277(.A1(new_n693), .A2(new_n694), .A3(new_n698), .A4(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT34), .Z(new_n704));
  NAND2_X1  g279(.A1(new_n688), .A2(G24), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n589), .A2(new_n593), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n706), .B2(new_n688), .ZN(new_n707));
  INV_X1    g282(.A(G1986), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n711));
  OR2_X1    g286(.A1(new_n710), .A2(KEYINPUT95), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT91), .B(G29), .Z(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G25), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT92), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n487), .A2(G119), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n473), .A2(G107), .ZN(new_n717));
  OAI21_X1  g292(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G131), .B2(new_n476), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT93), .ZN(new_n721));
  INV_X1    g296(.A(new_n713), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n715), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n723), .B(KEYINPUT94), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT35), .B(G1991), .Z(new_n725));
  INV_X1    g300(.A(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n724), .B(new_n726), .ZN(new_n727));
  NAND4_X1  g302(.A1(new_n704), .A2(new_n711), .A3(new_n712), .A4(new_n727), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT36), .ZN(new_n729));
  OR3_X1    g304(.A1(new_n728), .A2(KEYINPUT96), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(KEYINPUT96), .B(KEYINPUT36), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n713), .A2(G26), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  OR2_X1    g309(.A1(G104), .A2(G2105), .ZN(new_n735));
  OAI211_X1 g310(.A(new_n735), .B(G2104), .C1(G116), .C2(new_n473), .ZN(new_n736));
  INV_X1    g311(.A(G128), .ZN(new_n737));
  INV_X1    g312(.A(new_n476), .ZN(new_n738));
  INV_X1    g313(.A(G140), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n736), .B1(new_n737), .B2(new_n486), .C1(new_n738), .C2(new_n739), .ZN(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n734), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G2067), .ZN(new_n744));
  NOR2_X1   g319(.A1(G5), .A2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT99), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G301), .B2(new_n688), .ZN(new_n747));
  INV_X1    g322(.A(G1961), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  NOR2_X1   g324(.A1(G16), .A2(G19), .ZN(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n549), .B2(G16), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n744), .B(new_n749), .C1(G1341), .C2(new_n751), .ZN(new_n752));
  NOR2_X1   g327(.A1(G168), .A2(new_n688), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n753), .B1(new_n688), .B2(G21), .ZN(new_n754));
  XNOR2_X1  g329(.A(KEYINPUT98), .B(G1966), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n754), .A2(new_n755), .ZN(new_n757));
  NOR2_X1   g332(.A1(new_n722), .A2(G27), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(G164), .B2(new_n722), .ZN(new_n759));
  XNOR2_X1  g334(.A(new_n759), .B(new_n443), .ZN(new_n760));
  NAND4_X1  g335(.A1(new_n752), .A2(new_n756), .A3(new_n757), .A4(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n722), .A2(G35), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n722), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  OR2_X1    g339(.A1(new_n764), .A2(G2090), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(G2090), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n751), .A2(G1341), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n476), .A2(G139), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n473), .A2(G103), .A3(G2104), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT25), .ZN(new_n770));
  NAND2_X1  g345(.A1(G115), .A2(G2104), .ZN(new_n771));
  INV_X1    g346(.A(G127), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n771), .B1(new_n480), .B2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n770), .B1(G2105), .B2(new_n773), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n775), .A2(new_n742), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(new_n742), .B2(G33), .ZN(new_n777));
  OR2_X1    g352(.A1(new_n777), .A2(new_n442), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT24), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n779), .A2(G34), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n779), .A2(G34), .ZN(new_n781));
  NAND3_X1  g356(.A1(new_n713), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G160), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n782), .B1(new_n783), .B2(new_n742), .ZN(new_n784));
  INV_X1    g359(.A(G2084), .ZN(new_n785));
  NAND2_X1  g360(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n777), .A2(new_n442), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n784), .A2(new_n785), .ZN(new_n788));
  NAND4_X1  g363(.A1(new_n778), .A2(new_n786), .A3(new_n787), .A4(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n742), .A2(G32), .ZN(new_n790));
  NAND3_X1  g365(.A1(new_n473), .A2(G105), .A3(G2104), .ZN(new_n791));
  NAND3_X1  g366(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT97), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(KEYINPUT26), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n476), .A2(G141), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n487), .A2(G129), .ZN(new_n796));
  AND4_X1   g371(.A1(new_n791), .A2(new_n794), .A3(new_n795), .A4(new_n796), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n790), .B1(new_n797), .B2(new_n742), .ZN(new_n798));
  XOR2_X1   g373(.A(KEYINPUT27), .B(G1996), .Z(new_n799));
  NOR2_X1   g374(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n798), .A2(new_n799), .ZN(new_n801));
  INV_X1    g376(.A(KEYINPUT30), .ZN(new_n802));
  AND2_X1   g377(.A1(new_n802), .A2(G28), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n742), .B1(new_n802), .B2(G28), .ZN(new_n804));
  AND2_X1   g379(.A1(KEYINPUT31), .A2(G11), .ZN(new_n805));
  NOR2_X1   g380(.A1(KEYINPUT31), .A2(G11), .ZN(new_n806));
  OAI22_X1  g381(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n627), .B2(new_n722), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n801), .A2(new_n808), .ZN(new_n809));
  NOR4_X1   g384(.A1(new_n767), .A2(new_n789), .A3(new_n800), .A4(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n688), .A2(G4), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n603), .B2(new_n688), .ZN(new_n812));
  INV_X1    g387(.A(G1348), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND4_X1  g389(.A1(new_n765), .A2(new_n766), .A3(new_n810), .A4(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n688), .A2(G20), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT23), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n608), .B2(new_n688), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(G1956), .ZN(new_n819));
  NOR3_X1   g394(.A1(new_n761), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n730), .A2(new_n732), .A3(new_n820), .ZN(G150));
  INV_X1    g396(.A(G150), .ZN(G311));
  INV_X1    g397(.A(KEYINPUT100), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n523), .A2(G93), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n510), .B2(new_n825), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n826), .B1(new_n537), .B2(G55), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n549), .A2(new_n823), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n823), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n544), .A2(new_n545), .A3(new_n548), .ZN(new_n830));
  INV_X1    g405(.A(G55), .ZN(new_n831));
  OAI221_X1 g406(.A(new_n824), .B1(new_n510), .B2(new_n825), .C1(new_n533), .C2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(KEYINPUT100), .ZN(new_n833));
  NAND3_X1  g408(.A1(new_n829), .A2(new_n830), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n835), .B(KEYINPUT38), .Z(new_n836));
  NAND2_X1  g411(.A1(new_n603), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n836), .B(new_n837), .ZN(new_n838));
  OR2_X1    g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  INV_X1    g414(.A(G860), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n841));
  NAND3_X1  g416(.A1(new_n839), .A2(new_n840), .A3(new_n841), .ZN(new_n842));
  NOR2_X1   g417(.A1(new_n827), .A2(new_n840), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n843), .B(KEYINPUT37), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(G145));
  XNOR2_X1  g420(.A(new_n797), .B(new_n740), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n847));
  INV_X1    g422(.A(new_n503), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n847), .A2(new_n508), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n498), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n851), .A2(KEYINPUT101), .ZN(new_n852));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n853));
  NAND2_X1  g428(.A1(G164), .A2(new_n853), .ZN(new_n854));
  AND2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  XOR2_X1   g430(.A(new_n846), .B(new_n855), .Z(new_n856));
  AOI21_X1  g431(.A(new_n775), .B1(new_n856), .B2(KEYINPUT104), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(KEYINPUT104), .B2(new_n856), .ZN(new_n858));
  INV_X1    g433(.A(new_n775), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(KEYINPUT102), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n846), .B(new_n855), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n859), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g439(.A(new_n858), .B1(new_n864), .B2(KEYINPUT103), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n865), .B1(KEYINPUT103), .B2(new_n864), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n476), .A2(G142), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n487), .A2(G130), .ZN(new_n868));
  NOR3_X1   g443(.A1(new_n473), .A2(KEYINPUT105), .A3(G118), .ZN(new_n869));
  OAI21_X1  g444(.A(KEYINPUT105), .B1(new_n473), .B2(G118), .ZN(new_n870));
  OR2_X1    g445(.A1(G106), .A2(G2105), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n870), .A2(G2104), .A3(new_n871), .ZN(new_n872));
  OAI211_X1 g447(.A(new_n867), .B(new_n868), .C1(new_n869), .C2(new_n872), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n633), .Z(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(new_n721), .Z(new_n875));
  XOR2_X1   g450(.A(new_n875), .B(KEYINPUT106), .Z(new_n876));
  NAND2_X1  g451(.A1(new_n866), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G162), .B(new_n783), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n878), .B(new_n628), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  OAI211_X1 g455(.A(new_n877), .B(new_n879), .C1(new_n866), .C2(new_n880), .ZN(new_n881));
  INV_X1    g456(.A(G37), .ZN(new_n882));
  XOR2_X1   g457(.A(new_n866), .B(new_n876), .Z(new_n883));
  OAI211_X1 g458(.A(new_n881), .B(new_n882), .C1(new_n883), .C2(new_n879), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g460(.A1(new_n832), .A2(new_n606), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n706), .B(G288), .ZN(new_n887));
  XNOR2_X1  g462(.A(G303), .B(new_n583), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(KEYINPUT109), .ZN(new_n890));
  OR2_X1    g465(.A1(new_n887), .A2(new_n888), .ZN(new_n891));
  AND2_X1   g466(.A1(new_n891), .A2(KEYINPUT108), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n891), .A2(KEYINPUT108), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n890), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT42), .ZN(new_n895));
  NAND2_X1  g470(.A1(G299), .A2(KEYINPUT107), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT107), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n608), .A2(new_n897), .ZN(new_n898));
  INV_X1    g473(.A(new_n603), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n896), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n608), .A2(new_n897), .A3(new_n603), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  XNOR2_X1  g477(.A(new_n902), .B(KEYINPUT41), .ZN(new_n903));
  INV_X1    g478(.A(new_n902), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n835), .B(new_n614), .ZN(new_n905));
  MUX2_X1   g480(.A(new_n903), .B(new_n904), .S(new_n905), .Z(new_n906));
  XNOR2_X1  g481(.A(new_n895), .B(new_n906), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n886), .B1(new_n907), .B2(new_n606), .ZN(G295));
  OAI21_X1  g483(.A(new_n886), .B1(new_n907), .B2(new_n606), .ZN(G331));
  INV_X1    g484(.A(KEYINPUT43), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n835), .A2(G286), .ZN(new_n911));
  AOI21_X1  g486(.A(G168), .B1(new_n828), .B2(new_n834), .ZN(new_n912));
  OR3_X1    g487(.A1(new_n911), .A2(G301), .A3(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(G301), .B1(new_n911), .B2(new_n912), .ZN(new_n914));
  NAND2_X1  g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n903), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n904), .A2(new_n913), .A3(new_n914), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n916), .A2(new_n894), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(new_n882), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n894), .B1(new_n916), .B2(new_n917), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n910), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n917), .A2(KEYINPUT110), .ZN(new_n922));
  OR3_X1    g497(.A1(new_n915), .A2(KEYINPUT110), .A3(new_n902), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n916), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n894), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n882), .A3(new_n918), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n921), .B1(new_n927), .B2(new_n910), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT44), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT43), .B1(new_n919), .B2(new_n920), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n926), .A2(new_n910), .A3(new_n882), .A4(new_n918), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT44), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n855), .B2(new_n936), .ZN(new_n937));
  AND2_X1   g512(.A1(G160), .A2(G40), .ZN(new_n938));
  AND2_X1   g513(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(G1996), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  XOR2_X1   g516(.A(new_n941), .B(KEYINPUT111), .Z(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  OR2_X1    g518(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(KEYINPUT46), .ZN(new_n945));
  INV_X1    g520(.A(G2067), .ZN(new_n946));
  XNOR2_X1  g521(.A(new_n740), .B(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n797), .ZN(new_n948));
  AOI22_X1  g523(.A1(new_n944), .A2(new_n945), .B1(new_n939), .B2(new_n948), .ZN(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(KEYINPUT47), .ZN(new_n950));
  INV_X1    g525(.A(new_n939), .ZN(new_n951));
  NOR2_X1   g526(.A1(new_n721), .A2(new_n726), .ZN(new_n952));
  OAI21_X1  g527(.A(new_n947), .B1(new_n940), .B2(new_n797), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n939), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n942), .A2(new_n797), .ZN(new_n955));
  AND2_X1   g530(.A1(new_n955), .A2(KEYINPUT112), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n955), .A2(KEYINPUT112), .ZN(new_n957));
  OAI211_X1 g532(.A(new_n952), .B(new_n954), .C1(new_n956), .C2(new_n957), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n741), .A2(new_n946), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n951), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(new_n721), .B(new_n725), .ZN(new_n961));
  OAI221_X1 g536(.A(new_n954), .B1(new_n951), .B2(new_n961), .C1(new_n956), .C2(new_n957), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n706), .A2(new_n708), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n951), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g539(.A(new_n964), .B(KEYINPUT48), .ZN(new_n965));
  NOR2_X1   g540(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n950), .A2(new_n960), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT127), .ZN(new_n968));
  INV_X1    g543(.A(G8), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT113), .B1(new_n851), .B2(new_n936), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT113), .ZN(new_n971));
  AOI211_X1 g546(.A(new_n971), .B(G1384), .C1(new_n849), .C2(new_n850), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT50), .B1(new_n970), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n973), .A2(KEYINPUT117), .A3(new_n938), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT117), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n971), .B1(G164), .B2(G1384), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n504), .A2(new_n507), .A3(KEYINPUT4), .ZN(new_n978));
  AOI21_X1  g553(.A(new_n507), .B1(new_n504), .B2(KEYINPUT4), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n978), .A2(new_n979), .A3(new_n503), .ZN(new_n980));
  OAI211_X1 g555(.A(KEYINPUT113), .B(new_n936), .C1(new_n980), .C2(new_n498), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n976), .B1(new_n977), .B2(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(G160), .A2(G40), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n975), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n851), .A2(new_n976), .A3(new_n936), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n974), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n986), .A2(G2090), .ZN(new_n987));
  NAND4_X1  g562(.A1(new_n852), .A2(new_n854), .A3(KEYINPUT45), .A4(new_n936), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n988), .A2(new_n938), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n851), .A2(new_n936), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n993), .A2(new_n697), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n969), .B1(new_n987), .B2(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(G303), .A2(G8), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n996), .B(KEYINPUT55), .ZN(new_n997));
  INV_X1    g572(.A(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n995), .A2(new_n998), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n983), .B1(KEYINPUT50), .B2(new_n990), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n977), .A2(new_n981), .A3(new_n976), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n1002), .A2(G2090), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n969), .B1(new_n994), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(new_n998), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n938), .A2(new_n977), .A3(new_n981), .ZN(new_n1006));
  INV_X1    g581(.A(G1976), .ZN(new_n1007));
  OAI211_X1 g582(.A(G8), .B(new_n1006), .C1(G288), .C2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT52), .ZN(new_n1009));
  OR3_X1    g584(.A1(new_n580), .A2(G1981), .A3(new_n582), .ZN(new_n1010));
  OAI21_X1  g585(.A(G1981), .B1(new_n580), .B2(new_n582), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(KEYINPUT114), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT114), .ZN(new_n1013));
  NAND3_X1  g588(.A1(G305), .A2(new_n1013), .A3(G1981), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n1012), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1015), .A2(KEYINPUT49), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(KEYINPUT116), .ZN(new_n1017));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1015), .A2(new_n1018), .A3(KEYINPUT49), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT115), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1015), .B2(KEYINPUT49), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1012), .A2(new_n1014), .A3(KEYINPUT115), .A4(new_n1022), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1017), .A2(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1006), .A2(G8), .ZN(new_n1025));
  INV_X1    g600(.A(new_n1025), .ZN(new_n1026));
  INV_X1    g601(.A(new_n1008), .ZN(new_n1027));
  AOI21_X1  g602(.A(KEYINPUT52), .B1(G288), .B2(new_n1007), .ZN(new_n1028));
  AOI22_X1  g603(.A1(new_n1024), .A2(new_n1026), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1005), .A2(new_n1009), .A3(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n999), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT53), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1032), .B1(new_n993), .B2(G2078), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT126), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n938), .B1(new_n991), .B2(new_n990), .ZN(new_n1036));
  AOI21_X1  g611(.A(KEYINPUT45), .B1(new_n977), .B2(new_n981), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1038), .A2(KEYINPUT53), .A3(new_n443), .ZN(new_n1039));
  OAI211_X1 g614(.A(KEYINPUT126), .B(new_n1032), .C1(new_n993), .C2(G2078), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1002), .A2(new_n748), .ZN(new_n1041));
  NAND4_X1  g616(.A1(new_n1035), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1042), .A2(G171), .ZN(new_n1043));
  INV_X1    g618(.A(G1966), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1000), .A2(new_n785), .A3(new_n1001), .ZN(new_n1046));
  AND2_X1   g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1047), .A2(G168), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1045), .A2(G168), .A3(new_n1046), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT51), .B1(new_n1048), .B2(new_n1050), .ZN(new_n1051));
  OR2_X1    g626(.A1(new_n1050), .A2(KEYINPUT51), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT62), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1051), .A2(new_n1052), .A3(new_n1055), .ZN(new_n1056));
  NAND4_X1  g631(.A1(new_n1031), .A2(new_n1043), .A3(new_n1054), .A4(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1021), .A2(new_n1023), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  OAI211_X1 g635(.A(new_n1007), .B(new_n687), .C1(new_n1060), .C2(new_n1025), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1061), .A2(new_n1010), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n1026), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1064), .B(new_n1009), .C1(new_n1060), .C2(new_n1025), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  AOI211_X1 g641(.A(new_n969), .B(new_n997), .C1(new_n994), .C2(new_n1003), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1063), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1057), .A2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n1047), .A2(new_n969), .A3(G286), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1031), .A2(KEYINPUT118), .A3(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1073), .B(new_n1071), .C1(new_n998), .C2(new_n995), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT63), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1072), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1004), .ZN(new_n1079));
  AOI21_X1  g654(.A(new_n998), .B1(new_n1079), .B2(KEYINPUT119), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(KEYINPUT119), .B2(new_n1079), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(KEYINPUT63), .A3(new_n1073), .A4(new_n1071), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1070), .B1(new_n1078), .B2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT121), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n563), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1085), .A2(new_n571), .ZN(new_n1086));
  OAI211_X1 g661(.A(new_n563), .B(new_n570), .C1(new_n1084), .C2(KEYINPUT57), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT122), .B(KEYINPUT56), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1089), .B(new_n442), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n989), .A2(new_n992), .A3(new_n1090), .ZN(new_n1091));
  AND2_X1   g666(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT120), .ZN(new_n1093));
  INV_X1    g668(.A(G1956), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n986), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1093), .B1(new_n986), .B2(new_n1094), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1092), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n986), .A2(new_n1094), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(KEYINPUT120), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n986), .A2(new_n1093), .A3(new_n1094), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1088), .B1(new_n1101), .B2(new_n1091), .ZN(new_n1102));
  INV_X1    g677(.A(new_n1006), .ZN(new_n1103));
  AOI22_X1  g678(.A1(new_n1002), .A2(new_n813), .B1(new_n1103), .B2(new_n946), .ZN(new_n1104));
  NOR2_X1   g679(.A1(new_n1104), .A2(new_n899), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1097), .B1(new_n1102), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(new_n899), .ZN(new_n1109));
  NOR2_X1   g684(.A1(new_n1104), .A2(KEYINPUT60), .ZN(new_n1110));
  NOR2_X1   g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(new_n1091), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n1112), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1113));
  OAI211_X1 g688(.A(KEYINPUT61), .B(new_n1097), .C1(new_n1113), .C2(new_n1088), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  XOR2_X1   g690(.A(KEYINPUT58), .B(G1341), .Z(new_n1116));
  NAND2_X1  g691(.A1(new_n1006), .A2(new_n1116), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n988), .A2(new_n940), .A3(new_n938), .A4(new_n992), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1117), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1119), .A2(new_n549), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1115), .B1(new_n1120), .B2(KEYINPUT59), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(KEYINPUT123), .A3(KEYINPUT59), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n830), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1123));
  INV_X1    g698(.A(KEYINPUT59), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1123), .A2(KEYINPUT124), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT123), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1126), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1121), .A2(new_n1122), .A3(new_n1125), .A4(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1129));
  AOI21_X1  g704(.A(new_n1129), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1088), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1091), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1114), .B(new_n1128), .C1(new_n1133), .C2(KEYINPUT61), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT125), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1111), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1137), .B1(new_n1102), .B2(new_n1130), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1128), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1137), .B1(new_n1101), .B2(new_n1092), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1132), .A2(new_n1131), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1138), .A2(new_n1142), .A3(KEYINPUT125), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1107), .B1(new_n1136), .B2(new_n1143), .ZN(new_n1144));
  XNOR2_X1  g719(.A(G301), .B(KEYINPUT54), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1042), .A2(new_n1145), .ZN(new_n1146));
  NOR3_X1   g721(.A1(new_n937), .A2(new_n1032), .A3(G2078), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1145), .B1(new_n1147), .B2(new_n989), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1035), .A2(new_n1148), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1031), .A2(new_n1146), .A3(new_n1053), .A4(new_n1149), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1083), .B1(new_n1144), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(G290), .A2(G1986), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n951), .B1(new_n963), .B2(new_n1152), .ZN(new_n1153));
  NOR2_X1   g728(.A1(new_n962), .A2(new_n1153), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n968), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n1097), .A2(KEYINPUT61), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1128), .B1(new_n1102), .B2(new_n1156), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT61), .B1(new_n1141), .B2(new_n1097), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n1135), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1111), .ZN(new_n1160));
  NAND3_X1  g735(.A1(new_n1159), .A2(new_n1143), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1150), .B1(new_n1161), .B2(new_n1106), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1077), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1163));
  AOI21_X1  g738(.A(KEYINPUT118), .B1(new_n1031), .B2(new_n1071), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1082), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AND2_X1   g740(.A1(new_n1057), .A2(new_n1069), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1165), .A2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n968), .B(new_n1154), .C1(new_n1162), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  OAI21_X1  g744(.A(new_n967), .B1(new_n1155), .B2(new_n1169), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g745(.A1(G229), .A2(new_n466), .A3(G401), .A4(G227), .ZN(new_n1172));
  NAND3_X1  g746(.A1(new_n932), .A2(new_n884), .A3(new_n1172), .ZN(G225));
  INV_X1    g747(.A(G225), .ZN(G308));
endmodule


