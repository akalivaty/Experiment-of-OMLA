//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 0 1 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:05 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n824, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944;
  XNOR2_X1  g000(.A(G43gat), .B(G50gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT14), .ZN(new_n203));
  NOR3_X1   g002(.A1(new_n203), .A2(G29gat), .A3(G36gat), .ZN(new_n204));
  INV_X1    g003(.A(G29gat), .ZN(new_n205));
  INV_X1    g004(.A(G36gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT14), .B1(new_n205), .B2(new_n206), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n204), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n209), .A2(KEYINPUT15), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n202), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(new_n202), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n210), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(KEYINPUT87), .B(KEYINPUT17), .Z(new_n216));
  NAND3_X1  g015(.A1(new_n213), .A2(new_n215), .A3(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT88), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n213), .A2(new_n215), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(KEYINPUT17), .ZN(new_n221));
  NAND4_X1  g020(.A1(new_n213), .A2(KEYINPUT88), .A3(new_n215), .A4(new_n216), .ZN(new_n222));
  NAND2_X1  g021(.A1(G85gat), .A2(G92gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT7), .ZN(new_n224));
  NAND2_X1  g023(.A1(G99gat), .A2(G106gat), .ZN(new_n225));
  INV_X1    g024(.A(G85gat), .ZN(new_n226));
  INV_X1    g025(.A(G92gat), .ZN(new_n227));
  AOI22_X1  g026(.A1(KEYINPUT8), .A2(new_n225), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n224), .A2(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(G99gat), .B(G106gat), .Z(new_n230));
  OR3_X1    g029(.A1(new_n229), .A2(KEYINPUT94), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n230), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT94), .B1(new_n229), .B2(new_n230), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n231), .A2(new_n232), .A3(new_n233), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n221), .A3(new_n222), .A4(new_n234), .ZN(new_n235));
  NOR2_X1   g034(.A1(new_n220), .A2(new_n234), .ZN(new_n236));
  AND3_X1   g035(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(G190gat), .B(G218gat), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n239), .B(KEYINPUT95), .Z(new_n240));
  NAND3_X1  g039(.A1(new_n235), .A2(new_n238), .A3(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n240), .B1(new_n235), .B2(new_n238), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT96), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n235), .A2(new_n238), .ZN(new_n245));
  INV_X1    g044(.A(new_n240), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT96), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n247), .A2(new_n248), .A3(new_n241), .ZN(new_n249));
  XNOR2_X1  g048(.A(G134gat), .B(G162gat), .ZN(new_n250));
  AOI21_X1  g049(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n250), .B(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n244), .A2(new_n249), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(new_n252), .ZN(new_n254));
  OAI211_X1 g053(.A(KEYINPUT96), .B(new_n254), .C1(new_n242), .C2(new_n243), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G64gat), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n257), .A2(G57gat), .ZN(new_n258));
  AND2_X1   g057(.A1(new_n257), .A2(G57gat), .ZN(new_n259));
  INV_X1    g058(.A(G71gat), .ZN(new_n260));
  INV_X1    g059(.A(G78gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n258), .A2(new_n259), .B1(new_n262), .B2(KEYINPUT9), .ZN(new_n263));
  XOR2_X1   g062(.A(G71gat), .B(G78gat), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(new_n263), .B(new_n265), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(KEYINPUT21), .ZN(new_n267));
  XOR2_X1   g066(.A(G15gat), .B(G22gat), .Z(new_n268));
  INV_X1    g067(.A(G1gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(G8gat), .B1(new_n270), .B2(KEYINPUT89), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT16), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n272), .A2(G1gat), .ZN(new_n273));
  OAI21_X1  g072(.A(new_n270), .B1(new_n273), .B2(new_n268), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n271), .B(new_n274), .ZN(new_n275));
  XNOR2_X1  g074(.A(G127gat), .B(G155gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n266), .A2(KEYINPUT21), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n275), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G231gat), .A2(G233gat), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n275), .B2(new_n278), .ZN(new_n282));
  NOR3_X1   g081(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n275), .A2(new_n278), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n276), .ZN(new_n285));
  AOI22_X1  g084(.A1(new_n285), .A2(new_n279), .B1(G231gat), .B2(G233gat), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n267), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n281), .B1(new_n280), .B2(new_n282), .ZN(new_n288));
  NAND4_X1  g087(.A1(new_n285), .A2(G231gat), .A3(G233gat), .A4(new_n279), .ZN(new_n289));
  OAI211_X1 g088(.A(new_n288), .B(new_n289), .C1(KEYINPUT21), .C2(new_n266), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g090(.A(G183gat), .B(G211gat), .Z(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  XOR2_X1   g093(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n295));
  XOR2_X1   g094(.A(new_n294), .B(new_n295), .Z(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n291), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n287), .A2(new_n290), .A3(new_n296), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n256), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n301), .A2(KEYINPUT97), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT97), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n256), .A2(new_n300), .A3(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(G230gat), .ZN(new_n305));
  INV_X1    g104(.A(G233gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(new_n263), .B(new_n264), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n231), .A2(new_n309), .A3(new_n232), .A4(new_n233), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT98), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n229), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n230), .ZN(new_n313));
  INV_X1    g112(.A(new_n230), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n229), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n266), .A2(new_n313), .A3(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT10), .B1(new_n310), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n266), .A2(KEYINPUT10), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n234), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n308), .B1(new_n317), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n310), .A2(new_n307), .A3(new_n316), .ZN(new_n321));
  XNOR2_X1  g120(.A(G120gat), .B(G148gat), .ZN(new_n322));
  INV_X1    g121(.A(G176gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(G204gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n320), .A2(new_n321), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(KEYINPUT99), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n320), .A2(new_n321), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n330), .A2(new_n326), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n329), .B(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n302), .A2(new_n304), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT100), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n302), .A2(KEYINPUT100), .A3(new_n304), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT36), .ZN(new_n339));
  INV_X1    g138(.A(G227gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n340), .A2(new_n306), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  NOR2_X1   g141(.A1(G183gat), .A2(G190gat), .ZN(new_n343));
  AND2_X1   g142(.A1(G183gat), .A2(G190gat), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n343), .B1(new_n344), .B2(KEYINPUT24), .ZN(new_n345));
  NAND2_X1  g144(.A1(G183gat), .A2(G190gat), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT24), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT64), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n346), .A2(KEYINPUT64), .A3(new_n347), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n345), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NOR2_X1   g151(.A1(G169gat), .A2(G176gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n353), .A2(KEYINPUT23), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n355), .A2(new_n323), .ZN(new_n356));
  NOR2_X1   g155(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(KEYINPUT23), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n352), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(KEYINPUT25), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT65), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n353), .B(KEYINPUT66), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n345), .A2(new_n348), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n364), .A2(KEYINPUT25), .A3(new_n357), .A4(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT65), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n359), .A2(new_n367), .A3(new_n360), .ZN(new_n368));
  NAND3_X1  g167(.A1(new_n362), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT68), .ZN(new_n370));
  AND2_X1   g169(.A1(G127gat), .A2(G134gat), .ZN(new_n371));
  NOR2_X1   g170(.A1(G127gat), .A2(G134gat), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(G127gat), .ZN(new_n374));
  INV_X1    g173(.A(G134gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(G127gat), .A2(G134gat), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n376), .A2(KEYINPUT68), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n373), .A2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G120gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G113gat), .ZN(new_n381));
  INV_X1    g180(.A(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  AOI21_X1  g182(.A(KEYINPUT1), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(KEYINPUT69), .B1(new_n379), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n384), .B1(new_n372), .B2(new_n371), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n381), .A2(new_n383), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT1), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n389), .A2(new_n390), .A3(new_n373), .A4(new_n378), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n385), .A2(new_n386), .A3(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT26), .ZN(new_n393));
  AOI21_X1  g192(.A(new_n356), .B1(new_n363), .B2(new_n393), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n394), .B1(new_n393), .B2(new_n353), .ZN(new_n395));
  XNOR2_X1  g194(.A(KEYINPUT27), .B(G183gat), .ZN(new_n396));
  INV_X1    g195(.A(G190gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT67), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT28), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  OAI211_X1 g200(.A(new_n396), .B(new_n397), .C1(KEYINPUT67), .C2(KEYINPUT28), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n401), .B(new_n402), .C1(new_n399), .C2(new_n400), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n395), .A2(new_n403), .A3(new_n346), .ZN(new_n404));
  AND3_X1   g203(.A1(new_n369), .A2(new_n392), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n392), .B1(new_n369), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n342), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n407), .A2(KEYINPUT34), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT34), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n409), .B(new_n342), .C1(new_n405), .C2(new_n406), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n405), .A2(new_n406), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n414));
  AOI22_X1  g213(.A1(new_n413), .A2(new_n341), .B1(new_n414), .B2(KEYINPUT33), .ZN(new_n415));
  XNOR2_X1  g214(.A(G15gat), .B(G43gat), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n416), .B(KEYINPUT70), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n417), .B(G71gat), .ZN(new_n418));
  INV_X1    g217(.A(G99gat), .ZN(new_n419));
  XNOR2_X1  g218(.A(new_n418), .B(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT71), .B1(new_n415), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n369), .A2(new_n404), .ZN(new_n422));
  INV_X1    g221(.A(new_n392), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n369), .A2(new_n392), .A3(new_n404), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n341), .A3(new_n425), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n426), .B1(KEYINPUT32), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT71), .ZN(new_n429));
  INV_X1    g228(.A(new_n420), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n428), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n421), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n430), .A2(KEYINPUT33), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n426), .A2(new_n433), .A3(KEYINPUT32), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n412), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(new_n434), .ZN(new_n436));
  AOI211_X1 g235(.A(new_n411), .B(new_n436), .C1(new_n421), .C2(new_n431), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n339), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n415), .A2(KEYINPUT71), .A3(new_n420), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n429), .B1(new_n428), .B2(new_n430), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n434), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(new_n411), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n432), .A2(new_n412), .A3(new_n434), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n442), .A2(KEYINPUT36), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n438), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G155gat), .A2(G162gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT2), .ZN(new_n447));
  OR2_X1    g246(.A1(G141gat), .A2(G148gat), .ZN(new_n448));
  NAND2_X1  g247(.A1(G141gat), .A2(G148gat), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  OAI21_X1  g249(.A(KEYINPUT74), .B1(G155gat), .B2(G162gat), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  XNOR2_X1  g251(.A(G155gat), .B(G162gat), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n450), .A2(new_n453), .A3(new_n451), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n455), .A2(KEYINPUT77), .A3(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  AND3_X1   g257(.A1(new_n450), .A2(new_n453), .A3(new_n451), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n453), .B1(new_n450), .B2(new_n451), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n392), .B1(new_n457), .B2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT4), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT78), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n392), .B1(new_n455), .B2(new_n456), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(new_n463), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n461), .A2(new_n457), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n467), .B(KEYINPUT4), .C1(new_n468), .C2(new_n392), .ZN(new_n469));
  NAND3_X1  g268(.A1(new_n464), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT3), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n473), .B1(new_n459), .B2(new_n460), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n474), .A2(KEYINPUT76), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n455), .A2(new_n456), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT76), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n476), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n423), .B1(new_n475), .B2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n455), .A2(KEYINPUT3), .A3(new_n456), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT75), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n480), .B(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n472), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n470), .A2(new_n483), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n392), .B(new_n476), .ZN(new_n485));
  OAI21_X1  g284(.A(KEYINPUT5), .B1(new_n485), .B2(new_n471), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g287(.A(G1gat), .B(G29gat), .ZN(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT0), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(G57gat), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n491), .B(new_n226), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n479), .A2(new_n482), .ZN(new_n493));
  OAI21_X1  g292(.A(new_n463), .B1(new_n468), .B2(new_n392), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n465), .A2(KEYINPUT4), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n493), .A2(new_n494), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n488), .A2(new_n492), .A3(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499));
  INV_X1    g298(.A(new_n492), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n486), .B1(new_n470), .B2(new_n483), .ZN(new_n501));
  INV_X1    g300(.A(new_n497), .ZN(new_n502));
  OAI21_X1  g301(.A(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n498), .A2(new_n499), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n497), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT79), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT6), .A4(new_n500), .ZN(new_n507));
  OAI211_X1 g306(.A(KEYINPUT6), .B(new_n500), .C1(new_n501), .C2(new_n502), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT79), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n504), .A2(new_n507), .A3(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT73), .ZN(new_n511));
  AND2_X1   g310(.A1(G211gat), .A2(G218gat), .ZN(new_n512));
  NOR2_X1   g311(.A1(G211gat), .A2(G218gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G197gat), .B(G204gat), .ZN(new_n516));
  OAI211_X1 g315(.A(new_n515), .B(new_n516), .C1(KEYINPUT22), .C2(new_n512), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n516), .B1(KEYINPUT22), .B2(new_n512), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n514), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT29), .B1(new_n369), .B2(new_n404), .ZN(new_n522));
  AND2_X1   g321(.A1(G226gat), .A2(G233gat), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AND2_X1   g323(.A1(new_n422), .A2(new_n523), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n521), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n422), .A2(new_n523), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(new_n520), .C1(new_n523), .C2(new_n522), .ZN(new_n528));
  XNOR2_X1  g327(.A(G8gat), .B(G36gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n529), .B(KEYINPUT72), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(G64gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G92gat), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n526), .A2(KEYINPUT30), .A3(new_n528), .A4(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n532), .B1(new_n526), .B2(new_n528), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n511), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n526), .A2(new_n528), .ZN(new_n537));
  OAI211_X1 g336(.A(KEYINPUT73), .B(new_n533), .C1(new_n537), .C2(new_n532), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n532), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT30), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n510), .A2(new_n536), .A3(new_n538), .A4(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT81), .B(G106gat), .ZN(new_n543));
  INV_X1    g342(.A(G22gat), .ZN(new_n544));
  INV_X1    g343(.A(G228gat), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n545), .A2(new_n306), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n475), .A2(new_n478), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT29), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n520), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT3), .B1(new_n520), .B2(new_n549), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n461), .A2(new_n457), .ZN(new_n552));
  NOR2_X1   g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n547), .B1(new_n550), .B2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT80), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AOI21_X1  g355(.A(KEYINPUT29), .B1(new_n475), .B2(new_n478), .ZN(new_n557));
  OAI22_X1  g356(.A1(new_n557), .A2(new_n520), .B1(new_n552), .B2(new_n551), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n558), .A2(KEYINPUT80), .A3(new_n547), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  OR2_X1    g359(.A1(new_n551), .A2(new_n476), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n561), .B(new_n546), .C1(new_n557), .C2(new_n520), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n544), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n562), .ZN(new_n564));
  AOI211_X1 g363(.A(G22gat), .B(new_n564), .C1(new_n556), .C2(new_n559), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n543), .B1(new_n563), .B2(new_n565), .ZN(new_n566));
  XNOR2_X1  g365(.A(KEYINPUT31), .B(G50gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n567), .B(G78gat), .ZN(new_n568));
  AND3_X1   g367(.A1(new_n558), .A2(KEYINPUT80), .A3(new_n547), .ZN(new_n569));
  AOI21_X1  g368(.A(KEYINPUT80), .B1(new_n558), .B2(new_n547), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n562), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n571), .A2(G22gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n560), .A2(new_n544), .A3(new_n562), .ZN(new_n573));
  INV_X1    g372(.A(new_n543), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n566), .A2(new_n568), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n568), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n572), .A2(new_n573), .A3(new_n574), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n574), .B1(new_n572), .B2(new_n573), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n577), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n542), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n445), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT82), .ZN(new_n583));
  INV_X1    g382(.A(new_n510), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT37), .ZN(new_n585));
  OR2_X1    g384(.A1(new_n537), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n532), .B1(new_n537), .B2(new_n585), .ZN(new_n587));
  AND3_X1   g386(.A1(new_n586), .A2(KEYINPUT38), .A3(new_n587), .ZN(new_n588));
  OR4_X1    g387(.A1(KEYINPUT84), .A2(new_n524), .A3(new_n525), .A4(new_n521), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n526), .A2(KEYINPUT84), .A3(new_n528), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(KEYINPUT37), .A3(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(KEYINPUT38), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  OAI211_X1 g391(.A(new_n584), .B(new_n539), .C1(new_n588), .C2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n580), .A2(new_n576), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n534), .A2(new_n535), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n541), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n597), .A2(new_n472), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n485), .A2(new_n471), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT39), .A3(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(KEYINPUT83), .B(KEYINPUT39), .ZN(new_n601));
  NAND3_X1  g400(.A1(new_n597), .A2(new_n472), .A3(new_n601), .ZN(new_n602));
  AND3_X1   g401(.A1(new_n600), .A2(new_n492), .A3(new_n602), .ZN(new_n603));
  AOI22_X1  g402(.A1(new_n603), .A2(KEYINPUT40), .B1(new_n500), .B2(new_n505), .ZN(new_n604));
  OAI211_X1 g403(.A(new_n596), .B(new_n604), .C1(KEYINPUT40), .C2(new_n603), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n593), .A2(new_n594), .A3(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT82), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n445), .A2(new_n581), .A3(new_n607), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n583), .A2(new_n606), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n435), .A2(new_n437), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR3_X1   g411(.A1(new_n584), .A2(new_n596), .A3(KEYINPUT35), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT35), .B1(new_n611), .B2(new_n542), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n609), .A2(new_n616), .ZN(new_n617));
  NAND4_X1  g416(.A1(new_n219), .A2(new_n221), .A3(new_n275), .A4(new_n222), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n220), .A2(new_n275), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT90), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT18), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n621), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n220), .B(new_n275), .ZN(new_n625));
  XOR2_X1   g424(.A(new_n620), .B(KEYINPUT13), .Z(new_n626));
  NAND2_X1  g425(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n622), .A2(new_n623), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n618), .A2(new_n619), .A3(new_n620), .A4(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n627), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT86), .ZN(new_n631));
  XNOR2_X1  g430(.A(KEYINPUT85), .B(KEYINPUT11), .ZN(new_n632));
  XNOR2_X1  g431(.A(G113gat), .B(G141gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g433(.A(G169gat), .B(G197gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n631), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n637), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n630), .A2(KEYINPUT86), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g440(.A(KEYINPUT91), .B1(new_n617), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT91), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n643), .B(new_n644), .C1(new_n609), .C2(new_n616), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n338), .B1(new_n642), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  OAI211_X1 g447(.A(KEYINPUT101), .B(new_n338), .C1(new_n642), .C2(new_n645), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n584), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G1gat), .ZN(G1324gat));
  INV_X1    g451(.A(KEYINPUT42), .ZN(new_n653));
  XNOR2_X1  g452(.A(KEYINPUT102), .B(G8gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(new_n272), .ZN(new_n655));
  AND4_X1   g454(.A1(new_n653), .A2(new_n650), .A3(new_n596), .A4(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n644), .B1(new_n609), .B2(new_n616), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n657), .B(KEYINPUT91), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n658), .B2(new_n338), .ZN(new_n659));
  INV_X1    g458(.A(new_n649), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n596), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n653), .B1(new_n661), .B2(G8gat), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n650), .A2(new_n596), .A3(new_n655), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n656), .B1(new_n662), .B2(new_n663), .ZN(G1325gat));
  AOI21_X1  g463(.A(G15gat), .B1(new_n650), .B2(new_n610), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n445), .B1(new_n648), .B2(new_n649), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n665), .B1(G15gat), .B2(new_n666), .ZN(G1326gat));
  NOR3_X1   g466(.A1(new_n578), .A2(new_n579), .A3(new_n577), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n568), .B1(new_n566), .B2(new_n575), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n650), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT43), .B(G22gat), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n671), .B(new_n672), .ZN(G1327gat));
  NOR2_X1   g472(.A1(new_n642), .A2(new_n645), .ZN(new_n674));
  INV_X1    g473(.A(new_n300), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n333), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n256), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n205), .A3(new_n584), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(new_n256), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n617), .A2(KEYINPUT44), .A3(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n445), .A2(new_n581), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n614), .A2(new_n615), .B1(new_n685), .B2(new_n606), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n684), .B1(new_n686), .B2(new_n256), .ZN(new_n687));
  AND2_X1   g486(.A1(new_n683), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n644), .A2(new_n676), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  OAI21_X1  g489(.A(G29gat), .B1(new_n690), .B2(new_n510), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n681), .A2(new_n691), .ZN(G1328gat));
  NAND3_X1  g491(.A1(new_n679), .A2(new_n206), .A3(new_n596), .ZN(new_n693));
  OR2_X1    g492(.A1(new_n693), .A2(KEYINPUT46), .ZN(new_n694));
  INV_X1    g493(.A(new_n596), .ZN(new_n695));
  OAI21_X1  g494(.A(G36gat), .B1(new_n690), .B2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(KEYINPUT46), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n694), .A2(new_n696), .A3(new_n697), .ZN(G1329gat));
  OAI21_X1  g497(.A(G43gat), .B1(new_n690), .B2(new_n445), .ZN(new_n699));
  INV_X1    g498(.A(new_n679), .ZN(new_n700));
  INV_X1    g499(.A(new_n610), .ZN(new_n701));
  OR2_X1    g500(.A1(new_n701), .A2(G43gat), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n699), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT47), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n699), .B(KEYINPUT47), .C1(new_n700), .C2(new_n702), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(G1330gat));
  NAND4_X1  g506(.A1(new_n683), .A2(new_n670), .A3(new_n687), .A4(new_n689), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G50gat), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n594), .A2(G50gat), .ZN(new_n710));
  OAI211_X1 g509(.A(new_n677), .B(new_n710), .C1(new_n642), .C2(new_n645), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n709), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT48), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT104), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n709), .B1(new_n711), .B2(KEYINPUT103), .ZN(new_n716));
  INV_X1    g515(.A(new_n716), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n713), .B1(new_n711), .B2(KEYINPUT103), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  INV_X1    g518(.A(new_n718), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n716), .A3(KEYINPUT104), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n714), .B1(new_n719), .B2(new_n721), .ZN(G1331gat));
  AND3_X1   g521(.A1(new_n256), .A2(new_n300), .A3(new_n303), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n303), .B1(new_n256), .B2(new_n300), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n725), .A2(new_n332), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n686), .A2(new_n641), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(new_n584), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g528(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(new_n596), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT105), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n732), .B(new_n733), .Z(G1333gat));
  AND2_X1   g533(.A1(new_n727), .A2(new_n610), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n735), .A2(KEYINPUT106), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n736), .A2(new_n260), .A3(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(new_n445), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n727), .A2(G71gat), .A3(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT50), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT50), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n738), .A2(new_n743), .A3(new_n740), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n742), .A2(new_n744), .ZN(G1334gat));
  NAND2_X1  g544(.A1(new_n727), .A2(new_n670), .ZN(new_n746));
  XOR2_X1   g545(.A(KEYINPUT107), .B(G78gat), .Z(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1335gat));
  NOR2_X1   g547(.A1(new_n686), .A2(new_n256), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n641), .A2(new_n300), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT51), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT51), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n749), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n752), .A2(new_n332), .A3(new_n754), .ZN(new_n755));
  OR2_X1    g554(.A1(new_n755), .A2(G85gat), .ZN(new_n756));
  AND4_X1   g555(.A1(new_n584), .A2(new_n688), .A3(new_n332), .A4(new_n750), .ZN(new_n757));
  OAI22_X1  g556(.A1(new_n756), .A2(new_n510), .B1(new_n757), .B2(new_n226), .ZN(G1336gat));
  NAND4_X1  g557(.A1(new_n752), .A2(new_n227), .A3(new_n332), .A4(new_n754), .ZN(new_n759));
  OR2_X1    g558(.A1(new_n759), .A2(new_n695), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n688), .A2(new_n332), .A3(new_n750), .ZN(new_n761));
  OAI21_X1  g560(.A(G92gat), .B1(new_n761), .B2(new_n695), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  OAI21_X1  g562(.A(KEYINPUT108), .B1(new_n759), .B2(new_n695), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(KEYINPUT52), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n760), .B(new_n762), .C1(KEYINPUT108), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n765), .A2(new_n767), .ZN(G1337gat));
  NAND2_X1  g567(.A1(new_n739), .A2(G99gat), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n761), .A2(new_n769), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n419), .B1(new_n755), .B2(new_n701), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT109), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT109), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(new_n774), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1338gat));
  NAND2_X1  g575(.A1(new_n670), .A2(G106gat), .ZN(new_n777));
  OR2_X1    g576(.A1(new_n761), .A2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(G106gat), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n779), .B1(new_n755), .B2(new_n594), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n778), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n778), .A2(KEYINPUT53), .A3(new_n780), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(G1339gat));
  NOR3_X1   g584(.A1(new_n317), .A2(new_n319), .A3(new_n308), .ZN(new_n786));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OR2_X1    g587(.A1(new_n787), .A2(KEYINPUT110), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n320), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n320), .B(new_n789), .C1(new_n786), .C2(new_n787), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n327), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n328), .A2(KEYINPUT55), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n795), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n641), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g597(.A1(new_n624), .A2(new_n627), .A3(new_n629), .A4(new_n637), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n620), .B1(new_n618), .B2(new_n619), .ZN(new_n800));
  NOR2_X1   g599(.A1(new_n625), .A2(new_n626), .ZN(new_n801));
  OAI21_X1  g600(.A(new_n636), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n332), .A2(new_n799), .A3(new_n802), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n682), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n682), .A2(new_n797), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n799), .A2(new_n802), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT111), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n675), .B1(new_n804), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n725), .A2(new_n644), .A3(new_n333), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n596), .A2(new_n510), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n612), .A3(new_n813), .ZN(new_n814));
  XOR2_X1   g613(.A(new_n814), .B(KEYINPUT112), .Z(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n382), .A3(new_n641), .ZN(new_n816));
  OAI21_X1  g615(.A(G113gat), .B1(new_n814), .B2(new_n644), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1340gat));
  NAND2_X1  g617(.A1(new_n332), .A2(new_n380), .ZN(new_n819));
  XOR2_X1   g618(.A(new_n819), .B(KEYINPUT113), .Z(new_n820));
  NAND2_X1  g619(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G120gat), .B1(new_n814), .B2(new_n333), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1341gat));
  NOR2_X1   g622(.A1(new_n814), .A2(new_n675), .ZN(new_n824));
  XNOR2_X1  g623(.A(KEYINPUT114), .B(G127gat), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n824), .B(new_n825), .ZN(G1342gat));
  NOR2_X1   g625(.A1(new_n596), .A2(new_n256), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT115), .ZN(new_n828));
  AND3_X1   g627(.A1(new_n812), .A2(new_n584), .A3(new_n828), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n829), .A2(new_n375), .A3(new_n612), .ZN(new_n830));
  XOR2_X1   g629(.A(new_n830), .B(KEYINPUT56), .Z(new_n831));
  OAI21_X1  g630(.A(G134gat), .B1(new_n814), .B2(new_n256), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(G1343gat));
  AOI21_X1  g632(.A(new_n594), .B1(new_n810), .B2(new_n811), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT57), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n445), .A2(new_n813), .ZN(new_n837));
  INV_X1    g636(.A(new_n837), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT116), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n793), .A2(new_n796), .ZN(new_n840));
  AOI211_X1 g639(.A(KEYINPUT55), .B(new_n327), .C1(new_n791), .C2(new_n792), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n795), .B(KEYINPUT116), .C1(new_n793), .C2(new_n796), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n843), .A3(new_n641), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n682), .B1(new_n844), .B2(new_n803), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n675), .B1(new_n845), .B2(new_n809), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n594), .B1(new_n846), .B2(new_n811), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n836), .B(new_n838), .C1(new_n835), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g647(.A(G141gat), .B1(new_n848), .B2(new_n644), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT58), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n834), .A2(new_n838), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n644), .A2(G141gat), .ZN(new_n853));
  XNOR2_X1  g652(.A(new_n853), .B(KEYINPUT117), .ZN(new_n854));
  OAI221_X1 g653(.A(new_n849), .B1(KEYINPUT118), .B2(new_n850), .C1(new_n852), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(KEYINPUT118), .ZN(new_n856));
  XNOR2_X1  g655(.A(new_n855), .B(new_n856), .ZN(G1344gat));
  OR3_X1    g656(.A1(new_n852), .A2(G148gat), .A3(new_n333), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT120), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n803), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n256), .ZN(new_n862));
  INV_X1    g661(.A(new_n809), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n300), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n641), .B1(new_n336), .B2(new_n337), .ZN(new_n865));
  OAI21_X1  g664(.A(new_n860), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(KEYINPUT100), .B1(new_n725), .B2(new_n333), .ZN(new_n867));
  INV_X1    g666(.A(new_n337), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n644), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(KEYINPUT120), .A3(new_n846), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n866), .A2(new_n870), .A3(new_n670), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n835), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n873));
  AND3_X1   g672(.A1(new_n834), .A2(new_n873), .A3(KEYINPUT57), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n834), .B2(KEYINPUT57), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n872), .A2(new_n876), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n877), .A2(new_n332), .A3(new_n838), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n859), .B1(new_n878), .B2(G148gat), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n859), .B(G148gat), .C1(new_n848), .C2(new_n333), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n858), .B1(new_n879), .B2(new_n881), .ZN(G1345gat));
  OAI21_X1  g681(.A(G155gat), .B1(new_n848), .B2(new_n675), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n675), .A2(G155gat), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n883), .B1(new_n852), .B2(new_n884), .ZN(G1346gat));
  INV_X1    g684(.A(G162gat), .ZN(new_n886));
  NAND4_X1  g685(.A1(new_n829), .A2(new_n886), .A3(new_n670), .A4(new_n445), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n848), .A2(new_n256), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT121), .Z(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n889), .B2(new_n886), .ZN(G1347gat));
  NOR2_X1   g689(.A1(new_n695), .A2(new_n584), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n892), .B1(new_n810), .B2(new_n811), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n893), .A2(new_n612), .ZN(new_n894));
  OAI21_X1  g693(.A(G169gat), .B1(new_n894), .B2(new_n644), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n894), .B(KEYINPUT122), .Z(new_n896));
  NAND2_X1  g695(.A1(new_n641), .A2(new_n355), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n895), .B1(new_n896), .B2(new_n897), .ZN(G1348gat));
  INV_X1    g697(.A(new_n896), .ZN(new_n899));
  AOI21_X1  g698(.A(G176gat), .B1(new_n899), .B2(new_n332), .ZN(new_n900));
  AND2_X1   g699(.A1(new_n900), .A2(KEYINPUT123), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n900), .A2(KEYINPUT123), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n894), .A2(new_n323), .A3(new_n333), .ZN(new_n903));
  XNOR2_X1  g702(.A(new_n903), .B(KEYINPUT124), .ZN(new_n904));
  NOR3_X1   g703(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(G1349gat));
  NOR2_X1   g704(.A1(new_n894), .A2(new_n675), .ZN(new_n906));
  MUX2_X1   g705(.A(G183gat), .B(new_n396), .S(new_n906), .Z(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g707(.A1(new_n899), .A2(new_n397), .A3(new_n682), .ZN(new_n909));
  OAI21_X1  g708(.A(G190gat), .B1(new_n894), .B2(new_n256), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n911));
  INV_X1    g710(.A(new_n911), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT61), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n910), .A2(KEYINPUT125), .ZN(new_n914));
  AND3_X1   g713(.A1(new_n912), .A2(new_n913), .A3(new_n914), .ZN(new_n915));
  AOI21_X1  g714(.A(new_n913), .B1(new_n912), .B2(new_n914), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n909), .B1(new_n915), .B2(new_n916), .ZN(G1351gat));
  NOR2_X1   g716(.A1(new_n739), .A2(new_n892), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n834), .A2(new_n918), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  INV_X1    g719(.A(G197gat), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n641), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n872), .A2(new_n876), .ZN(new_n923));
  INV_X1    g722(.A(new_n918), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(new_n644), .A3(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n922), .B1(new_n925), .B2(new_n921), .ZN(G1352gat));
  NOR3_X1   g725(.A1(new_n919), .A2(G204gat), .A3(new_n333), .ZN(new_n927));
  XNOR2_X1  g726(.A(new_n927), .B(KEYINPUT62), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n923), .A2(new_n333), .A3(new_n924), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n928), .B1(new_n929), .B2(new_n325), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n877), .A2(new_n300), .A3(new_n918), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT127), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT127), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n877), .A2(new_n933), .A3(new_n300), .A4(new_n918), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n932), .A2(G211gat), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT63), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT63), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n932), .A2(new_n937), .A3(G211gat), .A4(new_n934), .ZN(new_n938));
  NOR3_X1   g737(.A1(new_n919), .A2(G211gat), .A3(new_n675), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT126), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n938), .A3(new_n940), .ZN(G1354gat));
  AOI21_X1  g740(.A(G218gat), .B1(new_n920), .B2(new_n682), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n923), .A2(new_n924), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n682), .A2(G218gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(G1355gat));
endmodule


