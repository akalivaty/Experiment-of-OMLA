//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 1 1 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 1 1 0 1 0 1 0 1 1 0 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n802, new_n803, new_n804, new_n806, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n819, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n955, new_n956, new_n957, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030;
  INV_X1    g000(.A(KEYINPUT85), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT4), .ZN(new_n203));
  INV_X1    g002(.A(G134gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G127gat), .ZN(new_n205));
  INV_X1    g004(.A(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(G134gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n205), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G113gat), .B(G120gat), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n208), .B1(new_n209), .B2(KEYINPUT1), .ZN(new_n210));
  INV_X1    g009(.A(G120gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n211), .A2(G113gat), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT70), .B(G120gat), .ZN(new_n213));
  AOI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(G113gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT1), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n205), .A2(new_n207), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n210), .B1(new_n214), .B2(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G155gat), .A2(G162gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G155gat), .A2(G162gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(G141gat), .B(G148gat), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT2), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n222), .B1(G155gat), .B2(G162gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G141gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(G148gat), .ZN(new_n226));
  INV_X1    g025(.A(G148gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G141gat), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n226), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(G155gat), .B(G162gat), .ZN(new_n230));
  INV_X1    g029(.A(G155gat), .ZN(new_n231));
  INV_X1    g030(.A(G162gat), .ZN(new_n232));
  OAI21_X1  g031(.A(KEYINPUT2), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n229), .A2(new_n230), .A3(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n224), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n203), .B1(new_n217), .B2(new_n235), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n224), .A2(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n211), .A2(KEYINPUT70), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT70), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(G120gat), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n238), .A2(new_n240), .A3(G113gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n212), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n216), .ZN(new_n244));
  INV_X1    g043(.A(G113gat), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n245), .A2(G120gat), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n215), .B1(new_n212), .B2(new_n246), .ZN(new_n247));
  AOI22_X1  g046(.A1(new_n243), .A2(new_n244), .B1(new_n247), .B2(new_n208), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n237), .A2(new_n248), .A3(KEYINPUT4), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n236), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n237), .A2(new_n248), .ZN(new_n251));
  NAND2_X1  g050(.A1(G225gat), .A2(G233gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n243), .A2(new_n244), .ZN(new_n255));
  AOI22_X1  g054(.A1(KEYINPUT3), .A2(new_n235), .B1(new_n255), .B2(new_n210), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT3), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n224), .A2(new_n234), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT79), .B1(new_n256), .B2(new_n258), .ZN(new_n259));
  NOR3_X1   g058(.A1(new_n220), .A2(new_n221), .A3(new_n223), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n230), .B1(new_n233), .B2(new_n229), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT3), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND4_X1   g061(.A1(KEYINPUT79), .A2(new_n262), .A3(new_n217), .A4(new_n258), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n250), .B(new_n254), .C1(new_n259), .C2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT5), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n217), .A2(new_n235), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n251), .A2(new_n266), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n265), .B1(new_n267), .B2(new_n253), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n236), .A2(new_n249), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n262), .A2(new_n217), .A3(new_n258), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT79), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n256), .A2(KEYINPUT79), .A3(new_n258), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n269), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n253), .A2(KEYINPUT5), .ZN(new_n275));
  AOI22_X1  g074(.A1(new_n264), .A2(new_n268), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G1gat), .B(G29gat), .ZN(new_n277));
  XNOR2_X1  g076(.A(new_n277), .B(KEYINPUT0), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(G57gat), .ZN(new_n279));
  INV_X1    g078(.A(G85gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(new_n279), .B(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(new_n202), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n274), .A2(new_n252), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT84), .B1(new_n267), .B2(new_n253), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT84), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n251), .A2(new_n266), .A3(new_n285), .A4(new_n252), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n284), .A2(KEYINPUT39), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n281), .B1(new_n283), .B2(new_n287), .ZN(new_n288));
  NOR3_X1   g087(.A1(new_n274), .A2(KEYINPUT39), .A3(new_n252), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT40), .ZN(new_n291));
  INV_X1    g090(.A(new_n281), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n267), .A2(new_n253), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT5), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n294), .B1(new_n274), .B2(new_n254), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n250), .B(new_n275), .C1(new_n259), .C2(new_n263), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(KEYINPUT85), .B(new_n292), .C1(new_n295), .C2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT40), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n288), .B2(new_n289), .ZN(new_n300));
  AND4_X1   g099(.A1(new_n282), .A2(new_n291), .A3(new_n298), .A4(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(G64gat), .B(G92gat), .ZN(new_n302));
  XNOR2_X1  g101(.A(new_n302), .B(G36gat), .ZN(new_n303));
  XNOR2_X1  g102(.A(KEYINPUT78), .B(G8gat), .ZN(new_n304));
  XOR2_X1   g103(.A(new_n303), .B(new_n304), .Z(new_n305));
  INV_X1    g104(.A(G226gat), .ZN(new_n306));
  INV_X1    g105(.A(G233gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT29), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(G169gat), .ZN(new_n312));
  INV_X1    g111(.A(G176gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT66), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  NOR2_X1   g115(.A1(G169gat), .A2(G176gat), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT66), .ZN(new_n318));
  NOR3_X1   g117(.A1(new_n317), .A2(new_n318), .A3(KEYINPUT23), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT25), .ZN(new_n321));
  NAND2_X1  g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT68), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n321), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT23), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n324), .B(new_n325), .C1(new_n323), .C2(new_n322), .ZN(new_n326));
  NOR2_X1   g125(.A1(G183gat), .A2(G190gat), .ZN(new_n327));
  INV_X1    g126(.A(G183gat), .ZN(new_n328));
  INV_X1    g127(.A(G190gat), .ZN(new_n329));
  OAI21_X1  g128(.A(KEYINPUT24), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT24), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n331), .A2(G183gat), .A3(G190gat), .ZN(new_n332));
  AOI21_X1  g131(.A(new_n327), .B1(new_n330), .B2(new_n332), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n320), .A2(new_n326), .A3(new_n333), .ZN(new_n334));
  AND2_X1   g133(.A1(G169gat), .A2(G176gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(KEYINPUT23), .B2(new_n317), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n336), .B1(new_n316), .B2(new_n319), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT67), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT67), .ZN(new_n339));
  OAI211_X1 g138(.A(new_n339), .B(new_n336), .C1(new_n316), .C2(new_n319), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT65), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n327), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n330), .A2(new_n332), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n338), .A2(new_n340), .A3(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n346));
  AOI21_X1  g145(.A(new_n334), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n348));
  OR2_X1    g147(.A1(new_n328), .A2(KEYINPUT27), .ZN(new_n349));
  AND2_X1   g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT28), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n350), .A2(new_n351), .A3(new_n329), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n329), .A3(new_n348), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n314), .A2(KEYINPUT26), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT26), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n322), .B1(new_n317), .B2(new_n357), .ZN(new_n358));
  OAI22_X1  g157(.A1(new_n356), .A2(new_n358), .B1(new_n328), .B2(new_n329), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(KEYINPUT69), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT69), .ZN(new_n361));
  OAI221_X1 g160(.A(new_n361), .B1(new_n328), .B2(new_n329), .C1(new_n356), .C2(new_n358), .ZN(new_n362));
  AOI21_X1  g161(.A(new_n355), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  OAI21_X1  g162(.A(new_n311), .B1(new_n347), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g163(.A(G197gat), .B(G204gat), .ZN(new_n365));
  INV_X1    g164(.A(G211gat), .ZN(new_n366));
  INV_X1    g165(.A(G218gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n365), .B1(KEYINPUT22), .B2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G211gat), .B(G218gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n360), .A2(new_n362), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n354), .A3(new_n352), .ZN(new_n374));
  INV_X1    g173(.A(new_n346), .ZN(new_n375));
  AOI22_X1  g174(.A1(new_n337), .A2(KEYINPUT67), .B1(new_n343), .B2(new_n342), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(new_n340), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n374), .B(new_n309), .C1(new_n377), .C2(new_n334), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n364), .A2(new_n372), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT76), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n372), .B1(new_n364), .B2(new_n378), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n325), .A2(new_n322), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n318), .B1(new_n317), .B2(KEYINPUT23), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n314), .A2(KEYINPUT66), .A3(new_n315), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n384), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n344), .B1(new_n387), .B2(new_n339), .ZN(new_n388));
  INV_X1    g187(.A(new_n340), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n346), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n334), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n392), .A2(new_n374), .B1(new_n310), .B2(new_n309), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n347), .A2(new_n363), .A3(new_n308), .ZN(new_n394));
  OAI211_X1 g193(.A(KEYINPUT76), .B(new_n371), .C1(new_n393), .C2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n305), .B1(new_n383), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n371), .B1(new_n393), .B2(new_n394), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n400), .A2(new_n380), .A3(new_n379), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n395), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n402), .A2(KEYINPUT30), .A3(new_n305), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT77), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n401), .A2(KEYINPUT77), .A3(new_n395), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n305), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n301), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(G228gat), .A2(G233gat), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n257), .B1(new_n371), .B2(KEYINPUT29), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n235), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n410), .B1(new_n412), .B2(KEYINPUT81), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n258), .A2(new_n310), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n371), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n412), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n413), .A2(new_n416), .ZN(new_n417));
  OAI211_X1 g216(.A(new_n412), .B(new_n415), .C1(KEYINPUT81), .C2(new_n410), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(G22gat), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n420), .A2(KEYINPUT82), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(G22gat), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n419), .A2(new_n421), .A3(new_n423), .ZN(new_n424));
  NAND4_X1  g223(.A1(new_n417), .A2(new_n422), .A3(G22gat), .A4(new_n418), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(KEYINPUT80), .A3(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(KEYINPUT83), .A2(G22gat), .ZN(new_n427));
  AND3_X1   g226(.A1(new_n417), .A2(new_n418), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n427), .B1(new_n417), .B2(new_n418), .ZN(new_n429));
  XNOR2_X1  g228(.A(G78gat), .B(G106gat), .ZN(new_n430));
  XNOR2_X1  g229(.A(new_n430), .B(KEYINPUT31), .ZN(new_n431));
  INV_X1    g230(.A(G50gat), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n428), .A2(new_n429), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT80), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n424), .A2(new_n435), .A3(new_n425), .ZN(new_n436));
  AOI22_X1  g235(.A1(new_n426), .A2(new_n434), .B1(new_n436), .B2(new_n433), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT38), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n401), .A2(KEYINPUT77), .A3(new_n395), .ZN(new_n439));
  AOI21_X1  g238(.A(KEYINPUT77), .B1(new_n401), .B2(new_n395), .ZN(new_n440));
  OAI21_X1  g239(.A(KEYINPUT37), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT37), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n442), .B1(new_n383), .B2(new_n396), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n438), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n305), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(new_n438), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n400), .A2(KEYINPUT87), .A3(new_n379), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT87), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n442), .B1(new_n382), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n446), .B1(new_n447), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n401), .A2(new_n438), .A3(new_n395), .ZN(new_n451));
  AOI22_X1  g250(.A1(new_n443), .A2(new_n450), .B1(new_n451), .B2(new_n305), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n292), .B1(new_n295), .B2(new_n297), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT6), .ZN(new_n454));
  NOR2_X1   g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT6), .B1(new_n276), .B2(new_n281), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n282), .A2(new_n456), .A3(new_n298), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n455), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n282), .A2(new_n456), .A3(KEYINPUT86), .A4(new_n298), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n452), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  OAI211_X1 g260(.A(new_n409), .B(new_n437), .C1(new_n444), .C2(new_n461), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n248), .B1(new_n347), .B2(new_n363), .ZN(new_n463));
  NAND2_X1  g262(.A1(G227gat), .A2(G233gat), .ZN(new_n464));
  INV_X1    g263(.A(new_n464), .ZN(new_n465));
  OAI211_X1 g264(.A(new_n374), .B(new_n217), .C1(new_n377), .C2(new_n334), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  XNOR2_X1  g266(.A(G15gat), .B(G43gat), .ZN(new_n468));
  INV_X1    g267(.A(G71gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(new_n470), .B(KEYINPUT72), .ZN(new_n471));
  OR2_X1    g270(.A1(new_n471), .A2(G99gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT71), .B(KEYINPUT33), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n471), .A2(G99gat), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n472), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n467), .A2(KEYINPUT32), .A3(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n467), .A2(KEYINPUT74), .A3(KEYINPUT32), .A4(new_n476), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n472), .A2(new_n475), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n482), .B1(new_n467), .B2(KEYINPUT32), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n473), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n483), .A2(KEYINPUT73), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT73), .B1(new_n483), .B2(new_n484), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n463), .A2(new_n466), .ZN(new_n488));
  OAI211_X1 g287(.A(KEYINPUT75), .B(KEYINPUT34), .C1(new_n488), .C2(new_n465), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT75), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n465), .B1(new_n463), .B2(new_n466), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT34), .ZN(new_n492));
  OAI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n492), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n489), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NOR2_X1   g295(.A1(new_n487), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n483), .A2(new_n484), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT73), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n483), .A2(KEYINPUT73), .A3(new_n484), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n495), .B1(new_n502), .B2(new_n481), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT36), .B1(new_n497), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n496), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT36), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n495), .B(new_n481), .C1(new_n486), .C2(new_n485), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n445), .B1(new_n439), .B2(new_n440), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n456), .A2(new_n453), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(new_n454), .B2(new_n453), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n509), .A2(new_n511), .A3(new_n399), .A4(new_n403), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n434), .A2(new_n426), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n436), .A2(new_n433), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n512), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n462), .A2(new_n504), .A3(new_n508), .A4(new_n516), .ZN(new_n517));
  AND3_X1   g316(.A1(new_n437), .A2(new_n505), .A3(new_n507), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n509), .A2(new_n399), .A3(new_n403), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT35), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n459), .A2(new_n460), .ZN(new_n521));
  INV_X1    g320(.A(new_n521), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n518), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n437), .A2(new_n505), .A3(new_n507), .ZN(new_n524));
  OAI21_X1  g323(.A(KEYINPUT35), .B1(new_n524), .B2(new_n512), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(KEYINPUT88), .B(KEYINPUT11), .ZN(new_n528));
  XNOR2_X1  g327(.A(G113gat), .B(G141gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(G169gat), .B(G197gat), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  XNOR2_X1  g331(.A(new_n532), .B(KEYINPUT12), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  XNOR2_X1  g333(.A(G15gat), .B(G22gat), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT16), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(G1gat), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n537), .B1(G1gat), .B2(new_n535), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(G8gat), .ZN(new_n539));
  INV_X1    g338(.A(G43gat), .ZN(new_n540));
  OAI21_X1  g339(.A(KEYINPUT15), .B1(new_n540), .B2(G50gat), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n432), .A2(G43gat), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT91), .B(G43gat), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(new_n432), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT92), .B(G50gat), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(new_n540), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT15), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  XOR2_X1   g349(.A(KEYINPUT90), .B(G29gat), .Z(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(G36gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT89), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n553), .A2(G29gat), .A3(G36gat), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n553), .B1(G29gat), .B2(G36gat), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(KEYINPUT14), .ZN(new_n556));
  OR2_X1    g355(.A1(new_n555), .A2(KEYINPUT14), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n544), .B1(new_n550), .B2(new_n558), .ZN(new_n559));
  AND3_X1   g358(.A1(new_n552), .A2(new_n556), .A3(new_n557), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n543), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n539), .B1(new_n562), .B2(KEYINPUT17), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT93), .ZN(new_n564));
  NOR3_X1   g363(.A1(new_n562), .A2(new_n564), .A3(KEYINPUT17), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n558), .A2(new_n544), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n545), .A2(G50gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(KEYINPUT92), .B(G50gat), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n569), .A2(G43gat), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n560), .A2(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n566), .B1(new_n572), .B2(new_n544), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT17), .ZN(new_n574));
  AOI21_X1  g373(.A(KEYINPUT93), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n563), .B1(new_n565), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(G229gat), .A2(G233gat), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n539), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n576), .A2(KEYINPUT18), .A3(new_n577), .A4(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n577), .B(KEYINPUT13), .Z(new_n580));
  OAI21_X1  g379(.A(KEYINPUT94), .B1(new_n573), .B2(new_n539), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(new_n578), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n573), .A2(KEYINPUT94), .A3(new_n539), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n580), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n577), .ZN(new_n586));
  INV_X1    g385(.A(new_n578), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n564), .B1(new_n562), .B2(KEYINPUT17), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n573), .A2(KEYINPUT93), .A3(new_n574), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI211_X1 g389(.A(new_n586), .B(new_n587), .C1(new_n590), .C2(new_n563), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n585), .A2(KEYINPUT95), .B1(KEYINPUT18), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT95), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n579), .B2(new_n584), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n534), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g394(.A(new_n533), .B1(new_n591), .B2(KEYINPUT18), .ZN(new_n596));
  OAI21_X1  g395(.A(KEYINPUT96), .B1(new_n596), .B2(new_n585), .ZN(new_n597));
  AND2_X1   g396(.A1(new_n579), .A2(new_n584), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT96), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n601));
  AOI21_X1  g400(.A(new_n534), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n598), .A2(new_n599), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n595), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G134gat), .B(G162gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  XOR2_X1   g406(.A(G99gat), .B(G106gat), .Z(new_n608));
  OR2_X1    g407(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(KEYINPUT99), .A2(G92gat), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n609), .A2(new_n280), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G85gat), .A2(G92gat), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT7), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n612), .A2(KEYINPUT98), .A3(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G99gat), .A2(G106gat), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT8), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n611), .A2(new_n614), .A3(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT7), .B1(new_n612), .B2(KEYINPUT98), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT98), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n619), .B1(G85gat), .B2(G92gat), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n608), .B1(new_n617), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n617), .A2(new_n621), .A3(new_n608), .ZN(new_n624));
  NOR2_X1   g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n625), .B1(new_n562), .B2(KEYINPUT17), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n590), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(KEYINPUT100), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n590), .A2(KEYINPUT100), .A3(new_n626), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  INV_X1    g432(.A(new_n625), .ZN(new_n634));
  OAI21_X1  g433(.A(new_n633), .B1(new_n634), .B2(new_n562), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n607), .B1(new_n631), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g437(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n639));
  XNOR2_X1  g438(.A(G190gat), .B(G218gat), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n631), .A2(new_n607), .A3(new_n636), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n638), .A2(new_n641), .A3(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(new_n641), .ZN(new_n644));
  AOI211_X1 g443(.A(new_n606), .B(new_n635), .C1(new_n629), .C2(new_n630), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n644), .B1(new_n637), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n643), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(G8gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n538), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT21), .ZN(new_n650));
  XNOR2_X1  g449(.A(G57gat), .B(G64gat), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n652));
  AND2_X1   g451(.A1(G71gat), .A2(G78gat), .ZN(new_n653));
  NOR2_X1   g452(.A1(G71gat), .A2(G78gat), .ZN(new_n654));
  OAI22_X1  g453(.A1(new_n651), .A2(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(KEYINPUT9), .ZN(new_n656));
  NOR2_X1   g455(.A1(new_n656), .A2(new_n651), .ZN(new_n657));
  AND2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n655), .A2(new_n657), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n649), .B1(new_n650), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(G183gat), .ZN(new_n662));
  XNOR2_X1  g461(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n663));
  NAND2_X1  g462(.A1(G231gat), .A2(G233gat), .ZN(new_n664));
  XOR2_X1   g463(.A(new_n663), .B(new_n664), .Z(new_n665));
  XNOR2_X1  g464(.A(new_n662), .B(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n660), .A2(new_n650), .ZN(new_n667));
  XNOR2_X1  g466(.A(G127gat), .B(G155gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(G211gat), .ZN(new_n670));
  OR2_X1    g469(.A1(new_n666), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n666), .A2(new_n670), .ZN(new_n672));
  AND2_X1   g471(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n647), .A2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(G230gat), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n675), .A2(new_n307), .ZN(new_n676));
  INV_X1    g475(.A(new_n676), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n660), .B1(new_n624), .B2(new_n623), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n655), .B(new_n657), .ZN(new_n679));
  INV_X1    g478(.A(new_n624), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n679), .A2(new_n680), .A3(new_n622), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n678), .A2(KEYINPUT101), .A3(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT101), .ZN(new_n683));
  OAI211_X1 g482(.A(new_n660), .B(new_n683), .C1(new_n624), .C2(new_n623), .ZN(new_n684));
  AOI21_X1  g483(.A(KEYINPUT10), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n625), .A2(KEYINPUT10), .A3(new_n679), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n677), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n682), .A2(new_n676), .A3(new_n684), .ZN(new_n689));
  XNOR2_X1  g488(.A(G120gat), .B(G148gat), .ZN(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(G176gat), .ZN(new_n691));
  INV_X1    g490(.A(G204gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n688), .A2(new_n689), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(KEYINPUT102), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT102), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n688), .A2(new_n689), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT103), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n688), .A2(new_n689), .ZN(new_n700));
  INV_X1    g499(.A(new_n693), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AND3_X1   g501(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n699), .B1(new_n698), .B2(new_n702), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g504(.A1(new_n527), .A2(new_n605), .A3(new_n674), .A4(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n511), .B(KEYINPUT104), .Z(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  XOR2_X1   g507(.A(new_n708), .B(G1gat), .Z(G1324gat));
  INV_X1    g508(.A(new_n519), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n706), .A2(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n648), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT105), .ZN(new_n713));
  XOR2_X1   g512(.A(KEYINPUT16), .B(G8gat), .Z(new_n714));
  NAND2_X1  g513(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT42), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1325gat));
  INV_X1    g516(.A(KEYINPUT106), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n506), .B1(new_n505), .B2(new_n507), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n504), .A2(KEYINPUT106), .A3(new_n508), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G15gat), .B1(new_n706), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n497), .A2(new_n503), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OR2_X1    g525(.A1(new_n726), .A2(G15gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n706), .B2(new_n727), .ZN(G1326gat));
  NOR2_X1   g527(.A1(new_n706), .A2(new_n437), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT43), .B(G22gat), .Z(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT107), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n729), .B(new_n731), .ZN(G1327gat));
  AND2_X1   g531(.A1(new_n643), .A2(new_n646), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n733), .B1(new_n517), .B2(new_n526), .ZN(new_n734));
  INV_X1    g533(.A(new_n705), .ZN(new_n735));
  INV_X1    g534(.A(new_n605), .ZN(new_n736));
  INV_X1    g535(.A(new_n673), .ZN(new_n737));
  NOR3_X1   g536(.A1(new_n735), .A2(new_n736), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n739), .A2(new_n551), .A3(new_n707), .ZN(new_n740));
  XNOR2_X1  g539(.A(KEYINPUT108), .B(KEYINPUT45), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n740), .B(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n743));
  AOI211_X1 g542(.A(new_n743), .B(new_n733), .C1(new_n517), .C2(new_n526), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n409), .A2(new_n437), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n444), .A2(new_n461), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n516), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  AOI21_X1  g546(.A(new_n747), .B1(new_n722), .B2(new_n721), .ZN(new_n748));
  INV_X1    g547(.A(new_n526), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n647), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g549(.A(new_n744), .B1(new_n750), .B2(new_n743), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n738), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n551), .B1(new_n752), .B2(new_n707), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n742), .A2(new_n753), .ZN(G1328gat));
  NOR3_X1   g553(.A1(new_n739), .A2(G36gat), .A3(new_n710), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(KEYINPUT46), .ZN(new_n756));
  OAI21_X1  g555(.A(G36gat), .B1(new_n752), .B2(new_n710), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(G1329gat));
  AOI21_X1  g557(.A(new_n442), .B1(new_n406), .B2(new_n407), .ZN(new_n759));
  INV_X1    g558(.A(new_n443), .ZN(new_n760));
  OAI21_X1  g559(.A(KEYINPUT38), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n761), .A2(new_n521), .A3(new_n452), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n515), .B1(new_n519), .B2(new_n301), .ZN(new_n763));
  AOI22_X1  g562(.A1(new_n762), .A2(new_n763), .B1(new_n512), .B2(new_n515), .ZN(new_n764));
  AOI22_X1  g563(.A1(new_n723), .A2(new_n764), .B1(new_n525), .B2(new_n523), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n743), .B1(new_n765), .B2(new_n733), .ZN(new_n766));
  INV_X1    g565(.A(new_n723), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n734), .A2(KEYINPUT44), .ZN(new_n768));
  NAND4_X1  g567(.A1(new_n766), .A2(new_n767), .A3(new_n768), .A4(new_n738), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n546), .ZN(new_n770));
  INV_X1    g569(.A(new_n739), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n726), .A2(new_n546), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT47), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT110), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT109), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n545), .B1(new_n769), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g578(.A1(new_n751), .A2(KEYINPUT109), .A3(new_n767), .A4(new_n738), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n773), .A2(KEYINPUT47), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n777), .B1(new_n781), .B2(new_n783), .ZN(new_n784));
  AOI211_X1 g583(.A(KEYINPUT110), .B(new_n782), .C1(new_n779), .C2(new_n780), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n776), .B1(new_n784), .B2(new_n785), .ZN(G1330gat));
  AOI21_X1  g585(.A(new_n437), .B1(new_n739), .B2(KEYINPUT111), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n787), .B1(KEYINPUT111), .B2(new_n739), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n569), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n751), .A2(new_n515), .A3(new_n548), .A4(new_n738), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g591(.A1(new_n735), .A2(new_n674), .A3(new_n736), .ZN(new_n793));
  NOR2_X1   g592(.A1(new_n765), .A2(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n707), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g596(.A1(new_n794), .A2(new_n519), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n799));
  XOR2_X1   g598(.A(KEYINPUT49), .B(G64gat), .Z(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n798), .B2(new_n800), .ZN(G1333gat));
  NAND3_X1  g600(.A1(new_n794), .A2(new_n469), .A3(new_n725), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n765), .A2(new_n723), .A3(new_n793), .ZN(new_n803));
  OAI21_X1  g602(.A(new_n802), .B1(new_n803), .B2(new_n469), .ZN(new_n804));
  XOR2_X1   g603(.A(new_n804), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g604(.A1(new_n794), .A2(new_n515), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g606(.A1(new_n736), .A2(new_n673), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n647), .B(new_n809), .C1(new_n748), .C2(new_n749), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n765), .A2(new_n733), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(KEYINPUT51), .A3(new_n809), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n705), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n280), .A3(new_n795), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n808), .A2(new_n705), .ZN(new_n817));
  AND3_X1   g616(.A1(new_n766), .A2(new_n768), .A3(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n818), .A2(new_n795), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n280), .B2(new_n819), .ZN(G1336gat));
  NOR2_X1   g619(.A1(new_n710), .A2(G92gat), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n815), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT52), .ZN(new_n823));
  NAND4_X1  g622(.A1(new_n766), .A2(new_n519), .A3(new_n768), .A4(new_n817), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n609), .A2(new_n610), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n823), .A3(new_n826), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT113), .ZN(new_n828));
  NOR2_X1   g627(.A1(KEYINPUT112), .A2(KEYINPUT51), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n813), .B2(new_n809), .ZN(new_n831));
  NOR4_X1   g630(.A1(new_n765), .A2(new_n733), .A3(new_n808), .A4(new_n829), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n735), .B(new_n821), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n826), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n828), .B1(new_n834), .B2(KEYINPUT52), .ZN(new_n835));
  AOI211_X1 g634(.A(KEYINPUT113), .B(new_n823), .C1(new_n833), .C2(new_n826), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n827), .B1(new_n835), .B2(new_n836), .ZN(G1337gat));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n767), .A2(G99gat), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n818), .A2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n814), .ZN(new_n841));
  AOI21_X1  g640(.A(KEYINPUT51), .B1(new_n813), .B2(new_n809), .ZN(new_n842));
  OAI211_X1 g641(.A(new_n725), .B(new_n735), .C1(new_n841), .C2(new_n842), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OAI211_X1 g643(.A(new_n838), .B(new_n840), .C1(new_n844), .C2(G99gat), .ZN(new_n845));
  AOI21_X1  g644(.A(G99gat), .B1(new_n815), .B2(new_n725), .ZN(new_n846));
  INV_X1    g645(.A(new_n840), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT114), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n845), .A2(new_n848), .ZN(G1338gat));
  NAND2_X1  g648(.A1(new_n818), .A2(new_n515), .ZN(new_n850));
  XNOR2_X1  g649(.A(KEYINPUT115), .B(G106gat), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT53), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n705), .A2(G106gat), .A3(new_n437), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n854), .B1(new_n841), .B2(new_n842), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n853), .A3(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n831), .A2(new_n832), .ZN(new_n857));
  AOI22_X1  g656(.A1(new_n857), .A2(new_n854), .B1(new_n850), .B2(new_n851), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n856), .B1(new_n858), .B2(new_n853), .ZN(G1339gat));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860));
  INV_X1    g659(.A(new_n685), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n676), .A3(new_n686), .ZN(new_n862));
  AND3_X1   g661(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n688), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n701), .B1(new_n688), .B2(KEYINPUT54), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n860), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g664(.A1(new_n862), .A2(KEYINPUT54), .A3(new_n688), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n688), .A2(KEYINPUT54), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT55), .A4(new_n701), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n865), .A2(new_n698), .A3(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n605), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n577), .B1(new_n576), .B2(new_n578), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n582), .A2(new_n580), .A3(new_n583), .ZN(new_n872));
  OR2_X1    g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  AOI22_X1  g672(.A1(new_n597), .A2(new_n603), .B1(new_n873), .B2(new_n532), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n874), .B1(new_n703), .B2(new_n704), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n647), .B1(new_n870), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n647), .A2(new_n869), .A3(new_n874), .ZN(new_n877));
  INV_X1    g676(.A(new_n877), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n673), .B1(new_n876), .B2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n674), .A2(new_n736), .A3(new_n705), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n881), .A2(new_n437), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT116), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n726), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n883), .B(new_n515), .C1(new_n879), .C2(new_n880), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n795), .A2(new_n710), .ZN(new_n888));
  NOR4_X1   g687(.A1(new_n887), .A2(new_n245), .A3(new_n736), .A4(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(new_n880), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n873), .A2(new_n532), .ZN(new_n891));
  NOR3_X1   g690(.A1(new_n596), .A2(new_n585), .A3(KEYINPUT96), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n599), .B1(new_n598), .B2(new_n602), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  INV_X1    g693(.A(new_n704), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n698), .A2(new_n699), .A3(new_n702), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n894), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n865), .A2(new_n698), .A3(new_n868), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n604), .B2(new_n595), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n733), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n877), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n890), .B1(new_n901), .B2(new_n673), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n707), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n710), .A3(new_n518), .ZN(new_n904));
  OR2_X1    g703(.A1(new_n904), .A2(new_n736), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n889), .B1(new_n245), .B2(new_n905), .ZN(G1340gat));
  NOR3_X1   g705(.A1(new_n887), .A2(new_n705), .A3(new_n888), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n735), .A2(new_n213), .ZN(new_n908));
  OAI22_X1  g707(.A1(new_n907), .A2(new_n211), .B1(new_n904), .B2(new_n908), .ZN(G1341gat));
  NOR3_X1   g708(.A1(new_n887), .A2(new_n673), .A3(new_n888), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n737), .A2(new_n206), .ZN(new_n911));
  OAI22_X1  g710(.A1(new_n910), .A2(new_n206), .B1(new_n904), .B2(new_n911), .ZN(G1342gat));
  NOR3_X1   g711(.A1(new_n733), .A2(G134gat), .A3(new_n519), .ZN(new_n913));
  NAND4_X1  g712(.A1(new_n881), .A2(new_n518), .A3(new_n795), .A4(new_n913), .ZN(new_n914));
  XOR2_X1   g713(.A(new_n914), .B(KEYINPUT56), .Z(new_n915));
  AOI21_X1  g714(.A(new_n515), .B1(new_n879), .B2(new_n880), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n725), .B1(new_n916), .B2(KEYINPUT116), .ZN(new_n917));
  NOR4_X1   g716(.A1(new_n917), .A2(new_n885), .A3(new_n733), .A4(new_n888), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n915), .B1(new_n918), .B2(new_n204), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(KEYINPUT117), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT117), .ZN(new_n921));
  OAI211_X1 g720(.A(new_n915), .B(new_n921), .C1(new_n204), .C2(new_n918), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(new_n922), .ZN(G1343gat));
  INV_X1    g722(.A(KEYINPUT118), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT58), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n767), .A2(new_n437), .ZN(new_n926));
  NAND4_X1  g725(.A1(new_n881), .A2(new_n926), .A3(new_n710), .A4(new_n795), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n736), .A2(G141gat), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  OAI21_X1  g728(.A(new_n925), .B1(new_n927), .B2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n931), .B1(new_n902), .B2(new_n437), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n881), .A2(KEYINPUT57), .A3(new_n515), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n767), .A2(new_n888), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n934), .A2(new_n605), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n930), .B1(new_n936), .B2(G141gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n924), .A2(KEYINPUT58), .ZN(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NOR2_X1   g738(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  AOI211_X1 g739(.A(new_n938), .B(new_n930), .C1(new_n936), .C2(G141gat), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n940), .A2(new_n941), .ZN(G1344gat));
  NOR3_X1   g741(.A1(new_n927), .A2(G148gat), .A3(new_n705), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT119), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT59), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n946), .B1(new_n932), .B2(new_n933), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n881), .B2(new_n515), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n948), .A2(KEYINPUT120), .ZN(new_n949));
  OAI211_X1 g748(.A(new_n735), .B(new_n935), .C1(new_n947), .C2(new_n949), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n945), .B1(new_n950), .B2(G148gat), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n934), .A2(new_n735), .A3(new_n935), .ZN(new_n952));
  AND3_X1   g751(.A1(new_n952), .A2(new_n945), .A3(G148gat), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n944), .B1(new_n951), .B2(new_n953), .ZN(G1345gat));
  NAND2_X1  g753(.A1(new_n934), .A2(new_n935), .ZN(new_n955));
  OAI21_X1  g754(.A(G155gat), .B1(new_n955), .B2(new_n673), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n737), .A2(new_n231), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n927), .B2(new_n957), .ZN(G1346gat));
  NOR3_X1   g757(.A1(new_n733), .A2(G162gat), .A3(new_n519), .ZN(new_n959));
  NAND3_X1  g758(.A1(new_n903), .A2(new_n926), .A3(new_n959), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT121), .ZN(new_n961));
  OAI21_X1  g760(.A(new_n961), .B1(new_n955), .B2(new_n733), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(G162gat), .ZN(new_n963));
  NOR3_X1   g762(.A1(new_n955), .A2(new_n961), .A3(new_n733), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n960), .B1(new_n963), .B2(new_n964), .ZN(G1347gat));
  NOR4_X1   g764(.A1(new_n902), .A2(new_n710), .A3(new_n524), .A4(new_n795), .ZN(new_n966));
  AOI21_X1  g765(.A(G169gat), .B1(new_n966), .B2(new_n605), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n795), .A2(new_n710), .ZN(new_n968));
  INV_X1    g767(.A(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n887), .A2(new_n969), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n736), .A2(new_n312), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n967), .B1(new_n970), .B2(new_n971), .ZN(G1348gat));
  AOI21_X1  g771(.A(new_n313), .B1(new_n970), .B2(new_n735), .ZN(new_n973));
  AND3_X1   g772(.A1(new_n966), .A2(new_n313), .A3(new_n735), .ZN(new_n974));
  OR2_X1    g773(.A1(new_n973), .A2(new_n974), .ZN(G1349gat));
  NAND3_X1  g774(.A1(new_n966), .A2(new_n350), .A3(new_n737), .ZN(new_n976));
  NOR4_X1   g775(.A1(new_n917), .A2(new_n885), .A3(new_n673), .A4(new_n969), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n976), .B1(new_n977), .B2(new_n328), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n978), .A2(KEYINPUT60), .ZN(new_n979));
  INV_X1    g778(.A(KEYINPUT60), .ZN(new_n980));
  OAI211_X1 g779(.A(new_n976), .B(new_n980), .C1(new_n977), .C2(new_n328), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n979), .A2(new_n981), .ZN(G1350gat));
  INV_X1    g781(.A(KEYINPUT122), .ZN(new_n983));
  NOR4_X1   g782(.A1(new_n917), .A2(new_n885), .A3(new_n733), .A4(new_n969), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n984), .B2(new_n329), .ZN(new_n985));
  NAND4_X1  g784(.A1(new_n884), .A2(new_n647), .A3(new_n886), .A4(new_n968), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n986), .A2(KEYINPUT122), .A3(G190gat), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n985), .A2(KEYINPUT61), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n966), .A2(new_n329), .A3(new_n647), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT61), .ZN(new_n990));
  OAI211_X1 g789(.A(new_n983), .B(new_n990), .C1(new_n984), .C2(new_n329), .ZN(new_n991));
  NAND3_X1  g790(.A1(new_n988), .A2(new_n989), .A3(new_n991), .ZN(G1351gat));
  INV_X1    g791(.A(G197gat), .ZN(new_n993));
  INV_X1    g792(.A(KEYINPUT124), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n767), .A2(new_n994), .A3(new_n969), .ZN(new_n995));
  AOI21_X1  g794(.A(KEYINPUT124), .B1(new_n723), .B2(new_n968), .ZN(new_n996));
  OR3_X1    g795(.A1(new_n995), .A2(KEYINPUT125), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g796(.A(KEYINPUT125), .B1(new_n995), .B2(new_n996), .ZN(new_n998));
  AOI211_X1 g797(.A(new_n993), .B(new_n736), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  OAI21_X1  g798(.A(KEYINPUT123), .B1(new_n947), .B2(new_n949), .ZN(new_n1000));
  AOI211_X1 g799(.A(new_n931), .B(new_n437), .C1(new_n879), .C2(new_n880), .ZN(new_n1001));
  OAI21_X1  g800(.A(KEYINPUT120), .B1(new_n948), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n932), .A2(new_n946), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT123), .ZN(new_n1004));
  NAND3_X1  g803(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n999), .A2(new_n1000), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g805(.A1(new_n902), .A2(new_n795), .ZN(new_n1007));
  NOR3_X1   g806(.A1(new_n767), .A2(new_n710), .A3(new_n437), .ZN(new_n1008));
  NAND2_X1  g807(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(new_n993), .B1(new_n1009), .B2(new_n736), .ZN(new_n1010));
  AND2_X1   g809(.A1(new_n1006), .A2(new_n1010), .ZN(G1352gat));
  AOI21_X1  g810(.A(new_n705), .B1(new_n997), .B2(new_n998), .ZN(new_n1012));
  NAND3_X1  g811(.A1(new_n1000), .A2(new_n1005), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g812(.A1(new_n1013), .A2(G204gat), .ZN(new_n1014));
  NOR3_X1   g813(.A1(new_n1009), .A2(G204gat), .A3(new_n705), .ZN(new_n1015));
  XNOR2_X1  g814(.A(new_n1015), .B(KEYINPUT62), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1014), .A2(new_n1016), .ZN(G1353gat));
  OAI21_X1  g816(.A(new_n737), .B1(new_n995), .B2(new_n996), .ZN(new_n1018));
  AOI21_X1  g817(.A(new_n1018), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1019));
  OR2_X1    g818(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1020));
  OR3_X1    g819(.A1(new_n1019), .A2(new_n366), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g820(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n1022));
  OAI211_X1 g821(.A(new_n1020), .B(new_n1022), .C1(new_n1019), .C2(new_n366), .ZN(new_n1023));
  NAND4_X1  g822(.A1(new_n1007), .A2(new_n366), .A3(new_n737), .A4(new_n1008), .ZN(new_n1024));
  NAND3_X1  g823(.A1(new_n1021), .A2(new_n1023), .A3(new_n1024), .ZN(G1354gat));
  NAND2_X1  g824(.A1(new_n647), .A2(G218gat), .ZN(new_n1026));
  XNOR2_X1  g825(.A(new_n1026), .B(KEYINPUT127), .ZN(new_n1027));
  AOI21_X1  g826(.A(new_n1027), .B1(new_n997), .B2(new_n998), .ZN(new_n1028));
  NAND3_X1  g827(.A1(new_n1000), .A2(new_n1005), .A3(new_n1028), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n367), .B1(new_n1009), .B2(new_n733), .ZN(new_n1030));
  AND2_X1   g829(.A1(new_n1029), .A2(new_n1030), .ZN(G1355gat));
endmodule


