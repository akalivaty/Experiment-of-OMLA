//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 1 0 0 0 1 0 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:53 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n803, new_n804, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n830, new_n831,
    new_n832, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1001, new_n1002;
  XOR2_X1   g000(.A(G1gat), .B(G29gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G57gat), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT86), .B(KEYINPUT0), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT5), .ZN(new_n208));
  NOR2_X1   g007(.A1(G127gat), .A2(G134gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G113gat), .B(G120gat), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n210), .B1(new_n211), .B2(KEYINPUT1), .ZN(new_n212));
  XNOR2_X1  g011(.A(KEYINPUT69), .B(G127gat), .ZN(new_n213));
  INV_X1    g012(.A(G134gat), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(KEYINPUT70), .B1(new_n212), .B2(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G127gat), .ZN(new_n217));
  AND2_X1   g016(.A1(new_n217), .A2(KEYINPUT69), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(KEYINPUT69), .ZN(new_n219));
  OAI21_X1  g018(.A(G134gat), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT1), .ZN(new_n221));
  INV_X1    g020(.A(G120gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n222), .A2(G113gat), .ZN(new_n223));
  INV_X1    g022(.A(G113gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n224), .A2(G120gat), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n221), .B1(new_n223), .B2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT70), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n220), .A2(new_n226), .A3(new_n227), .A4(new_n210), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n216), .A2(new_n228), .ZN(new_n229));
  OR2_X1    g028(.A1(new_n221), .A2(KEYINPUT73), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n221), .A2(KEYINPUT73), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n217), .A2(new_n214), .ZN(new_n232));
  OAI211_X1 g031(.A(new_n230), .B(new_n231), .C1(new_n232), .C2(new_n209), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n222), .A2(KEYINPUT71), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT71), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(G120gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n237), .A3(G113gat), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT72), .ZN(new_n239));
  INV_X1    g038(.A(new_n223), .ZN(new_n240));
  AND3_X1   g039(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n239), .B1(new_n238), .B2(new_n240), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n234), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n229), .A2(new_n243), .ZN(new_n244));
  NAND2_X1  g043(.A1(G155gat), .A2(G162gat), .ZN(new_n245));
  INV_X1    g044(.A(G155gat), .ZN(new_n246));
  INV_X1    g045(.A(G162gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n245), .B1(new_n248), .B2(KEYINPUT2), .ZN(new_n249));
  OR2_X1    g048(.A1(G141gat), .A2(G148gat), .ZN(new_n250));
  INV_X1    g049(.A(KEYINPUT85), .ZN(new_n251));
  NAND2_X1  g050(.A1(G141gat), .A2(G148gat), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n250), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AND2_X1   g052(.A1(G141gat), .A2(G148gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(G141gat), .A2(G148gat), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT85), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n249), .A2(new_n253), .A3(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n258));
  NOR2_X1   g057(.A1(KEYINPUT83), .A2(KEYINPUT2), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n245), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT84), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT84), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n262), .B(new_n245), .C1(new_n258), .C2(new_n259), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n250), .A2(new_n252), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n261), .A2(new_n263), .A3(new_n265), .ZN(new_n266));
  AND3_X1   g065(.A1(new_n246), .A2(new_n247), .A3(KEYINPUT82), .ZN(new_n267));
  AOI21_X1  g066(.A(KEYINPUT82), .B1(new_n246), .B2(new_n247), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n245), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(new_n269), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n266), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n244), .A2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n271), .A2(new_n229), .A3(new_n243), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G225gat), .A2(G233gat), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n208), .B1(new_n275), .B2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n264), .B1(new_n260), .B2(KEYINPUT84), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n269), .B1(new_n281), .B2(new_n263), .ZN(new_n282));
  OAI21_X1  g081(.A(KEYINPUT3), .B1(new_n282), .B2(new_n257), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n280), .A2(new_n244), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n274), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n238), .A2(new_n240), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT72), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n238), .A2(new_n239), .A3(new_n240), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n290), .A2(new_n234), .B1(new_n216), .B2(new_n228), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n291), .A2(KEYINPUT4), .A3(new_n271), .ZN(new_n292));
  NAND4_X1  g091(.A1(new_n284), .A2(new_n286), .A3(new_n292), .A4(new_n276), .ZN(new_n293));
  AND2_X1   g092(.A1(new_n278), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(new_n284), .A2(new_n208), .A3(new_n276), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n286), .A2(new_n292), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n286), .A2(new_n292), .A3(KEYINPUT87), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n295), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n207), .B1(new_n294), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT91), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n295), .ZN(new_n304));
  AND3_X1   g103(.A1(new_n286), .A2(new_n292), .A3(KEYINPUT87), .ZN(new_n305));
  AOI21_X1  g104(.A(KEYINPUT87), .B1(new_n286), .B2(new_n292), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n278), .A2(new_n293), .ZN(new_n308));
  AOI21_X1  g107(.A(new_n206), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT91), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n284), .B1(new_n305), .B2(new_n306), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n277), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n206), .B1(new_n313), .B2(KEYINPUT39), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n276), .B1(new_n315), .B2(new_n284), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT39), .B1(new_n275), .B2(new_n277), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(KEYINPUT90), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT90), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n319), .B(KEYINPUT39), .C1(new_n275), .C2(new_n277), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n316), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(KEYINPUT40), .B1(new_n314), .B2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT39), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n207), .B1(new_n316), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT40), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n313), .A2(new_n318), .A3(new_n320), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n325), .A2(new_n326), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n311), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n330));
  XNOR2_X1  g129(.A(G8gat), .B(G36gat), .ZN(new_n331));
  XNOR2_X1  g130(.A(G64gat), .B(G92gat), .ZN(new_n332));
  XOR2_X1   g131(.A(new_n331), .B(new_n332), .Z(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G197gat), .ZN(new_n335));
  INV_X1    g134(.A(G204gat), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(G197gat), .A2(G204gat), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n340));
  OAI21_X1  g139(.A(KEYINPUT78), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(G211gat), .ZN(new_n342));
  INV_X1    g141(.A(G218gat), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G211gat), .A2(G218gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT77), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n348));
  NAND3_X1  g147(.A1(new_n344), .A2(new_n348), .A3(new_n345), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n347), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT22), .ZN(new_n351));
  AOI22_X1  g150(.A1(new_n337), .A2(new_n338), .B1(new_n351), .B2(new_n345), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT78), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n341), .A2(new_n350), .A3(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n347), .A2(new_n352), .A3(new_n353), .A4(new_n349), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g156(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT67), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  OAI211_X1 g160(.A(KEYINPUT67), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT26), .ZN(new_n363));
  INV_X1    g162(.A(G169gat), .ZN(new_n364));
  INV_X1    g163(.A(G176gat), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n363), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  NAND4_X1  g165(.A1(new_n360), .A2(new_n361), .A3(new_n362), .A4(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(G183gat), .A2(G190gat), .ZN(new_n368));
  AND3_X1   g167(.A1(new_n367), .A2(KEYINPUT68), .A3(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT68), .B1(new_n367), .B2(new_n368), .ZN(new_n370));
  INV_X1    g169(.A(G190gat), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(KEYINPUT66), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(G190gat), .ZN(new_n374));
  INV_X1    g173(.A(G183gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT27), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT27), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(G183gat), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n372), .A2(new_n374), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT28), .ZN(new_n380));
  XNOR2_X1  g179(.A(KEYINPUT66), .B(G190gat), .ZN(new_n381));
  XNOR2_X1  g180(.A(KEYINPUT27), .B(G183gat), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT28), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  NOR3_X1   g184(.A1(new_n369), .A2(new_n370), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n368), .A2(KEYINPUT24), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT24), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n388), .A2(G183gat), .A3(G190gat), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n387), .A2(new_n389), .B1(new_n375), .B2(new_n371), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT23), .ZN(new_n392));
  AOI22_X1  g191(.A1(new_n392), .A2(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT65), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(KEYINPUT23), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n364), .A2(new_n365), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(KEYINPUT64), .B(G169gat), .ZN(new_n399));
  NOR2_X1   g198(.A1(new_n392), .A2(G176gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n391), .A2(new_n398), .A3(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT25), .ZN(new_n403));
  AOI22_X1  g202(.A1(new_n393), .A2(new_n395), .B1(new_n364), .B2(new_n365), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n400), .A2(new_n364), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT25), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n381), .A2(new_n375), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n389), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  AOI22_X1  g209(.A1(new_n402), .A2(new_n403), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  INV_X1    g210(.A(G226gat), .ZN(new_n412));
  INV_X1    g211(.A(G233gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NOR3_X1   g213(.A1(new_n386), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n367), .A2(new_n368), .ZN(new_n416));
  INV_X1    g215(.A(KEYINPUT68), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n379), .A2(KEYINPUT28), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n383), .B1(new_n381), .B2(new_n382), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n367), .A2(KEYINPUT68), .A3(new_n368), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n403), .B1(new_n400), .B2(new_n364), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n410), .A2(new_n398), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n364), .A2(KEYINPUT64), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT64), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(G169gat), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n400), .A2(new_n426), .A3(new_n428), .ZN(new_n429));
  NOR3_X1   g228(.A1(new_n404), .A2(new_n390), .A3(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n425), .B1(new_n430), .B2(KEYINPUT25), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT29), .ZN(new_n432));
  INV_X1    g231(.A(new_n414), .ZN(new_n433));
  AOI22_X1  g232(.A1(new_n423), .A2(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n357), .B1(new_n415), .B2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT79), .ZN(new_n436));
  OAI22_X1  g235(.A1(new_n386), .A2(new_n411), .B1(KEYINPUT29), .B2(new_n414), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n423), .A2(new_n431), .A3(new_n433), .ZN(new_n438));
  INV_X1    g237(.A(new_n357), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n436), .A3(new_n440), .ZN(new_n441));
  OAI211_X1 g240(.A(KEYINPUT79), .B(new_n357), .C1(new_n415), .C2(new_n434), .ZN(new_n442));
  AOI211_X1 g241(.A(new_n330), .B(new_n334), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  AND3_X1   g242(.A1(new_n441), .A2(KEYINPUT80), .A3(new_n442), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT80), .B1(new_n441), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n443), .B1(new_n446), .B2(new_n334), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n441), .A2(new_n442), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n448), .A2(new_n333), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT81), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n448), .A2(KEYINPUT81), .A3(new_n333), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n451), .A2(new_n330), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n447), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n329), .A2(new_n454), .ZN(new_n455));
  OAI211_X1 g254(.A(KEYINPUT6), .B(new_n207), .C1(new_n294), .C2(new_n300), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n456), .B(KEYINPUT92), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT37), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n448), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n440), .ZN(new_n460));
  AOI21_X1  g259(.A(KEYINPUT38), .B1(new_n460), .B2(KEYINPUT37), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n459), .A2(new_n334), .A3(new_n461), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n462), .A2(new_n451), .A3(new_n452), .ZN(new_n463));
  NOR3_X1   g262(.A1(new_n444), .A2(new_n445), .A3(new_n458), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n459), .A2(new_n334), .ZN(new_n465));
  OAI21_X1  g264(.A(KEYINPUT38), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n307), .A2(new_n308), .A3(new_n206), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n303), .A2(new_n467), .A3(new_n468), .A4(new_n310), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n457), .A2(new_n463), .A3(new_n466), .A4(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G78gat), .B(G106gat), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n471), .B(G50gat), .ZN(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n472), .B(new_n473), .ZN(new_n474));
  XOR2_X1   g273(.A(new_n474), .B(KEYINPUT89), .Z(new_n475));
  NAND3_X1  g274(.A1(new_n355), .A2(new_n432), .A3(new_n356), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n476), .A2(new_n279), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(new_n272), .ZN(new_n478));
  AOI21_X1  g277(.A(KEYINPUT29), .B1(new_n271), .B2(new_n279), .ZN(new_n479));
  OAI211_X1 g278(.A(new_n478), .B(G22gat), .C1(new_n439), .C2(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(G22gat), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n479), .A2(new_n439), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n271), .B1(new_n476), .B2(new_n279), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n481), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(G228gat), .A2(G233gat), .ZN(new_n485));
  AND3_X1   g284(.A1(new_n480), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n485), .B1(new_n480), .B2(new_n484), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n475), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n480), .A2(new_n484), .ZN(new_n489));
  AND2_X1   g288(.A1(G228gat), .A2(G233gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n474), .A2(KEYINPUT89), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n480), .A2(new_n484), .A3(new_n485), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n491), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n488), .A2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n455), .A2(new_n470), .A3(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(new_n291), .B1(new_n386), .B2(new_n411), .ZN(new_n498));
  NAND2_X1  g297(.A1(G227gat), .A2(G233gat), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n244), .A2(new_n431), .A3(new_n423), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n498), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT33), .ZN(new_n503));
  XNOR2_X1  g302(.A(G15gat), .B(G43gat), .ZN(new_n504));
  XNOR2_X1  g303(.A(G71gat), .B(G99gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n502), .B(KEYINPUT32), .C1(new_n503), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n506), .B1(new_n502), .B2(KEYINPUT32), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n502), .A2(KEYINPUT74), .A3(new_n503), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT74), .B1(new_n502), .B2(new_n503), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n507), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT75), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT34), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n501), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n499), .ZN(new_n517));
  AOI211_X1 g316(.A(KEYINPUT34), .B(new_n500), .C1(new_n498), .C2(new_n501), .ZN(new_n518));
  NOR2_X1   g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(new_n519), .ZN(new_n520));
  OAI211_X1 g319(.A(KEYINPUT75), .B(new_n507), .C1(new_n510), .C2(new_n511), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  OAI211_X1 g321(.A(new_n519), .B(new_n507), .C1(new_n510), .C2(new_n511), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n522), .A2(KEYINPUT36), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n512), .A2(new_n520), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(KEYINPUT76), .A3(new_n523), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT76), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n527), .A3(new_n520), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n526), .A2(new_n528), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n524), .B1(new_n529), .B2(KEYINPUT36), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n468), .A2(new_n467), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n456), .B1(new_n531), .B2(new_n309), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n495), .B1(new_n454), .B2(new_n533), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n497), .A2(new_n530), .A3(new_n534), .ZN(new_n535));
  INV_X1    g334(.A(new_n454), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n457), .A2(new_n469), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n495), .A2(KEYINPUT35), .ZN(new_n538));
  AND4_X1   g337(.A1(new_n529), .A2(new_n536), .A3(new_n537), .A4(new_n538), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n523), .A2(new_n488), .A3(new_n494), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n522), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT93), .ZN(new_n542));
  AND3_X1   g341(.A1(new_n447), .A2(new_n532), .A3(new_n453), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT93), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n522), .A2(new_n540), .A3(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n542), .A2(new_n543), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT35), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT94), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n539), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n546), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n535), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G8gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n553), .A2(G1gat), .ZN(new_n554));
  INV_X1    g353(.A(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(G1gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT16), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n552), .B1(new_n555), .B2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n558), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n560), .A2(new_n554), .A3(G8gat), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  INV_X1    g361(.A(G29gat), .ZN(new_n563));
  INV_X1    g362(.A(G36gat), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n563), .A2(new_n564), .A3(KEYINPUT14), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G29gat), .B2(G36gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n563), .A2(new_n564), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT96), .ZN(new_n571));
  AND2_X1   g370(.A1(G43gat), .A2(G50gat), .ZN(new_n572));
  NOR2_X1   g371(.A1(G43gat), .A2(G50gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT15), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  OR2_X1    g373(.A1(G43gat), .A2(G50gat), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT15), .ZN(new_n576));
  NAND2_X1  g375(.A1(G43gat), .A2(G50gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n570), .A2(new_n571), .A3(new_n574), .A4(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n574), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n565), .B(new_n567), .C1(new_n563), .C2(new_n564), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT96), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT17), .ZN(new_n584));
  INV_X1    g383(.A(new_n574), .ZN(new_n585));
  OAI22_X1  g384(.A1(new_n568), .A2(KEYINPUT95), .B1(new_n563), .B2(new_n564), .ZN(new_n586));
  AND2_X1   g385(.A1(new_n568), .A2(KEYINPUT95), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n583), .A2(new_n584), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n584), .B1(new_n583), .B2(new_n588), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n562), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n559), .A2(new_n561), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n583), .A2(new_n588), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g394(.A1(new_n591), .A2(new_n592), .A3(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n592), .A4(new_n595), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT97), .B1(new_n593), .B2(new_n594), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT97), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n562), .A2(new_n601), .A3(new_n583), .A4(new_n588), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n595), .A3(new_n602), .ZN(new_n603));
  XOR2_X1   g402(.A(new_n592), .B(KEYINPUT13), .Z(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n598), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(G113gat), .B(G141gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n607), .B(G197gat), .ZN(new_n608));
  XOR2_X1   g407(.A(KEYINPUT11), .B(G169gat), .Z(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT12), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n606), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g412(.A1(new_n596), .A2(new_n597), .B1(new_n604), .B2(new_n603), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n611), .B1(new_n614), .B2(new_n599), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT98), .ZN(new_n616));
  NOR3_X1   g415(.A1(new_n613), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n606), .A2(new_n612), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n614), .A2(new_n611), .A3(new_n599), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT98), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g420(.A(G57gat), .B(G64gat), .Z(new_n622));
  INV_X1    g421(.A(KEYINPUT99), .ZN(new_n623));
  NAND2_X1  g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT9), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n622), .A2(new_n623), .A3(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(G71gat), .B(G78gat), .Z(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NAND4_X1  g429(.A1(new_n630), .A2(new_n623), .A3(new_n626), .A4(new_n622), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  XOR2_X1   g431(.A(KEYINPUT100), .B(KEYINPUT21), .Z(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND2_X1  g433(.A1(G231gat), .A2(G233gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(G127gat), .ZN(new_n637));
  XOR2_X1   g436(.A(G183gat), .B(G211gat), .Z(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT21), .ZN(new_n640));
  OAI21_X1  g439(.A(new_n562), .B1(new_n640), .B2(new_n632), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT101), .ZN(new_n642));
  XNOR2_X1  g441(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(new_n246), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n642), .B(new_n644), .ZN(new_n645));
  OR2_X1    g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n639), .A2(new_n645), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  INV_X1    g447(.A(G85gat), .ZN(new_n649));
  INV_X1    g448(.A(G92gat), .ZN(new_n650));
  OAI21_X1  g449(.A(KEYINPUT7), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT7), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n652), .A2(G85gat), .A3(G92gat), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n650), .A2(KEYINPUT102), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT102), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(G92gat), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n655), .A2(new_n657), .A3(new_n649), .ZN(new_n658));
  NAND2_X1  g457(.A1(G99gat), .A2(G106gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(KEYINPUT8), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n654), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g460(.A(G99gat), .B(G106gat), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(KEYINPUT103), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n661), .A2(new_n662), .ZN(new_n664));
  XNOR2_X1  g463(.A(KEYINPUT102), .B(G92gat), .ZN(new_n665));
  AOI22_X1  g464(.A1(new_n665), .A2(new_n649), .B1(KEYINPUT8), .B2(new_n659), .ZN(new_n666));
  INV_X1    g465(.A(new_n662), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n666), .A2(new_n667), .A3(new_n654), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n664), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  OAI211_X1 g469(.A(new_n663), .B(new_n670), .C1(new_n589), .C2(new_n590), .ZN(new_n671));
  XOR2_X1   g470(.A(G190gat), .B(G218gat), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n670), .A2(new_n663), .ZN(new_n674));
  AND2_X1   g473(.A1(G232gat), .A2(G233gat), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n674), .A2(new_n594), .B1(KEYINPUT41), .B2(new_n675), .ZN(new_n676));
  AND3_X1   g475(.A1(new_n671), .A2(new_n673), .A3(new_n676), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n673), .B1(new_n671), .B2(new_n676), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n675), .A2(KEYINPUT41), .ZN(new_n679));
  XNOR2_X1  g478(.A(G134gat), .B(G162gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  OR3_X1    g481(.A1(new_n677), .A2(new_n678), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n682), .B1(new_n677), .B2(new_n678), .ZN(new_n684));
  AND2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n648), .A2(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n670), .A2(new_n632), .A3(new_n663), .ZN(new_n688));
  INV_X1    g487(.A(KEYINPUT10), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n664), .A2(new_n668), .A3(new_n629), .A4(new_n631), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n688), .A2(new_n689), .A3(new_n690), .ZN(new_n691));
  NAND4_X1  g490(.A1(new_n674), .A2(KEYINPUT10), .A3(new_n629), .A4(new_n631), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g492(.A1(G230gat), .A2(G233gat), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n688), .A2(new_n690), .ZN(new_n696));
  INV_X1    g495(.A(new_n694), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(G120gat), .B(G148gat), .ZN(new_n700));
  XNOR2_X1  g499(.A(G176gat), .B(G204gat), .ZN(new_n701));
  XOR2_X1   g500(.A(new_n700), .B(new_n701), .Z(new_n702));
  INV_X1    g501(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n695), .A2(new_n698), .A3(new_n702), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n687), .A2(new_n706), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n551), .A2(new_n621), .A3(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(new_n533), .ZN(new_n710));
  XNOR2_X1  g509(.A(KEYINPUT104), .B(G1gat), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n710), .B(new_n711), .ZN(G1324gat));
  NOR2_X1   g511(.A1(new_n551), .A2(new_n621), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n708), .A2(new_n536), .ZN(new_n714));
  XOR2_X1   g513(.A(KEYINPUT16), .B(G8gat), .Z(new_n715));
  AND3_X1   g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n552), .B1(new_n713), .B2(new_n714), .ZN(new_n717));
  OAI21_X1  g516(.A(KEYINPUT42), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n718), .B1(KEYINPUT42), .B2(new_n716), .ZN(G1325gat));
  INV_X1    g518(.A(new_n709), .ZN(new_n720));
  OAI21_X1  g519(.A(G15gat), .B1(new_n720), .B2(new_n530), .ZN(new_n721));
  INV_X1    g520(.A(new_n529), .ZN(new_n722));
  NOR3_X1   g521(.A1(new_n708), .A2(G15gat), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n713), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n721), .A2(new_n724), .ZN(G1326gat));
  NAND2_X1  g524(.A1(new_n709), .A2(new_n495), .ZN(new_n726));
  XNOR2_X1  g525(.A(KEYINPUT43), .B(G22gat), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n726), .B(new_n727), .ZN(G1327gat));
  NAND2_X1  g527(.A1(new_n549), .A2(new_n550), .ZN(new_n729));
  INV_X1    g528(.A(new_n535), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n621), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n648), .A2(new_n686), .A3(new_n706), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n532), .A2(G29gat), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT45), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT44), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n551), .B2(new_n686), .ZN(new_n738));
  AND3_X1   g537(.A1(new_n546), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n739));
  AOI21_X1  g538(.A(KEYINPUT94), .B1(new_n546), .B2(KEYINPUT35), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n739), .A2(new_n740), .A3(new_n539), .ZN(new_n741));
  OAI211_X1 g540(.A(KEYINPUT44), .B(new_n685), .C1(new_n741), .C2(new_n535), .ZN(new_n742));
  INV_X1    g541(.A(new_n648), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n618), .A2(new_n619), .ZN(new_n744));
  INV_X1    g543(.A(new_n706), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(new_n746), .B(KEYINPUT105), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n738), .A2(new_n742), .A3(new_n533), .A4(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(G29gat), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n736), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT106), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n736), .A2(KEYINPUT106), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(G1328gat));
  NAND2_X1  g553(.A1(new_n713), .A2(new_n733), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n755), .A2(G36gat), .A3(new_n536), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT46), .ZN(new_n757));
  AND2_X1   g556(.A1(new_n738), .A2(new_n742), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n454), .A3(new_n747), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(G36gat), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1329gat));
  INV_X1    g560(.A(new_n530), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n738), .A2(new_n742), .A3(new_n762), .A4(new_n747), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n763), .A2(G43gat), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n722), .A2(G43gat), .ZN(new_n765));
  AND4_X1   g564(.A1(new_n732), .A2(new_n731), .A3(new_n733), .A4(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT47), .B1(new_n768), .B2(KEYINPUT107), .ZN(new_n769));
  AOI21_X1  g568(.A(new_n766), .B1(new_n763), .B2(G43gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT47), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n770), .A2(new_n771), .A3(new_n772), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n769), .A2(new_n773), .ZN(G1330gat));
  NAND4_X1  g573(.A1(new_n738), .A2(new_n742), .A3(new_n495), .A4(new_n747), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(G50gat), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n496), .A2(G50gat), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n755), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(KEYINPUT48), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g579(.A(new_n776), .B(KEYINPUT48), .C1(new_n755), .C2(new_n777), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(G1331gat));
  INV_X1    g581(.A(new_n744), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n648), .A2(new_n783), .A3(new_n686), .A4(new_n706), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n551), .A2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n533), .ZN(new_n786));
  XOR2_X1   g585(.A(KEYINPUT108), .B(G57gat), .Z(new_n787));
  XNOR2_X1  g586(.A(new_n786), .B(new_n787), .ZN(G1332gat));
  AOI21_X1  g587(.A(new_n536), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n789));
  AND2_X1   g588(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g591(.A(KEYINPUT109), .B(KEYINPUT110), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n790), .A2(new_n791), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n792), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n792), .B2(new_n794), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(G1333gat));
  NAND3_X1  g596(.A1(new_n785), .A2(G71gat), .A3(new_n762), .ZN(new_n798));
  XOR2_X1   g597(.A(new_n529), .B(KEYINPUT111), .Z(new_n799));
  AND2_X1   g598(.A1(new_n785), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n798), .B1(new_n800), .B2(G71gat), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g601(.A1(new_n785), .A2(new_n495), .ZN(new_n803));
  XNOR2_X1  g602(.A(KEYINPUT112), .B(G78gat), .ZN(new_n804));
  XNOR2_X1  g603(.A(new_n803), .B(new_n804), .ZN(G1335gat));
  NOR3_X1   g604(.A1(new_n648), .A2(new_n744), .A3(new_n745), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n758), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G85gat), .B1(new_n807), .B2(new_n532), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n648), .A2(new_n744), .ZN(new_n809));
  OAI211_X1 g608(.A(new_n685), .B(new_n809), .C1(new_n741), .C2(new_n535), .ZN(new_n810));
  INV_X1    g609(.A(KEYINPUT51), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n731), .A2(KEYINPUT51), .A3(new_n685), .A4(new_n809), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  NAND4_X1  g613(.A1(new_n814), .A2(new_n649), .A3(new_n533), .A4(new_n706), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n808), .A2(new_n815), .ZN(G1336gat));
  NAND3_X1  g615(.A1(new_n812), .A2(KEYINPUT113), .A3(new_n813), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT113), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n810), .A2(new_n818), .A3(new_n811), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n536), .A2(G92gat), .A3(new_n745), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n738), .A2(new_n742), .A3(new_n454), .A4(new_n806), .ZN(new_n822));
  INV_X1    g621(.A(new_n665), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(new_n814), .B2(new_n820), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n824), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(G1337gat));
  OAI21_X1  g628(.A(G99gat), .B1(new_n807), .B2(new_n530), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n722), .A2(G99gat), .A3(new_n745), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1338gat));
  NOR3_X1   g632(.A1(new_n496), .A2(G106gat), .A3(new_n745), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n817), .A2(new_n819), .A3(new_n834), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n738), .A2(new_n742), .A3(new_n495), .A4(new_n806), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT53), .ZN(new_n839));
  AOI21_X1  g638(.A(KEYINPUT53), .B1(new_n814), .B2(new_n834), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n840), .A2(new_n837), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n839), .A2(new_n841), .ZN(G1339gat));
  NAND2_X1  g641(.A1(new_n744), .A2(new_n224), .ZN(new_n843));
  XOR2_X1   g642(.A(new_n843), .B(KEYINPUT116), .Z(new_n844));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n691), .A2(new_n692), .A3(new_n697), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n697), .B1(new_n691), .B2(new_n692), .ZN(new_n847));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n846), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n693), .A2(new_n848), .A3(new_n694), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n703), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n845), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n691), .A2(new_n692), .A3(new_n697), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n695), .A2(KEYINPUT54), .A3(new_n853), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n702), .B1(new_n847), .B2(new_n848), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n854), .A2(KEYINPUT55), .A3(new_n855), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n852), .A2(new_n705), .A3(new_n856), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n857), .A2(KEYINPUT114), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(KEYINPUT114), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n858), .A2(new_n744), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n603), .A2(new_n604), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n592), .B1(new_n591), .B2(new_n595), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n610), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n619), .A2(new_n863), .ZN(new_n864));
  INV_X1    g663(.A(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n706), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n685), .B1(new_n860), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n686), .A2(new_n864), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n868), .A2(new_n859), .A3(new_n858), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n743), .B1(new_n867), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n707), .A2(new_n783), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n532), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n542), .ZN(new_n873));
  INV_X1    g672(.A(new_n545), .ZN(new_n874));
  NOR3_X1   g673(.A1(new_n873), .A2(new_n454), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n876), .A2(KEYINPUT115), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n876), .A2(KEYINPUT115), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n844), .B1(new_n877), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n495), .B1(new_n870), .B2(new_n871), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n722), .A2(new_n532), .A3(new_n454), .ZN(new_n881));
  AND2_X1   g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(G113gat), .B1(new_n883), .B2(new_n621), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n879), .A2(new_n884), .ZN(G1340gat));
  NAND3_X1  g684(.A1(new_n706), .A2(new_n235), .A3(new_n237), .ZN(new_n886));
  XNOR2_X1  g685(.A(new_n886), .B(KEYINPUT117), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n887), .B1(new_n877), .B2(new_n878), .ZN(new_n888));
  OAI21_X1  g687(.A(G120gat), .B1(new_n883), .B2(new_n745), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n888), .A2(new_n889), .ZN(G1341gat));
  OAI211_X1 g689(.A(new_n882), .B(new_n648), .C1(new_n218), .C2(new_n219), .ZN(new_n891));
  OR2_X1    g690(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n213), .B1(new_n876), .B2(new_n743), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(KEYINPUT118), .ZN(new_n894));
  AND3_X1   g693(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(G1342gat));
  OAI21_X1  g694(.A(G134gat), .B1(new_n883), .B2(new_n686), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n686), .A2(G134gat), .ZN(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  OR3_X1    g697(.A1(new_n876), .A2(KEYINPUT56), .A3(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT56), .B1(new_n876), .B2(new_n898), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n896), .A2(new_n899), .A3(new_n900), .ZN(G1343gat));
  INV_X1    g700(.A(KEYINPUT58), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n762), .A2(new_n532), .A3(new_n454), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n870), .A2(new_n871), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT57), .B1(new_n904), .B2(new_n495), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n495), .A2(KEYINPUT57), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT119), .ZN(new_n907));
  NAND4_X1  g706(.A1(new_n852), .A2(new_n907), .A3(new_n705), .A4(new_n856), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n856), .A2(new_n705), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT55), .B1(new_n854), .B2(new_n855), .ZN(new_n910));
  OAI21_X1  g709(.A(KEYINPUT119), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n908), .B(new_n911), .C1(new_n617), .C2(new_n620), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n685), .B1(new_n912), .B2(new_n866), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n743), .B1(new_n913), .B2(new_n869), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n906), .B1(new_n914), .B2(new_n871), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n903), .B1(new_n905), .B2(new_n915), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n916), .A2(new_n783), .ZN(new_n917));
  AND4_X1   g716(.A1(new_n530), .A2(new_n872), .A3(new_n536), .A4(new_n495), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n621), .A2(G141gat), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n917), .A2(G141gat), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g719(.A(G141gat), .B1(new_n916), .B2(new_n621), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT120), .ZN(new_n922));
  AOI21_X1  g721(.A(KEYINPUT58), .B1(new_n918), .B2(new_n919), .ZN(new_n923));
  AND3_X1   g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n921), .B2(new_n923), .ZN(new_n925));
  OAI22_X1  g724(.A1(new_n902), .A2(new_n920), .B1(new_n924), .B2(new_n925), .ZN(G1344gat));
  INV_X1    g725(.A(KEYINPUT59), .ZN(new_n927));
  OAI211_X1 g726(.A(new_n927), .B(G148gat), .C1(new_n916), .C2(new_n745), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n904), .A2(KEYINPUT57), .A3(new_n495), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n686), .A2(new_n864), .A3(new_n857), .ZN(new_n932));
  INV_X1    g731(.A(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n616), .B1(new_n613), .B2(new_n615), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n618), .A2(KEYINPUT98), .A3(new_n619), .ZN(new_n935));
  AOI22_X1  g734(.A1(new_n934), .A2(new_n935), .B1(new_n857), .B2(KEYINPUT119), .ZN(new_n936));
  AOI22_X1  g735(.A1(new_n936), .A2(new_n908), .B1(new_n706), .B2(new_n865), .ZN(new_n937));
  OAI211_X1 g736(.A(new_n931), .B(new_n933), .C1(new_n937), .C2(new_n685), .ZN(new_n938));
  OAI21_X1  g737(.A(KEYINPUT121), .B1(new_n913), .B2(new_n932), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n743), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n707), .A2(new_n621), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n496), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n930), .B1(new_n942), .B2(KEYINPUT57), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n903), .A2(new_n706), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n945), .A2(G148gat), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n929), .B1(new_n946), .B2(KEYINPUT59), .ZN(new_n947));
  INV_X1    g746(.A(G148gat), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n948), .B1(new_n943), .B2(new_n944), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n949), .A2(KEYINPUT122), .A3(new_n927), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n928), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n918), .A2(new_n948), .A3(new_n706), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(new_n952), .ZN(G1345gat));
  OAI21_X1  g752(.A(G155gat), .B1(new_n916), .B2(new_n743), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n918), .A2(new_n246), .A3(new_n648), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1346gat));
  OR2_X1    g755(.A1(new_n916), .A2(new_n686), .ZN(new_n957));
  INV_X1    g756(.A(KEYINPUT123), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n247), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n959), .B1(new_n958), .B2(new_n957), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n918), .A2(new_n247), .A3(new_n685), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(G1347gat));
  NOR2_X1   g761(.A1(new_n536), .A2(new_n533), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n880), .A2(new_n799), .A3(new_n963), .ZN(new_n964));
  OAI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n621), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n533), .B1(new_n870), .B2(new_n871), .ZN(new_n966));
  NAND4_X1  g765(.A1(new_n966), .A2(new_n454), .A3(new_n542), .A4(new_n545), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n744), .A2(new_n399), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n965), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(KEYINPUT124), .ZN(G1348gat));
  OAI21_X1  g769(.A(G176gat), .B1(new_n964), .B2(new_n745), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n706), .A2(new_n365), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n967), .B2(new_n972), .ZN(G1349gat));
  OAI21_X1  g772(.A(G183gat), .B1(new_n964), .B2(new_n743), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n648), .A2(new_n382), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n974), .B1(new_n967), .B2(new_n975), .ZN(new_n976));
  XNOR2_X1  g775(.A(new_n976), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g776(.A(G190gat), .B1(new_n964), .B2(new_n686), .ZN(new_n978));
  AND2_X1   g777(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n979));
  NOR2_X1   g778(.A1(new_n978), .A2(KEYINPUT61), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n685), .A2(new_n381), .ZN(new_n981));
  OAI22_X1  g780(.A1(new_n979), .A2(new_n980), .B1(new_n967), .B2(new_n981), .ZN(G1351gat));
  AND4_X1   g781(.A1(new_n530), .A2(new_n966), .A3(new_n454), .A4(new_n495), .ZN(new_n983));
  AOI21_X1  g782(.A(G197gat), .B1(new_n983), .B2(new_n744), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n530), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT125), .ZN(new_n986));
  INV_X1    g785(.A(new_n986), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n943), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n621), .A2(new_n335), .ZN(new_n989));
  AOI21_X1  g788(.A(new_n984), .B1(new_n988), .B2(new_n989), .ZN(G1352gat));
  NAND3_X1  g789(.A1(new_n983), .A2(new_n336), .A3(new_n706), .ZN(new_n991));
  XOR2_X1   g790(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n992));
  XNOR2_X1  g791(.A(new_n991), .B(new_n992), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n988), .A2(new_n706), .ZN(new_n994));
  OAI21_X1  g793(.A(new_n993), .B1(new_n336), .B2(new_n994), .ZN(G1353gat));
  NAND3_X1  g794(.A1(new_n983), .A2(new_n342), .A3(new_n648), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n988), .A2(new_n648), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n996), .B1(new_n998), .B2(new_n999), .ZN(G1354gat));
  NAND3_X1  g799(.A1(new_n983), .A2(new_n343), .A3(new_n685), .ZN(new_n1001));
  AND2_X1   g800(.A1(new_n988), .A2(new_n685), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1001), .B1(new_n1002), .B2(new_n343), .ZN(G1355gat));
endmodule


