//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 1 1 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1326, new_n1327, new_n1328, new_n1329,
    new_n1330, new_n1331, new_n1332, new_n1333, new_n1334, new_n1335,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g0017(.A(KEYINPUT65), .B(G244), .Z(new_n218));
  XNOR2_X1  g0018(.A(KEYINPUT64), .B(G77), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G107), .A2(G264), .ZN(new_n224));
  NAND4_X1  g0024(.A1(new_n221), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n209), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT2), .B(G226), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XNOR2_X1  g0036(.A(G50), .B(G68), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G58), .B(G77), .ZN(new_n238));
  XOR2_X1   g0038(.A(new_n237), .B(new_n238), .Z(new_n239));
  XOR2_X1   g0039(.A(G87), .B(G97), .Z(new_n240));
  XNOR2_X1  g0040(.A(G107), .B(G116), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G351));
  NAND3_X1  g0043(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n244));
  AND2_X1   g0044(.A1(new_n244), .A2(new_n215), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n206), .A2(G20), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G50), .ZN(new_n249));
  OAI22_X1  g0049(.A1(new_n247), .A2(new_n249), .B1(G50), .B2(new_n246), .ZN(new_n250));
  XNOR2_X1  g0050(.A(KEYINPUT8), .B(G58), .ZN(new_n251));
  INV_X1    g0051(.A(new_n251), .ZN(new_n252));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(new_n253), .A2(G20), .ZN(new_n254));
  NOR2_X1   g0054(.A1(G20), .A2(G33), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n252), .A2(new_n254), .B1(G150), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n203), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n244), .A2(new_n215), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n250), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  XOR2_X1   g0060(.A(new_n260), .B(KEYINPUT9), .Z(new_n261));
  AND2_X1   g0061(.A1(KEYINPUT66), .A2(G41), .ZN(new_n262));
  NOR2_X1   g0062(.A1(KEYINPUT66), .A2(G41), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G45), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G274), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G1), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G41), .ZN(new_n271));
  OAI211_X1 g0071(.A(G1), .B(G13), .C1(new_n253), .C2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AOI21_X1  g0074(.A(new_n270), .B1(G226), .B2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n272), .B1(new_n279), .B2(new_n219), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G222), .A2(G1698), .ZN(new_n281));
  XOR2_X1   g0081(.A(KEYINPUT67), .B(G223), .Z(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G1698), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(new_n279), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n275), .A2(new_n284), .ZN(new_n285));
  XOR2_X1   g0085(.A(KEYINPUT68), .B(G200), .Z(new_n286));
  INV_X1    g0086(.A(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G190), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n261), .B(new_n288), .C1(new_n289), .C2(new_n285), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT10), .ZN(new_n291));
  INV_X1    g0091(.A(G169), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n260), .B1(new_n285), .B2(new_n292), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n293), .B1(G179), .B2(new_n285), .ZN(new_n294));
  AND2_X1   g0094(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(KEYINPUT16), .ZN(new_n296));
  INV_X1    g0096(.A(G58), .ZN(new_n297));
  INV_X1    g0097(.A(G68), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n299), .A2(new_n201), .ZN(new_n300));
  AOI22_X1  g0100(.A1(new_n300), .A2(G20), .B1(G159), .B2(new_n255), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  XOR2_X1   g0102(.A(KEYINPUT72), .B(KEYINPUT7), .Z(new_n303));
  XNOR2_X1  g0103(.A(KEYINPUT3), .B(G33), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(G20), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT7), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n306), .A2(KEYINPUT72), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n279), .A2(new_n207), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n298), .B1(new_n305), .B2(new_n308), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n296), .B1(new_n302), .B2(new_n309), .ZN(new_n310));
  NOR3_X1   g0110(.A1(new_n253), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n311), .B1(new_n304), .B2(KEYINPUT71), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n312), .A2(new_n306), .A3(new_n207), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(G68), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n306), .B1(new_n312), .B2(new_n207), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n301), .B1(new_n314), .B2(new_n315), .ZN(new_n316));
  OAI211_X1 g0116(.A(new_n310), .B(new_n259), .C1(new_n316), .C2(new_n296), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n252), .A2(new_n248), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n318), .A2(new_n247), .B1(new_n246), .B2(new_n252), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI22_X1  g0120(.A1(new_n274), .A2(G232), .B1(new_n266), .B2(new_n268), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n277), .A2(new_n278), .A3(KEYINPUT71), .ZN(new_n322));
  OR3_X1    g0122(.A1(new_n253), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  MUX2_X1   g0124(.A(G223), .B(G226), .S(G1698), .Z(new_n325));
  AOI22_X1  g0125(.A1(new_n324), .A2(new_n325), .B1(G33), .B2(G87), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n321), .B1(new_n326), .B2(new_n272), .ZN(new_n327));
  OR2_X1    g0127(.A1(new_n327), .A2(new_n289), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(G200), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n317), .A2(new_n320), .A3(new_n328), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT17), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n317), .A2(new_n320), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n327), .A2(G169), .ZN(new_n334));
  INV_X1    g0134(.A(G179), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n334), .B1(new_n335), .B2(new_n327), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(KEYINPUT18), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT18), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n333), .A2(new_n339), .A3(new_n336), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n330), .A2(new_n331), .ZN(new_n341));
  NAND4_X1  g0141(.A1(new_n332), .A2(new_n338), .A3(new_n340), .A4(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n246), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n298), .ZN(new_n345));
  XNOR2_X1  g0145(.A(new_n345), .B(KEYINPUT12), .ZN(new_n346));
  AOI22_X1  g0146(.A1(new_n255), .A2(G50), .B1(G20), .B2(new_n298), .ZN(new_n347));
  INV_X1    g0147(.A(new_n254), .ZN(new_n348));
  INV_X1    g0148(.A(G77), .ZN(new_n349));
  OAI21_X1  g0149(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n350), .A2(KEYINPUT11), .A3(new_n259), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n248), .A2(G68), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n346), .B(new_n351), .C1(new_n247), .C2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT11), .B1(new_n350), .B2(new_n259), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT13), .ZN(new_n357));
  INV_X1    g0157(.A(G1698), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n358), .A2(G232), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n304), .B(new_n359), .C1(G226), .C2(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(G33), .A2(G97), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  INV_X1    g0162(.A(new_n272), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n272), .A2(G238), .A3(new_n273), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n269), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n357), .B1(new_n364), .B2(new_n366), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n272), .B1(new_n360), .B2(new_n361), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n269), .A2(new_n365), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n368), .A2(new_n369), .A3(KEYINPUT13), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n367), .A2(new_n370), .A3(new_n289), .ZN(new_n371));
  INV_X1    g0171(.A(G200), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n364), .A2(new_n366), .A3(new_n357), .ZN(new_n373));
  OAI21_X1  g0173(.A(KEYINPUT13), .B1(new_n368), .B2(new_n369), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR3_X1   g0175(.A1(new_n356), .A2(new_n371), .A3(new_n375), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n373), .A2(new_n374), .A3(G179), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT70), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n377), .B(new_n378), .ZN(new_n379));
  OAI21_X1  g0179(.A(G169), .B1(new_n367), .B2(new_n370), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n380), .A2(KEYINPUT14), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g0183(.A(new_n376), .B1(new_n383), .B2(new_n356), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n248), .A2(G77), .ZN(new_n385));
  INV_X1    g0185(.A(new_n219), .ZN(new_n386));
  OAI22_X1  g0186(.A1(new_n247), .A2(new_n385), .B1(new_n386), .B2(new_n246), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT15), .B(G87), .ZN(new_n388));
  INV_X1    g0188(.A(new_n388), .ZN(new_n389));
  AOI22_X1  g0189(.A1(new_n386), .A2(G20), .B1(new_n389), .B2(new_n254), .ZN(new_n390));
  INV_X1    g0190(.A(new_n255), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n390), .B1(new_n391), .B2(new_n251), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n387), .B1(new_n392), .B2(new_n259), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G232), .A2(G1698), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n358), .A2(G238), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n304), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  OAI211_X1 g0196(.A(new_n396), .B(new_n363), .C1(G107), .C2(new_n304), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n272), .A2(new_n273), .ZN(new_n398));
  OAI211_X1 g0198(.A(new_n397), .B(new_n269), .C1(new_n218), .C2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n393), .B1(new_n292), .B2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n400), .B1(G179), .B2(new_n399), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n399), .A2(new_n287), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n402), .B(new_n393), .C1(new_n289), .C2(new_n399), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  XOR2_X1   g0204(.A(new_n404), .B(KEYINPUT69), .Z(new_n405));
  NAND4_X1  g0205(.A1(new_n295), .A2(new_n343), .A3(new_n384), .A4(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT6), .ZN(new_n408));
  INV_X1    g0208(.A(G97), .ZN(new_n409));
  NOR3_X1   g0209(.A1(new_n408), .A2(new_n409), .A3(G107), .ZN(new_n410));
  XNOR2_X1  g0210(.A(G97), .B(G107), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n410), .B1(new_n408), .B2(new_n411), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n412), .A2(new_n207), .B1(new_n349), .B2(new_n391), .ZN(new_n413));
  INV_X1    g0213(.A(G107), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(new_n305), .B2(new_n308), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n259), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n206), .A2(G33), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n246), .A2(new_n417), .A3(new_n215), .A4(new_n244), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G97), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n246), .A2(new_n409), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT73), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(KEYINPUT73), .A3(new_n420), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT5), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n427), .B1(new_n262), .B2(new_n263), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n271), .A2(KEYINPUT5), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n206), .A2(G45), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n428), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(G257), .A3(new_n272), .ZN(new_n433));
  NOR2_X1   g0233(.A1(new_n430), .A2(new_n267), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n428), .A2(new_n434), .A3(new_n272), .A4(new_n429), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n358), .A2(KEYINPUT4), .A3(G244), .ZN(new_n437));
  INV_X1    g0237(.A(G250), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n437), .B1(new_n438), .B2(new_n358), .ZN(new_n439));
  AOI22_X1  g0239(.A1(new_n439), .A2(new_n304), .B1(G33), .B2(G283), .ZN(new_n440));
  INV_X1    g0240(.A(G244), .ZN(new_n441));
  AOI211_X1 g0241(.A(new_n441), .B(G1698), .C1(new_n322), .C2(new_n323), .ZN(new_n442));
  XOR2_X1   g0242(.A(KEYINPUT74), .B(KEYINPUT4), .Z(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n440), .B1(new_n442), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n436), .B1(new_n445), .B2(new_n363), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n426), .B1(new_n446), .B2(G169), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n436), .A2(KEYINPUT75), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n441), .B1(new_n322), .B2(new_n323), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n444), .B1(new_n449), .B2(new_n358), .ZN(new_n450));
  INV_X1    g0250(.A(new_n440), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n363), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT75), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n433), .A2(new_n453), .A3(new_n435), .ZN(new_n454));
  AND4_X1   g0254(.A1(new_n335), .A2(new_n448), .A3(new_n452), .A4(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT77), .B1(new_n447), .B2(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n436), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  AOI22_X1  g0258(.A1(new_n458), .A2(new_n292), .B1(new_n416), .B2(new_n425), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n448), .A2(new_n452), .A3(new_n335), .A4(new_n454), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n448), .A2(new_n452), .A3(new_n454), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n464), .A2(KEYINPUT76), .A3(G200), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT76), .B1(new_n464), .B2(G200), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n416), .B(new_n425), .C1(new_n458), .C2(new_n289), .ZN(new_n467));
  NOR3_X1   g0267(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n463), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT80), .ZN(new_n470));
  AOI21_X1  g0270(.A(G20), .B1(new_n322), .B2(new_n323), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G68), .ZN(new_n472));
  NOR3_X1   g0272(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n473));
  AOI21_X1  g0273(.A(G20), .B1(G33), .B2(G97), .ZN(new_n474));
  OAI21_X1  g0274(.A(KEYINPUT19), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT19), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n254), .A2(new_n476), .A3(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n245), .B1(new_n472), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n389), .A2(new_n246), .ZN(new_n480));
  INV_X1    g0280(.A(G87), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n418), .A2(new_n481), .ZN(new_n482));
  NOR3_X1   g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n358), .A2(G238), .ZN(new_n484));
  INV_X1    g0284(.A(G116), .ZN(new_n485));
  OAI22_X1  g0285(.A1(new_n312), .A2(new_n484), .B1(new_n253), .B2(new_n485), .ZN(new_n486));
  AOI211_X1 g0286(.A(new_n441), .B(new_n358), .C1(new_n322), .C2(new_n323), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n363), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n434), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n430), .A2(G250), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n363), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g0291(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n488), .A2(G190), .A3(new_n492), .ZN(new_n493));
  NOR2_X1   g0293(.A1(new_n253), .A2(new_n485), .ZN(new_n494));
  INV_X1    g0294(.A(new_n484), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n494), .B1(new_n324), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n324), .A2(G244), .A3(G1698), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n272), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  OAI21_X1  g0298(.A(new_n287), .B1(new_n498), .B2(new_n491), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n483), .A2(new_n493), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n488), .A2(new_n335), .A3(new_n492), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT78), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n496), .A2(new_n497), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n491), .B1(new_n503), .B2(new_n363), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT78), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n504), .A2(new_n505), .A3(new_n335), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n488), .A2(new_n492), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n292), .ZN(new_n508));
  XNOR2_X1  g0308(.A(new_n388), .B(KEYINPUT79), .ZN(new_n509));
  INV_X1    g0309(.A(new_n418), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(new_n480), .ZN(new_n512));
  AOI22_X1  g0312(.A1(new_n471), .A2(G68), .B1(new_n475), .B2(new_n477), .ZN(new_n513));
  OAI211_X1 g0313(.A(new_n511), .B(new_n512), .C1(new_n513), .C2(new_n245), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n502), .A2(new_n506), .A3(new_n508), .A4(new_n514), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n469), .A2(new_n470), .A3(new_n500), .A4(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n464), .A2(G200), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT76), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n464), .A2(KEYINPUT76), .A3(G200), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n426), .B1(G190), .B2(new_n446), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(new_n456), .A3(new_n462), .A4(new_n500), .ZN(new_n523));
  INV_X1    g0323(.A(new_n515), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT80), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NOR4_X1   g0325(.A1(new_n279), .A2(KEYINPUT22), .A3(G20), .A4(new_n481), .ZN(new_n526));
  AOI211_X1 g0326(.A(G20), .B(new_n481), .C1(new_n322), .C2(new_n323), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT22), .ZN(new_n528));
  OAI21_X1  g0328(.A(KEYINPUT81), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n324), .A2(new_n207), .A3(G87), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT81), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n530), .A2(new_n531), .A3(KEYINPUT22), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n526), .B1(new_n529), .B2(new_n532), .ZN(new_n533));
  AOI21_X1  g0333(.A(KEYINPUT23), .B1(new_n414), .B2(G20), .ZN(new_n534));
  INV_X1    g0334(.A(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n414), .A2(KEYINPUT23), .A3(G20), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n535), .A2(new_n536), .B1(new_n494), .B2(new_n207), .ZN(new_n537));
  INV_X1    g0337(.A(new_n537), .ZN(new_n538));
  NOR3_X1   g0338(.A1(new_n533), .A2(KEYINPUT24), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT24), .ZN(new_n540));
  INV_X1    g0340(.A(new_n526), .ZN(new_n541));
  AOI211_X1 g0341(.A(KEYINPUT81), .B(new_n528), .C1(new_n471), .C2(G87), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n531), .B1(new_n530), .B2(KEYINPUT22), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n540), .B1(new_n544), .B2(new_n537), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n259), .B1(new_n539), .B2(new_n545), .ZN(new_n546));
  AOI21_X1  g0346(.A(KEYINPUT25), .B1(new_n344), .B2(new_n414), .ZN(new_n547));
  INV_X1    g0347(.A(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n344), .A2(KEYINPUT25), .A3(new_n414), .ZN(new_n549));
  AOI22_X1  g0349(.A1(new_n548), .A2(new_n549), .B1(G107), .B2(new_n510), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n432), .A2(G264), .A3(new_n272), .ZN(new_n551));
  NOR2_X1   g0351(.A1(G250), .A2(G1698), .ZN(new_n552));
  INV_X1    g0352(.A(G257), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G1698), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n324), .A2(new_n554), .B1(G33), .B2(G294), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n435), .B(new_n551), .C1(new_n555), .C2(new_n272), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n556), .A2(G190), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n372), .B2(new_n556), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n546), .A2(new_n550), .A3(new_n559), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n556), .A2(G179), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n561), .B1(new_n292), .B2(new_n556), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT24), .B1(new_n533), .B2(new_n538), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n544), .A2(new_n540), .A3(new_n537), .ZN(new_n564));
  AOI21_X1  g0364(.A(new_n245), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n550), .ZN(new_n566));
  OAI21_X1  g0366(.A(new_n562), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT21), .ZN(new_n568));
  NAND2_X1  g0368(.A1(G33), .A2(G283), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n569), .B(new_n207), .C1(G33), .C2(new_n409), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n570), .B(new_n259), .C1(new_n207), .C2(G116), .ZN(new_n571));
  XNOR2_X1  g0371(.A(new_n571), .B(KEYINPUT20), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n344), .A2(new_n485), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n573), .B1(new_n418), .B2(new_n485), .ZN(new_n574));
  OAI21_X1  g0374(.A(G169), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n553), .A2(new_n358), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n576), .B1(G264), .B2(new_n358), .ZN(new_n577));
  AOI21_X1  g0377(.A(new_n577), .B1(new_n323), .B2(new_n322), .ZN(new_n578));
  INV_X1    g0378(.A(G303), .ZN(new_n579));
  NOR2_X1   g0379(.A1(new_n304), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n363), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n432), .A2(G270), .A3(new_n272), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n581), .A2(new_n435), .A3(new_n582), .ZN(new_n583));
  INV_X1    g0383(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n568), .B1(new_n575), .B2(new_n584), .ZN(new_n585));
  INV_X1    g0385(.A(new_n575), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n586), .A2(KEYINPUT21), .A3(new_n583), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n583), .A2(G200), .ZN(new_n588));
  NOR2_X1   g0388(.A1(new_n572), .A2(new_n574), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n588), .B(new_n589), .C1(new_n289), .C2(new_n583), .ZN(new_n590));
  NOR2_X1   g0390(.A1(new_n583), .A2(new_n335), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n591), .B1(new_n572), .B2(new_n574), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n585), .A2(new_n587), .A3(new_n590), .A4(new_n592), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n560), .A2(new_n567), .A3(new_n593), .ZN(new_n594));
  AND4_X1   g0394(.A1(new_n407), .A2(new_n516), .A3(new_n525), .A4(new_n594), .ZN(G372));
  NAND2_X1  g0395(.A1(new_n383), .A2(new_n356), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n596), .B1(new_n376), .B2(new_n401), .ZN(new_n597));
  XNOR2_X1  g0397(.A(new_n330), .B(KEYINPUT17), .ZN(new_n598));
  AND2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n333), .A2(new_n339), .A3(new_n336), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n339), .B1(new_n333), .B2(new_n336), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n291), .B1(new_n599), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n294), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n483), .A2(new_n493), .A3(new_n499), .ZN(new_n607));
  OAI21_X1  g0407(.A(new_n514), .B1(new_n504), .B2(G169), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n505), .B1(new_n504), .B2(new_n335), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n607), .B1(new_n610), .B2(new_n506), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n463), .A2(new_n611), .A3(KEYINPUT26), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT26), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n508), .A2(new_n501), .A3(new_n514), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(new_n500), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n459), .A2(new_n461), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n613), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n612), .A2(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n324), .A2(G244), .A3(new_n358), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(new_n443), .ZN(new_n621));
  AOI21_X1  g0421(.A(new_n272), .B1(new_n621), .B2(new_n440), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n292), .B1(new_n622), .B2(new_n436), .ZN(new_n623));
  AND4_X1   g0423(.A1(new_n460), .A2(new_n623), .A3(new_n461), .A4(new_n426), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n560), .A2(new_n625), .A3(new_n522), .A4(new_n500), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n587), .A2(new_n585), .A3(new_n592), .ZN(new_n627));
  AND2_X1   g0427(.A1(new_n567), .A2(new_n627), .ZN(new_n628));
  OAI211_X1 g0428(.A(new_n618), .B(new_n614), .C1(new_n626), .C2(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(new_n629), .ZN(new_n630));
  OAI21_X1  g0430(.A(new_n606), .B1(new_n406), .B2(new_n630), .ZN(G369));
  NAND3_X1  g0431(.A1(new_n206), .A2(new_n207), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(new_n634), .A3(G213), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n637), .B1(new_n565), .B2(new_n566), .ZN(new_n638));
  NAND3_X1  g0438(.A1(new_n560), .A2(new_n567), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT82), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT82), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n560), .A2(new_n567), .A3(new_n638), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n640), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n562), .B(new_n637), .C1(new_n565), .C2(new_n566), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n637), .B1(new_n572), .B2(new_n574), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n593), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n627), .B2(new_n647), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n649), .A2(G330), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n646), .A2(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n627), .A2(new_n637), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n640), .A2(new_n642), .A3(new_n652), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n567), .A2(new_n637), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  OR2_X1    g0455(.A1(new_n651), .A2(new_n655), .ZN(G399));
  NAND2_X1  g0456(.A1(new_n210), .A2(new_n264), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n473), .A2(new_n485), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n658), .A2(new_n206), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n214), .B2(new_n658), .ZN(new_n661));
  XOR2_X1   g0461(.A(new_n661), .B(KEYINPUT28), .Z(new_n662));
  INV_X1    g0462(.A(KEYINPUT29), .ZN(new_n663));
  INV_X1    g0463(.A(new_n637), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n629), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n614), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n565), .A2(new_n558), .A3(new_n566), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n523), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n567), .A2(new_n627), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n666), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n614), .A2(new_n500), .ZN(new_n671));
  INV_X1    g0471(.A(new_n616), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n613), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n515), .A2(new_n500), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n674), .B1(new_n456), .B2(new_n462), .ZN(new_n675));
  AOI21_X1  g0475(.A(new_n673), .B1(new_n675), .B2(new_n613), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n637), .B1(new_n670), .B2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n665), .B1(new_n677), .B2(new_n663), .ZN(new_n678));
  INV_X1    g0478(.A(G330), .ZN(new_n679));
  NAND4_X1  g0479(.A1(new_n516), .A2(new_n525), .A3(new_n594), .A4(new_n664), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n555), .A2(new_n272), .ZN(new_n681));
  INV_X1    g0481(.A(new_n551), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND4_X1  g0483(.A1(new_n591), .A2(new_n446), .A3(new_n504), .A4(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(KEYINPUT30), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g0486(.A1(new_n584), .A2(new_n504), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n687), .A2(new_n335), .A3(new_n464), .A4(new_n556), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(KEYINPUT83), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n690), .B1(new_n684), .B2(new_n685), .ZN(new_n691));
  AND3_X1   g0491(.A1(new_n591), .A2(new_n504), .A3(new_n683), .ZN(new_n692));
  NAND4_X1  g0492(.A1(new_n692), .A2(KEYINPUT83), .A3(KEYINPUT30), .A4(new_n446), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n689), .B1(new_n691), .B2(new_n693), .ZN(new_n694));
  OAI21_X1  g0494(.A(KEYINPUT31), .B1(new_n694), .B2(new_n664), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT31), .ZN(new_n696));
  AND2_X1   g0496(.A1(new_n693), .A2(new_n691), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n696), .B(new_n637), .C1(new_n697), .C2(new_n689), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n695), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n679), .B1(new_n680), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g0500(.A(KEYINPUT84), .B1(new_n678), .B2(new_n700), .ZN(new_n701));
  OAI211_X1 g0501(.A(new_n676), .B(new_n614), .C1(new_n628), .C2(new_n626), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n663), .B1(new_n702), .B2(new_n664), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n680), .A2(new_n699), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n705), .A2(G330), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT84), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n704), .A2(new_n706), .A3(new_n707), .A4(new_n665), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n701), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n662), .B1(new_n709), .B2(G1), .ZN(G364));
  NOR2_X1   g0510(.A1(new_n649), .A2(G330), .ZN(new_n711));
  XOR2_X1   g0511(.A(new_n711), .B(KEYINPUT85), .Z(new_n712));
  INV_X1    g0512(.A(G13), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(G20), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n206), .B1(new_n714), .B2(G45), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n658), .A2(new_n716), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n650), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n210), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n720), .A2(new_n279), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G355), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n722), .B1(G116), .B2(new_n210), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n720), .A2(new_n324), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n265), .B2(new_n214), .ZN(new_n726));
  OR2_X1    g0526(.A1(new_n239), .A2(new_n265), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n723), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(G13), .A2(G33), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT86), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n730), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n215), .B1(G20), .B2(new_n292), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n717), .B1(new_n728), .B2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G179), .A2(G200), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n736), .A2(G190), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G294), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n736), .A2(G20), .A3(new_n289), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  AOI211_X1 g0543(.A(new_n304), .B(new_n741), .C1(G329), .C2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G283), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n207), .A2(G179), .ZN(new_n746));
  NAND3_X1  g0546(.A1(new_n287), .A2(new_n289), .A3(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n287), .A2(G190), .A3(new_n746), .ZN(new_n748));
  OAI221_X1 g0548(.A(new_n744), .B1(new_n745), .B2(new_n747), .C1(new_n579), .C2(new_n748), .ZN(new_n749));
  NAND2_X1  g0549(.A1(G20), .A2(G179), .ZN(new_n750));
  AOI21_X1  g0550(.A(G200), .B1(new_n750), .B2(KEYINPUT87), .ZN(new_n751));
  OAI21_X1  g0551(.A(new_n751), .B1(KEYINPUT87), .B2(new_n750), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n752), .A2(new_n289), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G311), .A2(new_n753), .B1(new_n754), .B2(G322), .ZN(new_n755));
  NAND3_X1  g0555(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n756));
  OR2_X1    g0556(.A1(new_n756), .A2(KEYINPUT88), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(KEYINPUT88), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n757), .A2(G190), .A3(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n760), .A2(G326), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n757), .A2(new_n289), .A3(new_n758), .ZN(new_n762));
  XOR2_X1   g0562(.A(KEYINPUT33), .B(G317), .Z(new_n763));
  OAI211_X1 g0563(.A(new_n755), .B(new_n761), .C1(new_n762), .C2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n747), .A2(new_n414), .ZN(new_n765));
  XNOR2_X1  g0565(.A(KEYINPUT89), .B(G159), .ZN(new_n766));
  INV_X1    g0566(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(new_n743), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT32), .ZN(new_n769));
  OAI21_X1  g0569(.A(new_n304), .B1(new_n739), .B2(new_n409), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n748), .A2(new_n481), .ZN(new_n771));
  OR4_X1    g0571(.A1(new_n765), .A2(new_n769), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  AOI22_X1  g0572(.A1(G50), .A2(new_n760), .B1(new_n754), .B2(G58), .ZN(new_n773));
  INV_X1    g0573(.A(new_n753), .ZN(new_n774));
  OAI221_X1 g0574(.A(new_n773), .B1(new_n298), .B2(new_n762), .C1(new_n219), .C2(new_n774), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n749), .A2(new_n764), .B1(new_n772), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n735), .B1(new_n776), .B2(new_n732), .ZN(new_n777));
  INV_X1    g0577(.A(new_n731), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n649), .B2(new_n778), .ZN(new_n779));
  AND2_X1   g0579(.A1(new_n719), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(G396));
  INV_X1    g0581(.A(G311), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n279), .B1(new_n742), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n747), .A2(new_n481), .ZN(new_n784));
  AOI211_X1 g0584(.A(new_n783), .B(new_n784), .C1(G97), .C2(new_n738), .ZN(new_n785));
  INV_X1    g0585(.A(new_n748), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n786), .A2(G107), .ZN(new_n787));
  INV_X1    g0587(.A(new_n762), .ZN(new_n788));
  AOI22_X1  g0588(.A1(G283), .A2(new_n788), .B1(new_n754), .B2(G294), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G303), .A2(new_n760), .B1(new_n753), .B2(G116), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n785), .A2(new_n787), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G137), .A2(new_n760), .B1(new_n788), .B2(G150), .ZN(new_n792));
  INV_X1    g0592(.A(new_n754), .ZN(new_n793));
  XOR2_X1   g0593(.A(KEYINPUT92), .B(G143), .Z(new_n794));
  OAI221_X1 g0594(.A(new_n792), .B1(new_n774), .B2(new_n766), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT34), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n797), .A2(KEYINPUT93), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n747), .A2(new_n298), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n312), .B1(G132), .B2(new_n743), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n800), .B1(new_n297), .B2(new_n739), .ZN(new_n801));
  AOI211_X1 g0601(.A(new_n799), .B(new_n801), .C1(G50), .C2(new_n786), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n797), .B2(KEYINPUT93), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n791), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n732), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n401), .A2(new_n637), .ZN(new_n806));
  OAI21_X1  g0606(.A(new_n403), .B1(new_n393), .B2(new_n664), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n401), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n730), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n732), .ZN(new_n812));
  INV_X1    g0612(.A(new_n729), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  XOR2_X1   g0614(.A(new_n814), .B(KEYINPUT90), .Z(new_n815));
  OAI21_X1  g0615(.A(new_n717), .B1(new_n815), .B2(G77), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT91), .Z(new_n817));
  NAND3_X1  g0617(.A1(new_n805), .A2(new_n811), .A3(new_n817), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n629), .A2(new_n664), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n809), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n404), .A2(new_n637), .ZN(new_n822));
  AND3_X1   g0622(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(KEYINPUT94), .B1(new_n629), .B2(new_n822), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n821), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AND3_X1   g0625(.A1(new_n825), .A2(KEYINPUT95), .A3(new_n706), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n718), .B1(new_n825), .B2(new_n706), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n629), .A2(new_n822), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT94), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n629), .A2(KEYINPUT94), .A3(new_n822), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n700), .B1(new_n833), .B2(new_n821), .ZN(new_n834));
  OR2_X1    g0634(.A1(new_n834), .A2(KEYINPUT95), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n819), .B1(new_n828), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(G384));
  NOR2_X1   g0637(.A1(new_n714), .A2(new_n206), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT37), .ZN(new_n839));
  INV_X1    g0639(.A(new_n635), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n333), .A2(new_n840), .ZN(new_n841));
  AND4_X1   g0641(.A1(new_n839), .A2(new_n337), .A3(new_n841), .A4(new_n330), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n259), .B1(new_n316), .B2(new_n296), .ZN(new_n843));
  OR2_X1    g0643(.A1(new_n316), .A2(KEYINPUT98), .ZN(new_n844));
  AOI21_X1  g0644(.A(KEYINPUT16), .B1(new_n316), .B2(KEYINPUT98), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n840), .B1(new_n846), .B2(new_n319), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n336), .B1(new_n846), .B2(new_n319), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n847), .A2(new_n848), .A3(new_n330), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n842), .B1(new_n849), .B2(KEYINPUT37), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n847), .B1(new_n598), .B2(new_n602), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT38), .ZN(new_n852));
  NOR3_X1   g0652(.A1(new_n850), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n342), .A2(new_n333), .A3(new_n840), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n337), .A2(new_n841), .A3(new_n330), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n337), .A2(new_n841), .A3(new_n839), .A4(new_n330), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT38), .B1(new_n854), .B2(new_n858), .ZN(new_n859));
  OAI21_X1  g0659(.A(KEYINPUT99), .B1(new_n853), .B2(new_n859), .ZN(new_n860));
  OR2_X1    g0660(.A1(new_n846), .A2(new_n319), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n342), .A2(new_n840), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g0662(.A1(new_n849), .A2(KEYINPUT37), .ZN(new_n863));
  OAI211_X1 g0663(.A(KEYINPUT38), .B(new_n862), .C1(new_n863), .C2(new_n842), .ZN(new_n864));
  INV_X1    g0664(.A(new_n858), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n841), .B1(new_n598), .B2(new_n602), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n852), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT99), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n864), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n860), .A2(new_n869), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT40), .ZN(new_n871));
  INV_X1    g0671(.A(KEYINPUT97), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n355), .A2(new_n664), .ZN(new_n873));
  OAI211_X1 g0673(.A(new_n872), .B(new_n873), .C1(new_n383), .C2(new_n376), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n383), .B2(new_n376), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT97), .ZN(new_n876));
  AOI211_X1 g0676(.A(new_n376), .B(new_n873), .C1(new_n383), .C2(new_n356), .ZN(new_n877));
  OAI211_X1 g0677(.A(new_n808), .B(new_n874), .C1(new_n876), .C2(new_n877), .ZN(new_n878));
  AOI211_X1 g0678(.A(new_n871), .B(new_n878), .C1(new_n680), .C2(new_n699), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n878), .B1(new_n680), .B2(new_n699), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n852), .B1(new_n850), .B2(new_n851), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n864), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  AOI22_X1  g0683(.A1(new_n870), .A2(new_n879), .B1(new_n883), .B2(new_n871), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n884), .B(KEYINPUT100), .Z(new_n885));
  NAND2_X1  g0685(.A1(new_n407), .A2(new_n705), .ZN(new_n886));
  OR2_X1    g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n887), .A2(G330), .A3(new_n888), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT39), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(new_n853), .B2(new_n859), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n596), .A2(new_n637), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n864), .A2(new_n881), .A3(KEYINPUT39), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n891), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n603), .A2(new_n635), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n874), .B1(new_n876), .B2(new_n877), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n806), .B(KEYINPUT96), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n897), .B1(new_n833), .B2(new_n898), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n896), .B1(new_n882), .B2(new_n899), .ZN(new_n900));
  AND3_X1   g0700(.A1(new_n629), .A2(new_n663), .A3(new_n664), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n407), .B1(new_n703), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n902), .A2(new_n606), .ZN(new_n903));
  XOR2_X1   g0703(.A(new_n900), .B(new_n903), .Z(new_n904));
  AOI21_X1  g0704(.A(new_n838), .B1(new_n889), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n904), .B2(new_n889), .ZN(new_n906));
  INV_X1    g0706(.A(new_n412), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n907), .A2(KEYINPUT35), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(KEYINPUT35), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n908), .A2(G116), .A3(new_n216), .A4(new_n909), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n910), .B(KEYINPUT36), .ZN(new_n911));
  NOR3_X1   g0711(.A1(new_n219), .A2(new_n213), .A3(new_n299), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n298), .A2(G50), .ZN(new_n913));
  OAI211_X1 g0713(.A(G1), .B(new_n713), .C1(new_n912), .C2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n906), .A2(new_n911), .A3(new_n914), .ZN(G367));
  NOR2_X1   g0715(.A1(new_n725), .A2(new_n235), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n733), .B1(new_n210), .B2(new_n388), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n717), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  OAI22_X1  g0718(.A1(new_n745), .A2(new_n774), .B1(new_n793), .B2(new_n579), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n786), .A2(G116), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT46), .Z(new_n921));
  AOI21_X1  g0721(.A(new_n324), .B1(G317), .B2(new_n743), .ZN(new_n922));
  OAI221_X1 g0722(.A(new_n922), .B1(new_n414), .B2(new_n739), .C1(new_n409), .C2(new_n747), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n740), .A2(new_n762), .B1(new_n759), .B2(new_n782), .ZN(new_n924));
  OR4_X1    g0724(.A1(new_n919), .A2(new_n921), .A3(new_n923), .A4(new_n924), .ZN(new_n925));
  OAI22_X1  g0725(.A1(new_n774), .A2(new_n202), .B1(new_n759), .B2(new_n794), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n788), .B2(new_n767), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n304), .B1(new_n747), .B2(new_n219), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT104), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n928), .A2(new_n929), .ZN(new_n931));
  AOI22_X1  g0731(.A1(G137), .A2(new_n743), .B1(new_n738), .B2(G68), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n932), .B1(new_n748), .B2(new_n297), .ZN(new_n933));
  AOI21_X1  g0733(.A(new_n933), .B1(G150), .B2(new_n754), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n927), .A2(new_n930), .A3(new_n931), .A4(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n925), .A2(new_n935), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n936), .B(KEYINPUT47), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n918), .B1(new_n937), .B2(new_n732), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n483), .A2(new_n664), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n614), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n671), .B2(new_n939), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT101), .Z(new_n942));
  NAND2_X1  g0742(.A1(new_n942), .A2(new_n731), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n938), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n644), .ZN(new_n945));
  AOI211_X1 g0745(.A(new_n945), .B(new_n652), .C1(new_n640), .C2(new_n642), .ZN(new_n946));
  INV_X1    g0746(.A(new_n650), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n640), .A2(new_n642), .A3(new_n652), .ZN(new_n948));
  NOR3_X1   g0748(.A1(new_n946), .A2(new_n947), .A3(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(new_n652), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n643), .A2(new_n644), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n650), .B1(new_n951), .B2(new_n653), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n949), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g0753(.A(new_n953), .B1(new_n701), .B2(new_n708), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n426), .A2(new_n637), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n469), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n672), .A2(new_n637), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n653), .B2(new_n654), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT44), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n959), .B(new_n960), .ZN(new_n961));
  XOR2_X1   g0761(.A(KEYINPUT102), .B(KEYINPUT45), .Z(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n958), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n963), .B1(new_n655), .B2(new_n964), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n653), .A2(new_n654), .A3(new_n958), .A4(new_n962), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n651), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n959), .B(KEYINPUT44), .ZN(new_n969));
  INV_X1    g0769(.A(new_n651), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n969), .A2(new_n970), .A3(new_n966), .A4(new_n965), .ZN(new_n971));
  NAND3_X1  g0771(.A1(new_n954), .A2(new_n968), .A3(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n972), .A2(new_n709), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n657), .B(KEYINPUT41), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT103), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n973), .A2(KEYINPUT103), .A3(new_n975), .ZN(new_n979));
  AOI21_X1  g0779(.A(new_n716), .B1(new_n978), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT43), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n942), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n948), .A2(new_n958), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n983), .A2(KEYINPUT42), .B1(new_n463), .B2(new_n664), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n654), .A2(KEYINPUT42), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n655), .A2(new_n958), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n982), .B1(new_n984), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n942), .A2(new_n981), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n987), .B(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n970), .A2(new_n964), .ZN(new_n990));
  XNOR2_X1  g0790(.A(new_n989), .B(new_n990), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n944), .B1(new_n980), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT105), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n993), .B(new_n994), .ZN(new_n995));
  INV_X1    g0795(.A(new_n995), .ZN(G387));
  INV_X1    g0796(.A(new_n953), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n703), .A2(new_n901), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n707), .B1(new_n998), .B2(new_n706), .ZN(new_n999));
  NOR3_X1   g0799(.A1(new_n678), .A2(KEYINPUT84), .A3(new_n700), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n997), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n1001), .A2(KEYINPUT108), .A3(new_n658), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT108), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n1003), .B1(new_n954), .B2(new_n657), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n701), .A2(new_n708), .A3(new_n953), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1004), .A3(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n786), .A2(new_n386), .ZN(new_n1007));
  INV_X1    g0807(.A(G150), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1007), .B1(new_n1008), .B2(new_n742), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT106), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n509), .A2(new_n738), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n324), .B1(new_n747), .B2(new_n409), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n793), .A2(new_n202), .B1(new_n762), .B2(new_n251), .ZN(new_n1014));
  INV_X1    g0814(.A(G159), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n774), .A2(new_n298), .B1(new_n759), .B2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1009), .A2(KEYINPUT106), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1010), .A2(new_n1013), .A3(new_n1017), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n324), .B1(G326), .B2(new_n743), .ZN(new_n1020));
  OAI22_X1  g0820(.A1(new_n748), .A2(new_n740), .B1(new_n739), .B2(new_n745), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(G303), .A2(new_n753), .B1(new_n754), .B2(G317), .ZN(new_n1022));
  INV_X1    g0822(.A(G322), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n1022), .B1(new_n782), .B2(new_n762), .C1(new_n1023), .C2(new_n759), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT48), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1021), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n1025), .B2(new_n1024), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT49), .ZN(new_n1028));
  OAI221_X1 g0828(.A(new_n1020), .B1(new_n485), .B2(new_n747), .C1(new_n1027), .C2(new_n1028), .ZN(new_n1029));
  AND2_X1   g0829(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1019), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT107), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n812), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1033), .B1(new_n1032), .B2(new_n1031), .ZN(new_n1034));
  AOI22_X1  g0834(.A1(new_n721), .A2(new_n659), .B1(new_n414), .B2(new_n720), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n232), .A2(new_n265), .ZN(new_n1036));
  AOI211_X1 g0836(.A(G45), .B(new_n659), .C1(G68), .C2(G77), .ZN(new_n1037));
  AOI21_X1  g0837(.A(KEYINPUT50), .B1(new_n252), .B2(new_n202), .ZN(new_n1038));
  AND3_X1   g0838(.A1(new_n252), .A2(KEYINPUT50), .A3(new_n202), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n1037), .B1(new_n1038), .B2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n724), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1035), .B1(new_n1036), .B2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n718), .B1(new_n1042), .B2(new_n733), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1034), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n646), .B2(new_n731), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n716), .B2(new_n997), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1006), .A2(new_n1046), .ZN(G393));
  NAND2_X1  g0847(.A1(new_n968), .A2(new_n971), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(KEYINPUT109), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT109), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n968), .A2(new_n1050), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1049), .A2(new_n1051), .A3(new_n716), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n725), .A2(new_n242), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n733), .B1(new_n409), .B2(new_n210), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n717), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n279), .B1(new_n742), .B2(new_n1023), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n1056), .B(new_n765), .C1(G116), .C2(new_n738), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n745), .B2(new_n748), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G317), .A2(new_n760), .B1(new_n754), .B2(G311), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT52), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n774), .A2(new_n740), .B1(new_n762), .B2(new_n579), .ZN(new_n1061));
  NOR3_X1   g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1062), .A2(KEYINPUT110), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1062), .A2(KEYINPUT110), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n793), .A2(new_n1015), .B1(new_n759), .B2(new_n1008), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT51), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n324), .B1(new_n742), .B2(new_n794), .C1(new_n739), .C2(new_n349), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1067), .B(new_n784), .C1(G68), .C2(new_n786), .ZN(new_n1068));
  AOI22_X1  g0868(.A1(G50), .A2(new_n788), .B1(new_n753), .B2(new_n252), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n1066), .A2(new_n1068), .A3(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n1063), .A2(new_n1064), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1055), .B1(new_n1071), .B2(new_n732), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n958), .B2(new_n778), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n954), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n972), .A2(new_n658), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1052), .B(new_n1073), .C1(new_n1074), .C2(new_n1075), .ZN(G390));
  OAI21_X1  g0876(.A(new_n898), .B1(new_n823), .B2(new_n824), .ZN(new_n1077));
  INV_X1    g0877(.A(new_n897), .ZN(new_n1078));
  AND3_X1   g0878(.A1(new_n700), .A2(new_n808), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1078), .B1(new_n700), .B2(new_n808), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1077), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n705), .A2(G330), .A3(new_n808), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n897), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n700), .A2(new_n808), .A3(new_n1078), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n898), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n1085), .B1(new_n677), .B2(new_n808), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1081), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n407), .A2(new_n700), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n902), .A2(new_n606), .A3(new_n1089), .ZN(new_n1090));
  INV_X1    g0890(.A(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1079), .A2(KEYINPUT111), .ZN(new_n1093));
  OR2_X1    g0893(.A1(new_n1079), .A2(KEYINPUT111), .ZN(new_n1094));
  AND2_X1   g0894(.A1(new_n891), .A2(new_n893), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1096));
  INV_X1    g0896(.A(new_n892), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1095), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n860), .A2(new_n869), .A3(new_n1097), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n702), .A2(new_n664), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n898), .B1(new_n1100), .B2(new_n809), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1099), .B1(new_n1078), .B2(new_n1101), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1093), .B(new_n1094), .C1(new_n1098), .C2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n891), .A2(new_n893), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n899), .B2(new_n892), .ZN(new_n1105));
  OAI211_X1 g0905(.A(new_n870), .B(new_n1097), .C1(new_n897), .C2(new_n1086), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1105), .A2(KEYINPUT111), .A3(new_n1106), .A4(new_n1079), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1092), .B1(new_n1103), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1103), .A2(new_n1107), .A3(new_n1092), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1109), .A2(new_n658), .A3(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(new_n716), .ZN(new_n1113));
  INV_X1    g0913(.A(G125), .ZN(new_n1114));
  OAI221_X1 g0914(.A(new_n304), .B1(new_n1114), .B2(new_n742), .C1(new_n747), .C2(new_n202), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(G128), .A2(new_n760), .B1(new_n754), .B2(G132), .ZN(new_n1116));
  NOR2_X1   g0916(.A1(new_n748), .A2(new_n1008), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(KEYINPUT53), .ZN(new_n1119));
  AOI211_X1 g0919(.A(new_n1115), .B(new_n1119), .C1(KEYINPUT53), .C2(new_n1118), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n788), .A2(G137), .ZN(new_n1121));
  XNOR2_X1  g0921(.A(KEYINPUT54), .B(G143), .ZN(new_n1122));
  OAI221_X1 g0922(.A(new_n1121), .B1(new_n1015), .B2(new_n739), .C1(new_n774), .C2(new_n1122), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT112), .Z(new_n1124));
  NAND2_X1  g0924(.A1(new_n1120), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  AND2_X1   g0926(.A1(new_n1126), .A2(KEYINPUT113), .ZN(new_n1127));
  NOR2_X1   g0927(.A1(new_n1126), .A2(KEYINPUT113), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(G97), .A2(new_n753), .B1(new_n754), .B2(G116), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n414), .B2(new_n762), .C1(new_n745), .C2(new_n759), .ZN(new_n1130));
  OAI221_X1 g0930(.A(new_n279), .B1(new_n740), .B2(new_n742), .C1(new_n739), .C2(new_n349), .ZN(new_n1131));
  NOR4_X1   g0931(.A1(new_n1130), .A2(new_n771), .A3(new_n799), .A4(new_n1131), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n1127), .A2(new_n1128), .A3(new_n1132), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n717), .B1(new_n252), .B2(new_n815), .C1(new_n1133), .C2(new_n812), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1134), .B1(new_n1104), .B2(new_n810), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT114), .B1(new_n1113), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT114), .ZN(new_n1138));
  AOI211_X1 g0938(.A(new_n1138), .B(new_n1135), .C1(new_n1112), .C2(new_n716), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1111), .B1(new_n1137), .B2(new_n1139), .ZN(G378));
  INV_X1    g0940(.A(KEYINPUT57), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1090), .B1(new_n1112), .B2(new_n1088), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n883), .A2(new_n871), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n880), .A2(new_n860), .A3(KEYINPUT40), .A4(new_n869), .ZN(new_n1144));
  NAND3_X1  g0944(.A1(new_n1143), .A2(new_n1144), .A3(G330), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n291), .A2(new_n294), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n260), .A2(new_n635), .ZN(new_n1147));
  XNOR2_X1  g0947(.A(new_n1146), .B(new_n1147), .ZN(new_n1148));
  XNOR2_X1  g0948(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1148), .B(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1145), .A2(new_n1152), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1151), .A2(new_n1143), .A3(G330), .A4(new_n1144), .ZN(new_n1154));
  AND3_X1   g0954(.A1(new_n1153), .A2(new_n900), .A3(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(new_n900), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1156));
  NOR2_X1   g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1141), .B1(new_n1142), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n900), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1151), .B1(new_n884), .B2(G330), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1154), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1159), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1153), .A2(new_n900), .A3(new_n1154), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1162), .A2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1164), .B(KEYINPUT57), .C1(new_n1090), .C2(new_n1108), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1158), .A2(new_n658), .A3(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT116), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n715), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1152), .A2(new_n810), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n717), .B1(new_n815), .B2(G50), .ZN(new_n1170));
  OAI22_X1  g0970(.A1(new_n748), .A2(new_n1122), .B1(new_n739), .B2(new_n1008), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(G128), .A2(new_n754), .B1(new_n753), .B2(G137), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n1114), .B2(new_n759), .ZN(new_n1173));
  AOI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(G132), .C2(new_n788), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(G33), .A2(G41), .ZN(new_n1178));
  XNOR2_X1  g0978(.A(new_n1178), .B(KEYINPUT115), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n747), .A2(new_n766), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G124), .C2(new_n743), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1176), .A2(new_n1177), .A3(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n509), .A2(new_n753), .B1(new_n760), .B2(G116), .ZN(new_n1183));
  OAI221_X1 g0983(.A(new_n1183), .B1(new_n409), .B2(new_n762), .C1(new_n414), .C2(new_n793), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1007), .B1(new_n298), .B2(new_n739), .C1(new_n745), .C2(new_n742), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n312), .A2(new_n264), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n747), .A2(new_n297), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .A4(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1186), .A2(new_n202), .A3(new_n1179), .ZN(new_n1190));
  OR2_X1    g0990(.A1(new_n1188), .A2(KEYINPUT58), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1182), .A2(new_n1189), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1170), .B1(new_n1192), .B2(new_n732), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1169), .A2(new_n1193), .ZN(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1167), .B1(new_n1168), .B2(new_n1195), .ZN(new_n1196));
  OAI211_X1 g0996(.A(KEYINPUT116), .B(new_n1194), .C1(new_n1157), .C2(new_n715), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(new_n1197), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1166), .A2(new_n1198), .ZN(G375));
  XOR2_X1   g0999(.A(new_n715), .B(KEYINPUT117), .Z(new_n1200));
  NOR3_X1   g1000(.A1(new_n1079), .A2(new_n1080), .A3(new_n1101), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n1083), .A2(new_n1084), .B1(new_n833), .B2(new_n898), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1200), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G116), .A2(new_n788), .B1(new_n753), .B2(G107), .ZN(new_n1204));
  OAI221_X1 g1004(.A(new_n1204), .B1(new_n745), .B2(new_n793), .C1(new_n740), .C2(new_n759), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n279), .B1(new_n742), .B2(new_n579), .ZN(new_n1206));
  OAI22_X1  g1006(.A1(new_n349), .A2(new_n747), .B1(new_n748), .B2(new_n409), .ZN(new_n1207));
  NOR4_X1   g1007(.A1(new_n1205), .A2(new_n1011), .A3(new_n1206), .A4(new_n1207), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT118), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n739), .A2(new_n202), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n312), .B(new_n1211), .C1(G128), .C2(new_n743), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1187), .B1(G159), .B2(new_n786), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G132), .A2(new_n760), .B1(new_n754), .B2(G137), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1122), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n788), .A2(new_n1215), .B1(new_n753), .B2(G150), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1216), .ZN(new_n1217));
  INV_X1    g1017(.A(KEYINPUT118), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1217), .B1(new_n1208), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n732), .B1(new_n1210), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n815), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n718), .B1(new_n1221), .B2(new_n298), .ZN(new_n1222));
  OAI211_X1 g1022(.A(new_n1220), .B(new_n1222), .C1(new_n1078), .C2(new_n813), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1203), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1081), .A2(new_n1090), .A3(new_n1087), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1092), .A2(new_n975), .A3(new_n1226), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1225), .A2(new_n1227), .ZN(G381));
  AND3_X1   g1028(.A1(new_n1006), .A2(new_n780), .A3(new_n1046), .ZN(new_n1229));
  NOR3_X1   g1029(.A1(G390), .A2(G384), .A3(G381), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n995), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT119), .ZN(new_n1232));
  OR2_X1    g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1135), .B1(new_n1112), .B2(new_n716), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1111), .A2(new_n1235), .ZN(new_n1236));
  NOR2_X1   g1036(.A1(G375), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1233), .A2(new_n1234), .A3(new_n1237), .ZN(G407));
  INV_X1    g1038(.A(G213), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1239), .B1(new_n1237), .B2(new_n636), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(G407), .A2(new_n1240), .ZN(G409));
  AOI21_X1  g1041(.A(new_n780), .B1(new_n1006), .B2(new_n1046), .ZN(new_n1242));
  OAI21_X1  g1042(.A(G390), .B1(new_n1229), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(G393), .A2(G396), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1006), .A2(new_n780), .A3(new_n1046), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n994), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1246), .B2(G390), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n944), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n978), .A2(new_n979), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n715), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1248), .B1(new_n1250), .B2(new_n991), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g1052(.A(KEYINPUT105), .B1(new_n1229), .B2(new_n1242), .ZN(new_n1253));
  INV_X1    g1053(.A(G390), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n993), .A2(new_n1255), .A3(new_n1243), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1239), .A2(G343), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1166), .A2(G378), .A3(new_n1198), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1195), .B1(new_n1164), .B2(new_n1200), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1164), .B1(new_n1090), .B2(new_n1108), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1260), .B1(new_n1261), .B2(new_n974), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1262), .A2(new_n1111), .A3(new_n1235), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1258), .B1(new_n1259), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1090), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT60), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1226), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND4_X1  g1067(.A1(new_n1081), .A2(new_n1090), .A3(new_n1087), .A4(KEYINPUT60), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1268), .A2(new_n658), .ZN(new_n1269));
  AOI211_X1 g1069(.A(new_n836), .B(new_n1224), .C1(new_n1267), .C2(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G384), .B1(new_n1271), .B2(new_n1225), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1270), .A2(new_n1272), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1264), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1257), .B1(new_n1274), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1268), .A2(new_n658), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1092), .A2(KEYINPUT60), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1277), .B1(new_n1278), .B2(new_n1226), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n836), .B1(new_n1279), .B2(new_n1224), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1271), .A2(G384), .A3(new_n1225), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1258), .A2(KEYINPUT120), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1280), .A2(new_n1281), .A3(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(KEYINPUT121), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1258), .A2(G2897), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1285), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT121), .ZN(new_n1287));
  NAND4_X1  g1087(.A1(new_n1280), .A2(new_n1281), .A3(new_n1287), .A4(new_n1282), .ZN(new_n1288));
  AND3_X1   g1088(.A1(new_n1284), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1286), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1289), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1264), .ZN(new_n1292));
  AOI21_X1  g1092(.A(KEYINPUT61), .B1(new_n1291), .B2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1264), .A2(KEYINPUT63), .A3(new_n1273), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1276), .A2(new_n1293), .A3(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT61), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1287), .B1(new_n1273), .B2(new_n1282), .ZN(new_n1297));
  INV_X1    g1097(.A(new_n1288), .ZN(new_n1298));
  OAI21_X1  g1098(.A(new_n1285), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1284), .A2(new_n1286), .A3(new_n1288), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  OAI21_X1  g1101(.A(new_n1296), .B1(new_n1301), .B2(new_n1264), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1259), .A2(new_n1263), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1258), .ZN(new_n1304));
  XOR2_X1   g1104(.A(KEYINPUT122), .B(KEYINPUT62), .Z(new_n1305));
  AND4_X1   g1105(.A1(new_n1273), .A2(new_n1303), .A3(new_n1304), .A4(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(KEYINPUT122), .A2(KEYINPUT62), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(new_n1264), .B2(new_n1273), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1302), .A2(new_n1306), .A3(new_n1308), .ZN(new_n1309));
  AND3_X1   g1109(.A1(new_n1252), .A2(KEYINPUT123), .A3(new_n1256), .ZN(new_n1310));
  AOI21_X1  g1110(.A(KEYINPUT123), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1311));
  OAI21_X1  g1111(.A(KEYINPUT124), .B1(new_n1310), .B2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT123), .ZN(new_n1313));
  NOR2_X1   g1113(.A1(new_n1247), .A2(new_n1251), .ZN(new_n1314));
  AOI21_X1  g1114(.A(new_n993), .B1(new_n1255), .B2(new_n1243), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1313), .B1(new_n1314), .B2(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(KEYINPUT124), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1252), .A2(KEYINPUT123), .A3(new_n1256), .ZN(new_n1318));
  NAND3_X1  g1118(.A1(new_n1316), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1312), .A2(new_n1319), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1295), .B1(new_n1309), .B2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1321), .A2(KEYINPUT125), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT125), .ZN(new_n1323));
  OAI211_X1 g1123(.A(new_n1323), .B(new_n1295), .C1(new_n1309), .C2(new_n1320), .ZN(new_n1324));
  NAND2_X1  g1124(.A1(new_n1322), .A2(new_n1324), .ZN(G405));
  INV_X1    g1125(.A(G375), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1259), .B1(new_n1326), .B2(new_n1236), .ZN(new_n1327));
  OAI21_X1  g1127(.A(KEYINPUT126), .B1(new_n1270), .B2(new_n1272), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1327), .A2(new_n1328), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT126), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1273), .A2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1331), .A2(new_n1328), .ZN(new_n1332));
  OAI211_X1 g1132(.A(new_n1332), .B(new_n1259), .C1(new_n1326), .C2(new_n1236), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1329), .A2(new_n1333), .ZN(new_n1334));
  INV_X1    g1134(.A(new_n1334), .ZN(new_n1335));
  NAND2_X1  g1135(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1336));
  OAI21_X1  g1136(.A(KEYINPUT127), .B1(new_n1335), .B2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1339));
  NOR3_X1   g1139(.A1(new_n1335), .A2(KEYINPUT127), .A3(new_n1336), .ZN(new_n1340));
  NOR2_X1   g1140(.A1(new_n1339), .A2(new_n1340), .ZN(G402));
endmodule


