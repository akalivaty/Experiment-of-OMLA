

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596;

  INV_X1 U324 ( .A(G22GAT), .ZN(n371) );
  XNOR2_X1 U325 ( .A(n425), .B(n424), .ZN(n524) );
  XNOR2_X1 U326 ( .A(KEYINPUT37), .B(KEYINPUT105), .ZN(n424) );
  XNOR2_X1 U327 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U328 ( .A(n482), .B(n481), .ZN(n548) );
  XNOR2_X1 U329 ( .A(KEYINPUT38), .B(n461), .ZN(n510) );
  NOR2_X1 U330 ( .A1(n470), .A2(n558), .ZN(n471) );
  XNOR2_X1 U331 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U332 ( .A(n374), .B(n373), .ZN(n375) );
  INV_X1 U333 ( .A(KEYINPUT116), .ZN(n480) );
  INV_X1 U334 ( .A(n442), .ZN(n385) );
  XNOR2_X1 U335 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n483) );
  XNOR2_X1 U336 ( .A(n480), .B(KEYINPUT48), .ZN(n481) );
  NOR2_X1 U337 ( .A1(n422), .A2(n421), .ZN(n491) );
  XNOR2_X1 U338 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U339 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U340 ( .A(n388), .B(n387), .ZN(n486) );
  XNOR2_X1 U341 ( .A(n440), .B(n439), .ZN(n444) );
  INV_X1 U342 ( .A(G43GAT), .ZN(n462) );
  NOR2_X1 U343 ( .A1(n589), .A2(n567), .ZN(n568) );
  XNOR2_X1 U344 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U345 ( .A(n465), .B(n464), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT83), .B(KEYINPUT20), .Z(n293) );
  XNOR2_X1 U347 ( .A(G169GAT), .B(KEYINPUT84), .ZN(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U349 ( .A(KEYINPUT85), .B(G176GAT), .Z(n295) );
  XNOR2_X1 U350 ( .A(G99GAT), .B(KEYINPUT86), .ZN(n294) );
  XNOR2_X1 U351 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U352 ( .A(n297), .B(n296), .Z(n303) );
  XOR2_X1 U353 ( .A(KEYINPUT82), .B(KEYINPUT0), .Z(n299) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(G134GAT), .ZN(n298) );
  XNOR2_X1 U355 ( .A(n299), .B(n298), .ZN(n407) );
  XOR2_X1 U356 ( .A(G183GAT), .B(KEYINPUT19), .Z(n301) );
  XNOR2_X1 U357 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n300) );
  XNOR2_X1 U358 ( .A(n301), .B(n300), .ZN(n366) );
  XNOR2_X1 U359 ( .A(n407), .B(n366), .ZN(n302) );
  XNOR2_X1 U360 ( .A(n303), .B(n302), .ZN(n307) );
  XOR2_X1 U361 ( .A(G15GAT), .B(G127GAT), .Z(n350) );
  XOR2_X1 U362 ( .A(G120GAT), .B(G71GAT), .Z(n434) );
  XOR2_X1 U363 ( .A(n350), .B(n434), .Z(n305) );
  NAND2_X1 U364 ( .A1(G227GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U365 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U366 ( .A(n307), .B(n306), .Z(n309) );
  XNOR2_X1 U367 ( .A(G43GAT), .B(G190GAT), .ZN(n308) );
  XNOR2_X1 U368 ( .A(n309), .B(n308), .ZN(n569) );
  XOR2_X1 U369 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n311) );
  XNOR2_X1 U370 ( .A(G92GAT), .B(KEYINPUT10), .ZN(n310) );
  XNOR2_X1 U371 ( .A(n311), .B(n310), .ZN(n316) );
  INV_X1 U372 ( .A(G85GAT), .ZN(n312) );
  NAND2_X1 U373 ( .A1(G99GAT), .A2(n312), .ZN(n315) );
  INV_X1 U374 ( .A(G99GAT), .ZN(n313) );
  NAND2_X1 U375 ( .A1(n313), .A2(G85GAT), .ZN(n314) );
  NAND2_X1 U376 ( .A1(n315), .A2(n314), .ZN(n427) );
  XOR2_X1 U377 ( .A(n316), .B(n427), .Z(n318) );
  XNOR2_X1 U378 ( .A(G218GAT), .B(G106GAT), .ZN(n317) );
  XNOR2_X1 U379 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U380 ( .A(G36GAT), .B(G190GAT), .Z(n355) );
  XNOR2_X1 U381 ( .A(G50GAT), .B(KEYINPUT76), .ZN(n319) );
  XNOR2_X1 U382 ( .A(n319), .B(G162GAT), .ZN(n382) );
  XOR2_X1 U383 ( .A(n355), .B(n382), .Z(n321) );
  NAND2_X1 U384 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U385 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U386 ( .A(n323), .B(n322), .Z(n331) );
  XOR2_X1 U387 ( .A(KEYINPUT7), .B(KEYINPUT8), .Z(n325) );
  XNOR2_X1 U388 ( .A(G43GAT), .B(G29GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U390 ( .A(KEYINPUT68), .B(n326), .Z(n460) );
  XOR2_X1 U391 ( .A(KEYINPUT78), .B(KEYINPUT11), .Z(n328) );
  XNOR2_X1 U392 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n460), .B(n329), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n571) );
  XOR2_X1 U396 ( .A(KEYINPUT36), .B(n571), .Z(n592) );
  XOR2_X1 U397 ( .A(KEYINPUT80), .B(G64GAT), .Z(n333) );
  XNOR2_X1 U398 ( .A(G8GAT), .B(G183GAT), .ZN(n332) );
  XNOR2_X1 U399 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U400 ( .A(KEYINPUT79), .B(KEYINPUT81), .Z(n335) );
  XNOR2_X1 U401 ( .A(KEYINPUT14), .B(KEYINPUT12), .ZN(n334) );
  XNOR2_X1 U402 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U403 ( .A(n337), .B(n336), .ZN(n354) );
  XOR2_X1 U404 ( .A(G78GAT), .B(G155GAT), .Z(n339) );
  XNOR2_X1 U405 ( .A(G71GAT), .B(G211GAT), .ZN(n338) );
  XNOR2_X1 U406 ( .A(n339), .B(n338), .ZN(n345) );
  XOR2_X1 U407 ( .A(KEYINPUT69), .B(KEYINPUT70), .Z(n341) );
  XNOR2_X1 U408 ( .A(G22GAT), .B(G1GAT), .ZN(n340) );
  XNOR2_X1 U409 ( .A(n341), .B(n340), .ZN(n454) );
  XOR2_X1 U410 ( .A(KEYINPUT15), .B(n454), .Z(n343) );
  NAND2_X1 U411 ( .A1(G231GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U412 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U413 ( .A(n345), .B(n344), .Z(n352) );
  INV_X1 U414 ( .A(KEYINPUT13), .ZN(n346) );
  NAND2_X1 U415 ( .A1(n346), .A2(G57GAT), .ZN(n349) );
  INV_X1 U416 ( .A(G57GAT), .ZN(n347) );
  NAND2_X1 U417 ( .A1(n347), .A2(KEYINPUT13), .ZN(n348) );
  NAND2_X1 U418 ( .A1(n349), .A2(n348), .ZN(n426) );
  XNOR2_X1 U419 ( .A(n350), .B(n426), .ZN(n351) );
  XNOR2_X1 U420 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U421 ( .A(n354), .B(n353), .ZN(n558) );
  XOR2_X1 U422 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n359) );
  XOR2_X1 U423 ( .A(G169GAT), .B(G8GAT), .Z(n450) );
  NAND2_X1 U424 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U426 ( .A(n450), .B(n357), .ZN(n358) );
  XNOR2_X1 U427 ( .A(n359), .B(n358), .ZN(n361) );
  XNOR2_X1 U428 ( .A(G176GAT), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U429 ( .A(n360), .B(G64GAT), .ZN(n441) );
  XOR2_X1 U430 ( .A(n361), .B(n441), .Z(n368) );
  XNOR2_X1 U431 ( .A(G211GAT), .B(G218GAT), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n362), .B(KEYINPUT21), .ZN(n363) );
  XOR2_X1 U433 ( .A(n363), .B(KEYINPUT89), .Z(n365) );
  XNOR2_X1 U434 ( .A(G197GAT), .B(G204GAT), .ZN(n364) );
  XNOR2_X1 U435 ( .A(n365), .B(n364), .ZN(n383) );
  XNOR2_X1 U436 ( .A(n366), .B(n383), .ZN(n367) );
  XNOR2_X1 U437 ( .A(n368), .B(n367), .ZN(n529) );
  XNOR2_X1 U438 ( .A(n529), .B(KEYINPUT27), .ZN(n419) );
  XOR2_X1 U439 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n370) );
  XNOR2_X1 U440 ( .A(KEYINPUT87), .B(KEYINPUT88), .ZN(n369) );
  XNOR2_X1 U441 ( .A(n370), .B(n369), .ZN(n374) );
  NAND2_X1 U442 ( .A1(G228GAT), .A2(G233GAT), .ZN(n372) );
  XOR2_X1 U443 ( .A(n375), .B(KEYINPUT22), .Z(n381) );
  XNOR2_X1 U444 ( .A(KEYINPUT91), .B(KEYINPUT2), .ZN(n376) );
  XNOR2_X1 U445 ( .A(n376), .B(KEYINPUT3), .ZN(n377) );
  XOR2_X1 U446 ( .A(n377), .B(KEYINPUT90), .Z(n379) );
  XNOR2_X1 U447 ( .A(G141GAT), .B(G155GAT), .ZN(n378) );
  XNOR2_X1 U448 ( .A(n379), .B(n378), .ZN(n411) );
  XNOR2_X1 U449 ( .A(n411), .B(KEYINPUT92), .ZN(n380) );
  XNOR2_X1 U450 ( .A(n381), .B(n380), .ZN(n388) );
  XNOR2_X1 U451 ( .A(n383), .B(n382), .ZN(n386) );
  XNOR2_X1 U452 ( .A(G106GAT), .B(G78GAT), .ZN(n384) );
  XNOR2_X1 U453 ( .A(n384), .B(G148GAT), .ZN(n442) );
  NOR2_X1 U454 ( .A1(n569), .A2(n486), .ZN(n389) );
  XOR2_X1 U455 ( .A(KEYINPUT101), .B(n389), .Z(n390) );
  XNOR2_X1 U456 ( .A(KEYINPUT26), .B(n390), .ZN(n577) );
  NAND2_X1 U457 ( .A1(n419), .A2(n577), .ZN(n394) );
  NAND2_X1 U458 ( .A1(n569), .A2(n529), .ZN(n391) );
  NAND2_X1 U459 ( .A1(n486), .A2(n391), .ZN(n392) );
  XOR2_X1 U460 ( .A(KEYINPUT25), .B(n392), .Z(n393) );
  NAND2_X1 U461 ( .A1(n394), .A2(n393), .ZN(n417) );
  XOR2_X1 U462 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n396) );
  XNOR2_X1 U463 ( .A(G127GAT), .B(G120GAT), .ZN(n395) );
  XNOR2_X1 U464 ( .A(n396), .B(n395), .ZN(n400) );
  XOR2_X1 U465 ( .A(G85GAT), .B(G148GAT), .Z(n398) );
  XNOR2_X1 U466 ( .A(G29GAT), .B(G162GAT), .ZN(n397) );
  XNOR2_X1 U467 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U468 ( .A(n400), .B(n399), .ZN(n415) );
  XOR2_X1 U469 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n402) );
  XNOR2_X1 U470 ( .A(KEYINPUT4), .B(KEYINPUT97), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n406) );
  XOR2_X1 U472 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n404) );
  XNOR2_X1 U473 ( .A(G1GAT), .B(G57GAT), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U475 ( .A(n406), .B(n405), .Z(n413) );
  XOR2_X1 U476 ( .A(n407), .B(KEYINPUT6), .Z(n409) );
  NAND2_X1 U477 ( .A1(G225GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U478 ( .A(n409), .B(n408), .ZN(n410) );
  XNOR2_X1 U479 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n413), .B(n412), .ZN(n414) );
  XNOR2_X1 U481 ( .A(n415), .B(n414), .ZN(n527) );
  INV_X1 U482 ( .A(n527), .ZN(n416) );
  NAND2_X1 U483 ( .A1(n417), .A2(n416), .ZN(n418) );
  XOR2_X1 U484 ( .A(KEYINPUT102), .B(n418), .Z(n422) );
  AND2_X1 U485 ( .A1(n419), .A2(n527), .ZN(n549) );
  XNOR2_X1 U486 ( .A(n486), .B(KEYINPUT28), .ZN(n501) );
  NAND2_X1 U487 ( .A1(n549), .A2(n501), .ZN(n538) );
  NOR2_X1 U488 ( .A1(n569), .A2(n538), .ZN(n420) );
  XNOR2_X1 U489 ( .A(n420), .B(KEYINPUT100), .ZN(n421) );
  NOR2_X1 U490 ( .A1(n558), .A2(n491), .ZN(n423) );
  NAND2_X1 U491 ( .A1(n592), .A2(n423), .ZN(n425) );
  XOR2_X1 U492 ( .A(KEYINPUT73), .B(n426), .Z(n429) );
  XNOR2_X1 U493 ( .A(G204GAT), .B(n427), .ZN(n428) );
  XNOR2_X1 U494 ( .A(n429), .B(n428), .ZN(n433) );
  XOR2_X1 U495 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n431) );
  NAND2_X1 U496 ( .A1(G230GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n440) );
  XOR2_X1 U499 ( .A(n434), .B(KEYINPUT31), .Z(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT32), .B(KEYINPUT75), .Z(n436) );
  XNOR2_X1 U501 ( .A(KEYINPUT71), .B(KEYINPUT74), .ZN(n435) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U503 ( .A(n442), .B(n441), .Z(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n584) );
  XOR2_X1 U505 ( .A(KEYINPUT29), .B(KEYINPUT66), .Z(n446) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(G113GAT), .ZN(n445) );
  XNOR2_X1 U507 ( .A(n446), .B(n445), .ZN(n458) );
  XOR2_X1 U508 ( .A(G141GAT), .B(G197GAT), .Z(n448) );
  XNOR2_X1 U509 ( .A(G50GAT), .B(G36GAT), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U511 ( .A(n450), .B(n449), .Z(n452) );
  NAND2_X1 U512 ( .A1(G229GAT), .A2(G233GAT), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U514 ( .A(n453), .B(KEYINPUT30), .Z(n456) );
  XNOR2_X1 U515 ( .A(n454), .B(KEYINPUT67), .ZN(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U518 ( .A(n460), .B(n459), .ZN(n579) );
  INV_X1 U519 ( .A(n579), .ZN(n552) );
  NAND2_X1 U520 ( .A1(n584), .A2(n552), .ZN(n494) );
  NOR2_X1 U521 ( .A1(n524), .A2(n494), .ZN(n461) );
  NAND2_X1 U522 ( .A1(n569), .A2(n510), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT108), .B(KEYINPUT40), .Z(n463) );
  XOR2_X1 U524 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n467) );
  XNOR2_X1 U525 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n466) );
  XOR2_X1 U526 ( .A(n467), .B(n466), .Z(n489) );
  XOR2_X1 U527 ( .A(n584), .B(KEYINPUT64), .Z(n468) );
  XNOR2_X1 U528 ( .A(KEYINPUT41), .B(n468), .ZN(n513) );
  NOR2_X1 U529 ( .A1(n579), .A2(n513), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT46), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n471), .B(KEYINPUT114), .ZN(n472) );
  NAND2_X1 U532 ( .A1(n472), .A2(n571), .ZN(n473) );
  XNOR2_X1 U533 ( .A(n473), .B(KEYINPUT47), .ZN(n479) );
  XOR2_X1 U534 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n475) );
  NAND2_X1 U535 ( .A1(n558), .A2(n592), .ZN(n474) );
  XNOR2_X1 U536 ( .A(n475), .B(n474), .ZN(n477) );
  NAND2_X1 U537 ( .A1(n584), .A2(n579), .ZN(n476) );
  NOR2_X1 U538 ( .A1(n477), .A2(n476), .ZN(n478) );
  NOR2_X1 U539 ( .A1(n479), .A2(n478), .ZN(n482) );
  NAND2_X1 U540 ( .A1(n548), .A2(n529), .ZN(n484) );
  NOR2_X1 U541 ( .A1(n527), .A2(n485), .ZN(n578) );
  NAND2_X1 U542 ( .A1(n486), .A2(n578), .ZN(n487) );
  XNOR2_X1 U543 ( .A(n487), .B(KEYINPUT55), .ZN(n573) );
  NAND2_X1 U544 ( .A1(n573), .A2(n569), .ZN(n567) );
  NOR2_X1 U545 ( .A1(n567), .A2(n513), .ZN(n488) );
  XNOR2_X1 U546 ( .A(n489), .B(n488), .ZN(G1349GAT) );
  INV_X1 U547 ( .A(n571), .ZN(n561) );
  INV_X1 U548 ( .A(n558), .ZN(n589) );
  NOR2_X1 U549 ( .A1(n561), .A2(n589), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n490), .B(KEYINPUT16), .ZN(n493) );
  INV_X1 U551 ( .A(n491), .ZN(n492) );
  NAND2_X1 U552 ( .A1(n493), .A2(n492), .ZN(n514) );
  NOR2_X1 U553 ( .A1(n494), .A2(n514), .ZN(n502) );
  NAND2_X1 U554 ( .A1(n502), .A2(n527), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(KEYINPUT34), .ZN(n496) );
  XNOR2_X1 U556 ( .A(G1GAT), .B(n496), .ZN(G1324GAT) );
  XOR2_X1 U557 ( .A(G8GAT), .B(KEYINPUT103), .Z(n498) );
  NAND2_X1 U558 ( .A1(n502), .A2(n529), .ZN(n497) );
  XNOR2_X1 U559 ( .A(n498), .B(n497), .ZN(G1325GAT) );
  XOR2_X1 U560 ( .A(G15GAT), .B(KEYINPUT35), .Z(n500) );
  NAND2_X1 U561 ( .A1(n502), .A2(n569), .ZN(n499) );
  XNOR2_X1 U562 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  INV_X1 U563 ( .A(n501), .ZN(n533) );
  NAND2_X1 U564 ( .A1(n502), .A2(n533), .ZN(n503) );
  XNOR2_X1 U565 ( .A(n503), .B(KEYINPUT104), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G22GAT), .B(n504), .ZN(G1327GAT) );
  XOR2_X1 U567 ( .A(G29GAT), .B(KEYINPUT39), .Z(n506) );
  NAND2_X1 U568 ( .A1(n527), .A2(n510), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(KEYINPUT106), .B(n507), .ZN(G1328GAT) );
  XOR2_X1 U571 ( .A(G36GAT), .B(KEYINPUT107), .Z(n509) );
  NAND2_X1 U572 ( .A1(n529), .A2(n510), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(G1329GAT) );
  XOR2_X1 U574 ( .A(G50GAT), .B(KEYINPUT109), .Z(n512) );
  NAND2_X1 U575 ( .A1(n533), .A2(n510), .ZN(n511) );
  XNOR2_X1 U576 ( .A(n512), .B(n511), .ZN(G1331GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT42), .B(KEYINPUT110), .Z(n516) );
  INV_X1 U578 ( .A(n513), .ZN(n554) );
  NAND2_X1 U579 ( .A1(n579), .A2(n554), .ZN(n525) );
  NOR2_X1 U580 ( .A1(n525), .A2(n514), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n521), .A2(n527), .ZN(n515) );
  XNOR2_X1 U582 ( .A(n516), .B(n515), .ZN(n517) );
  XOR2_X1 U583 ( .A(G57GAT), .B(n517), .Z(G1332GAT) );
  XOR2_X1 U584 ( .A(G64GAT), .B(KEYINPUT111), .Z(n519) );
  NAND2_X1 U585 ( .A1(n521), .A2(n529), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(G1333GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n569), .ZN(n520) );
  XNOR2_X1 U588 ( .A(n520), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U589 ( .A(G78GAT), .B(KEYINPUT43), .Z(n523) );
  NAND2_X1 U590 ( .A1(n521), .A2(n533), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n526), .B(KEYINPUT112), .ZN(n532) );
  NAND2_X1 U594 ( .A1(n527), .A2(n532), .ZN(n528) );
  XNOR2_X1 U595 ( .A(G85GAT), .B(n528), .ZN(G1336GAT) );
  NAND2_X1 U596 ( .A1(n532), .A2(n529), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n530), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U598 ( .A1(n532), .A2(n569), .ZN(n531) );
  XNOR2_X1 U599 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U600 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n535) );
  NAND2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(G106GAT), .B(n536), .ZN(G1339GAT) );
  NAND2_X1 U604 ( .A1(n569), .A2(n548), .ZN(n537) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n552), .A2(n544), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U609 ( .A1(n544), .A2(n554), .ZN(n540) );
  XNOR2_X1 U610 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  NAND2_X1 U611 ( .A1(n544), .A2(n558), .ZN(n542) );
  XNOR2_X1 U612 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U613 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n546) );
  NAND2_X1 U615 ( .A1(n544), .A2(n561), .ZN(n545) );
  XNOR2_X1 U616 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U617 ( .A(G134GAT), .B(n547), .Z(G1343GAT) );
  INV_X1 U618 ( .A(n548), .ZN(n551) );
  NAND2_X1 U619 ( .A1(n549), .A2(n577), .ZN(n550) );
  NOR2_X1 U620 ( .A1(n551), .A2(n550), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n562), .A2(n552), .ZN(n553) );
  XNOR2_X1 U622 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U624 ( .A1(n562), .A2(n554), .ZN(n555) );
  XNOR2_X1 U625 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n558), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n559), .B(KEYINPUT118), .ZN(n560) );
  XNOR2_X1 U629 ( .A(G155GAT), .B(n560), .ZN(G1346GAT) );
  XOR2_X1 U630 ( .A(G162GAT), .B(KEYINPUT119), .Z(n564) );
  NAND2_X1 U631 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U632 ( .A(n564), .B(n563), .ZN(G1347GAT) );
  NOR2_X1 U633 ( .A1(n579), .A2(n567), .ZN(n566) );
  XNOR2_X1 U634 ( .A(G169GAT), .B(KEYINPUT121), .ZN(n565) );
  XNOR2_X1 U635 ( .A(n566), .B(n565), .ZN(G1348GAT) );
  XOR2_X1 U636 ( .A(G183GAT), .B(n568), .Z(G1350GAT) );
  INV_X1 U637 ( .A(n569), .ZN(n570) );
  NOR2_X1 U638 ( .A1(n571), .A2(n570), .ZN(n572) );
  AND2_X1 U639 ( .A1(n573), .A2(n572), .ZN(n575) );
  XNOR2_X1 U640 ( .A(KEYINPUT123), .B(KEYINPUT58), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(G190GAT), .B(n576), .ZN(G1351GAT) );
  XNOR2_X1 U643 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n583) );
  NAND2_X1 U644 ( .A1(n578), .A2(n577), .ZN(n591) );
  NOR2_X1 U645 ( .A1(n579), .A2(n591), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(G1352GAT) );
  NOR2_X1 U649 ( .A1(n591), .A2(n584), .ZN(n588) );
  XOR2_X1 U650 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n586) );
  XNOR2_X1 U651 ( .A(G204GAT), .B(KEYINPUT126), .ZN(n585) );
  XNOR2_X1 U652 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(G1353GAT) );
  NOR2_X1 U654 ( .A1(n589), .A2(n591), .ZN(n590) );
  XOR2_X1 U655 ( .A(G211GAT), .B(n590), .Z(G1354GAT) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n595) );
  INV_X1 U657 ( .A(n591), .ZN(n593) );
  NAND2_X1 U658 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U659 ( .A(n595), .B(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(G218GAT), .B(n596), .ZN(G1355GAT) );
endmodule

