//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 1 0 1 0 1 0 1 0 0 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:45 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n578, new_n579, new_n581,
    new_n582, new_n583, new_n584, new_n585, new_n586, new_n587, new_n588,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n598, new_n599, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1252, new_n1253, new_n1254,
    new_n1255, new_n1256, new_n1257, new_n1258, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1264, new_n1267;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G125), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n461), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  AND2_X1   g040(.A1(G113), .A2(G2104), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G137), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  OAI21_X1  g046(.A(KEYINPUT64), .B1(new_n471), .B2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT64), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n473), .A2(new_n474), .A3(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n470), .B1(new_n476), .B2(G101), .ZN(new_n477));
  INV_X1    g052(.A(G101), .ZN(new_n478));
  AOI211_X1 g053(.A(KEYINPUT65), .B(new_n478), .C1(new_n472), .C2(new_n475), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n467), .B(new_n469), .C1(new_n477), .C2(new_n479), .ZN(new_n480));
  INV_X1    g055(.A(new_n480), .ZN(G160));
  OAI21_X1  g056(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n482));
  INV_X1    g057(.A(G112), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n482), .B1(new_n483), .B2(G2105), .ZN(new_n484));
  AOI21_X1  g059(.A(new_n484), .B1(new_n468), .B2(G136), .ZN(new_n485));
  XNOR2_X1  g060(.A(KEYINPUT3), .B(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT66), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n486), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G124), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n485), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  XNOR2_X1  g068(.A(new_n493), .B(KEYINPUT67), .ZN(G162));
  AND2_X1   g069(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n495));
  OAI211_X1 g070(.A(G138), .B(new_n474), .C1(new_n495), .C2(new_n462), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n486), .A2(KEYINPUT4), .A3(G138), .A4(new_n474), .ZN(new_n499));
  NAND3_X1  g074(.A1(new_n486), .A2(G126), .A3(G2105), .ZN(new_n500));
  OAI21_X1  g075(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(G114), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n503), .A2(KEYINPUT68), .A3(G2105), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n503), .B2(G2105), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n502), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND4_X1  g081(.A1(new_n498), .A2(new_n499), .A3(new_n500), .A4(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(G164));
  INV_X1    g083(.A(G62), .ZN(new_n509));
  OR2_X1    g084(.A1(KEYINPUT5), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT5), .A2(G543), .ZN(new_n511));
  AOI21_X1  g086(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g087(.A1(G75), .A2(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT71), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g090(.A1(new_n515), .A2(G75), .A3(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(G651), .B1(new_n512), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(KEYINPUT72), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT72), .ZN(new_n520));
  OAI211_X1 g095(.A(new_n520), .B(G651), .C1(new_n512), .C2(new_n517), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT69), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(KEYINPUT69), .ZN(new_n526));
  OAI21_X1  g101(.A(G651), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G651), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n510), .A2(new_n511), .B1(KEYINPUT6), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n527), .A2(new_n529), .A3(KEYINPUT70), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT70), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(KEYINPUT69), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n523), .A2(KEYINPUT6), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n528), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n528), .A2(KEYINPUT6), .ZN(new_n535));
  AND2_X1   g110(.A1(KEYINPUT5), .A2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(KEYINPUT5), .A2(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(new_n535), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  OAI21_X1  g113(.A(new_n531), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n530), .A2(new_n539), .A3(G88), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  AOI21_X1  g116(.A(new_n541), .B1(KEYINPUT6), .B2(new_n528), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n534), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G50), .ZN(new_n545));
  NAND3_X1  g120(.A1(new_n522), .A2(new_n540), .A3(new_n545), .ZN(G303));
  INV_X1    g121(.A(G303), .ZN(G166));
  NAND3_X1  g122(.A1(new_n527), .A2(G51), .A3(new_n542), .ZN(new_n548));
  NAND3_X1  g123(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n549), .B(KEYINPUT7), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n510), .A2(new_n511), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT73), .ZN(new_n552));
  AND2_X1   g127(.A1(G63), .A2(G651), .ZN(new_n553));
  NAND3_X1  g128(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g130(.A(new_n552), .B1(new_n551), .B2(new_n553), .ZN(new_n556));
  OAI211_X1 g131(.A(new_n548), .B(new_n550), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  AND2_X1   g132(.A1(new_n530), .A2(new_n539), .ZN(new_n558));
  AOI21_X1  g133(.A(new_n557), .B1(G89), .B2(new_n558), .ZN(G168));
  NAND2_X1  g134(.A1(G77), .A2(G543), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n536), .A2(new_n537), .ZN(new_n561));
  INV_X1    g136(.A(G64), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n560), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n544), .A2(G52), .B1(new_n563), .B2(G651), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n530), .A2(new_n539), .A3(G90), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(G301));
  INV_X1    g141(.A(G301), .ZN(G171));
  AOI22_X1  g142(.A1(new_n551), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n568));
  OR2_X1    g143(.A1(new_n568), .A2(new_n528), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n530), .A2(new_n539), .A3(G81), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n544), .A2(G43), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n570), .A2(KEYINPUT74), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT74), .B1(new_n570), .B2(new_n571), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n569), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(G860), .ZN(G153));
  NAND4_X1  g151(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g152(.A1(G1), .A2(G3), .ZN(new_n578));
  XNOR2_X1  g153(.A(new_n578), .B(KEYINPUT8), .ZN(new_n579));
  NAND4_X1  g154(.A1(G319), .A2(G483), .A3(G661), .A4(new_n579), .ZN(G188));
  INV_X1    g155(.A(KEYINPUT9), .ZN(new_n581));
  AOI21_X1  g156(.A(new_n581), .B1(new_n544), .B2(G53), .ZN(new_n582));
  NAND4_X1  g157(.A1(new_n527), .A2(new_n581), .A3(G53), .A4(new_n542), .ZN(new_n583));
  INV_X1    g158(.A(new_n583), .ZN(new_n584));
  OAI21_X1  g159(.A(KEYINPUT75), .B1(new_n582), .B2(new_n584), .ZN(new_n585));
  XNOR2_X1  g160(.A(KEYINPUT69), .B(KEYINPUT6), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n542), .B1(new_n586), .B2(new_n528), .ZN(new_n587));
  INV_X1    g162(.A(G53), .ZN(new_n588));
  OAI21_X1  g163(.A(KEYINPUT9), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT75), .ZN(new_n590));
  NAND3_X1  g165(.A1(new_n589), .A2(new_n590), .A3(new_n583), .ZN(new_n591));
  NAND2_X1  g166(.A1(G78), .A2(G543), .ZN(new_n592));
  XOR2_X1   g167(.A(KEYINPUT76), .B(G65), .Z(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n593), .B2(new_n561), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(G651), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n530), .A2(new_n539), .A3(G91), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n585), .A2(new_n591), .A3(new_n595), .A4(new_n596), .ZN(G299));
  INV_X1    g172(.A(new_n557), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n530), .A2(new_n539), .A3(G89), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n598), .A2(new_n599), .ZN(G286));
  NAND3_X1  g175(.A1(new_n530), .A2(new_n539), .A3(G87), .ZN(new_n601));
  INV_X1    g176(.A(G74), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n528), .B1(new_n561), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g178(.A(new_n603), .B1(new_n544), .B2(G49), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n601), .A2(new_n604), .ZN(G288));
  NAND3_X1  g180(.A1(new_n544), .A2(KEYINPUT77), .A3(G48), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT77), .ZN(new_n607));
  INV_X1    g182(.A(G48), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n587), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n606), .A2(new_n609), .ZN(new_n610));
  NAND3_X1  g185(.A1(new_n530), .A2(new_n539), .A3(G86), .ZN(new_n611));
  NAND2_X1  g186(.A1(G73), .A2(G543), .ZN(new_n612));
  INV_X1    g187(.A(G61), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n561), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n614), .A2(G651), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n610), .A2(new_n611), .A3(new_n615), .ZN(G305));
  NAND2_X1  g191(.A1(new_n558), .A2(G85), .ZN(new_n617));
  NAND2_X1  g192(.A1(G72), .A2(G543), .ZN(new_n618));
  INV_X1    g193(.A(G60), .ZN(new_n619));
  OAI21_X1  g194(.A(new_n618), .B1(new_n561), .B2(new_n619), .ZN(new_n620));
  AOI22_X1  g195(.A1(new_n544), .A2(G47), .B1(new_n620), .B2(G651), .ZN(new_n621));
  NAND2_X1  g196(.A1(new_n617), .A2(new_n621), .ZN(G290));
  NAND2_X1  g197(.A1(G301), .A2(G868), .ZN(new_n623));
  NAND2_X1  g198(.A1(G79), .A2(G543), .ZN(new_n624));
  INV_X1    g199(.A(G66), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n561), .B2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n626), .A2(G651), .ZN(new_n627));
  INV_X1    g202(.A(G54), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(new_n587), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n530), .A2(new_n539), .A3(G92), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND4_X1  g207(.A1(new_n530), .A2(new_n539), .A3(KEYINPUT10), .A4(G92), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n629), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n623), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n623), .B1(new_n634), .B2(G868), .ZN(G321));
  NAND2_X1  g211(.A1(G286), .A2(G868), .ZN(new_n637));
  INV_X1    g212(.A(G299), .ZN(new_n638));
  OAI21_X1  g213(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G297));
  OAI21_X1  g214(.A(new_n637), .B1(new_n638), .B2(G868), .ZN(G280));
  INV_X1    g215(.A(G559), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n634), .B1(new_n641), .B2(G860), .ZN(G148));
  INV_X1    g217(.A(G868), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n574), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g219(.A1(new_n632), .A2(new_n633), .ZN(new_n645));
  INV_X1    g220(.A(new_n629), .ZN(new_n646));
  NAND2_X1  g221(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n647), .A2(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(new_n643), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g225(.A1(new_n476), .A2(new_n486), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT12), .Z(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT13), .Z(new_n653));
  INV_X1    g228(.A(G2100), .ZN(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  OAI21_X1  g231(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n657));
  INV_X1    g232(.A(G111), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n657), .B1(new_n658), .B2(G2105), .ZN(new_n659));
  NAND2_X1  g234(.A1(new_n468), .A2(G135), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  AND2_X1   g236(.A1(new_n489), .A2(new_n490), .ZN(new_n662));
  AOI211_X1 g237(.A(new_n659), .B(new_n661), .C1(new_n662), .C2(G123), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(G2096), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n655), .A2(new_n656), .A3(new_n664), .ZN(G156));
  XOR2_X1   g240(.A(G1341), .B(G1348), .Z(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT78), .ZN(new_n667));
  XOR2_X1   g242(.A(G2451), .B(G2454), .Z(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT16), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n667), .B(new_n669), .ZN(new_n670));
  INV_X1    g245(.A(KEYINPUT14), .ZN(new_n671));
  XNOR2_X1  g246(.A(G2427), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2430), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT15), .B(G2435), .ZN(new_n674));
  AOI21_X1  g249(.A(new_n671), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  OAI21_X1  g250(.A(new_n675), .B1(new_n674), .B2(new_n673), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n670), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(G2443), .B(G2446), .ZN(new_n679));
  OR2_X1    g254(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g255(.A1(new_n678), .A2(new_n679), .ZN(new_n681));
  AND3_X1   g256(.A1(new_n680), .A2(G14), .A3(new_n681), .ZN(G401));
  XOR2_X1   g257(.A(G2084), .B(G2090), .Z(new_n683));
  XNOR2_X1  g258(.A(G2067), .B(G2678), .ZN(new_n684));
  XNOR2_X1  g259(.A(G2072), .B(G2078), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT18), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT79), .B(KEYINPUT17), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n685), .B(new_n688), .ZN(new_n689));
  INV_X1    g264(.A(new_n684), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(new_n684), .A2(new_n685), .ZN(new_n692));
  NOR3_X1   g267(.A1(new_n691), .A2(new_n683), .A3(new_n692), .ZN(new_n693));
  AND2_X1   g268(.A1(new_n690), .A2(new_n683), .ZN(new_n694));
  AOI211_X1 g269(.A(new_n687), .B(new_n693), .C1(new_n689), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(G2096), .ZN(new_n696));
  XNOR2_X1  g271(.A(KEYINPUT80), .B(G2100), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(G227));
  XOR2_X1   g273(.A(G1971), .B(G1976), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT19), .ZN(new_n700));
  XOR2_X1   g275(.A(G1956), .B(G2474), .Z(new_n701));
  XOR2_X1   g276(.A(G1961), .B(G1966), .Z(new_n702));
  AND2_X1   g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(KEYINPUT20), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n704), .B(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n701), .A2(new_n702), .ZN(new_n707));
  NOR2_X1   g282(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  MUX2_X1   g283(.A(new_n708), .B(new_n707), .S(new_n700), .Z(new_n709));
  NOR2_X1   g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1991), .B(G1996), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(G1981), .B(G1986), .ZN(new_n715));
  XNOR2_X1  g290(.A(new_n714), .B(new_n715), .ZN(G229));
  NAND2_X1  g291(.A1(G162), .A2(G29), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT29), .ZN(new_n718));
  OR2_X1    g293(.A1(G29), .A2(G35), .ZN(new_n719));
  AND3_X1   g294(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n718), .B1(new_n717), .B2(new_n719), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  INV_X1    g297(.A(G2090), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n722), .A2(KEYINPUT95), .A3(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n720), .B2(new_n721), .ZN(new_n725));
  INV_X1    g300(.A(KEYINPUT95), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G4), .A2(G16), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n634), .B2(G16), .ZN(new_n729));
  OR2_X1    g304(.A1(new_n729), .A2(G1348), .ZN(new_n730));
  INV_X1    g305(.A(G16), .ZN(new_n731));
  AND2_X1   g306(.A1(new_n731), .A2(G21), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G286), .B2(G16), .ZN(new_n733));
  INV_X1    g308(.A(G1966), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OR2_X1    g310(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(KEYINPUT94), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n736), .A2(new_n737), .B1(G1348), .B2(new_n729), .ZN(new_n738));
  NAND4_X1  g313(.A1(new_n724), .A2(new_n727), .A3(new_n730), .A4(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(KEYINPUT88), .B(KEYINPUT24), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AOI21_X1  g316(.A(G29), .B1(new_n741), .B2(G34), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G34), .B2(new_n741), .ZN(new_n743));
  INV_X1    g318(.A(G29), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n743), .B1(G160), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G2084), .ZN(new_n746));
  AND2_X1   g321(.A1(new_n744), .A2(G33), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT87), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n749), .B(KEYINPUT25), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n468), .A2(G139), .ZN(new_n751));
  AOI22_X1  g326(.A1(new_n486), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n750), .B(new_n751), .C1(new_n474), .C2(new_n752), .ZN(new_n753));
  AOI21_X1  g328(.A(new_n747), .B1(new_n753), .B2(G29), .ZN(new_n754));
  INV_X1    g329(.A(G2072), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT31), .B(G11), .Z(new_n757));
  INV_X1    g332(.A(KEYINPUT30), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n758), .A2(G28), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n744), .B1(new_n758), .B2(G28), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n761));
  OAI21_X1  g336(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  AOI211_X1 g338(.A(new_n757), .B(new_n763), .C1(new_n663), .C2(G29), .ZN(new_n764));
  NOR2_X1   g339(.A1(G27), .A2(G29), .ZN(new_n765));
  AOI21_X1  g340(.A(new_n765), .B1(G164), .B2(G29), .ZN(new_n766));
  INV_X1    g341(.A(G2078), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n756), .A2(new_n764), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT89), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n770), .B1(new_n754), .B2(new_n755), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n753), .A2(G29), .ZN(new_n772));
  OAI211_X1 g347(.A(KEYINPUT89), .B(G2072), .C1(new_n772), .C2(new_n747), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n746), .B(new_n769), .C1(new_n771), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(KEYINPUT27), .B(G1996), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n662), .A2(G129), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT90), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT26), .ZN(new_n779));
  AND2_X1   g354(.A1(new_n476), .A2(G105), .ZN(new_n780));
  AOI211_X1 g355(.A(new_n779), .B(new_n780), .C1(G141), .C2(new_n468), .ZN(new_n781));
  NAND4_X1  g356(.A1(new_n777), .A2(KEYINPUT91), .A3(G29), .A4(new_n781), .ZN(new_n782));
  AND3_X1   g357(.A1(new_n777), .A2(G29), .A3(new_n781), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT91), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n784), .B1(G29), .B2(G32), .ZN(new_n785));
  OAI211_X1 g360(.A(new_n775), .B(new_n782), .C1(new_n783), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n744), .A2(G26), .ZN(new_n787));
  XOR2_X1   g362(.A(new_n787), .B(KEYINPUT28), .Z(new_n788));
  NAND2_X1  g363(.A1(new_n468), .A2(G140), .ZN(new_n789));
  NOR2_X1   g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT86), .Z(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(new_n474), .B2(G116), .ZN(new_n792));
  INV_X1    g367(.A(G128), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n789), .B1(new_n791), .B2(new_n792), .C1(new_n491), .C2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n788), .B1(new_n794), .B2(G29), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(G2067), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n731), .A2(G5), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(G171), .B2(new_n731), .ZN(new_n798));
  INV_X1    g373(.A(G1961), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n798), .B(new_n799), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n786), .A2(new_n796), .A3(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n782), .B1(new_n783), .B2(new_n785), .ZN(new_n802));
  INV_X1    g377(.A(new_n775), .ZN(new_n803));
  INV_X1    g378(.A(KEYINPUT92), .ZN(new_n804));
  OR3_X1    g379(.A1(new_n733), .A2(new_n804), .A3(new_n734), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n804), .B1(new_n733), .B2(new_n734), .ZN(new_n806));
  AOI22_X1  g381(.A1(new_n802), .A2(new_n803), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  XNOR2_X1  g382(.A(KEYINPUT81), .B(G16), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(G20), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT23), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n638), .B2(new_n731), .ZN(new_n811));
  INV_X1    g386(.A(G1956), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n774), .A2(new_n801), .A3(new_n807), .A4(new_n813), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n808), .A2(G19), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(new_n575), .B2(new_n808), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1341), .Z(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n722), .B2(new_n723), .ZN(new_n818));
  NOR3_X1   g393(.A1(new_n739), .A2(new_n814), .A3(new_n818), .ZN(new_n819));
  MUX2_X1   g394(.A(G6), .B(G305), .S(G16), .Z(new_n820));
  XOR2_X1   g395(.A(KEYINPUT32), .B(G1981), .Z(new_n821));
  XNOR2_X1  g396(.A(new_n821), .B(KEYINPUT82), .ZN(new_n822));
  XNOR2_X1  g397(.A(new_n820), .B(new_n822), .ZN(new_n823));
  INV_X1    g398(.A(new_n808), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n824), .A2(G22), .ZN(new_n825));
  AOI21_X1  g400(.A(new_n825), .B1(G166), .B2(new_n824), .ZN(new_n826));
  INV_X1    g401(.A(G1971), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(KEYINPUT83), .B1(new_n601), .B2(new_n604), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n601), .A2(new_n604), .A3(KEYINPUT83), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n830), .A2(G16), .A3(new_n831), .ZN(new_n832));
  OAI21_X1  g407(.A(new_n832), .B1(G16), .B2(G23), .ZN(new_n833));
  XOR2_X1   g408(.A(KEYINPUT33), .B(G1976), .Z(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT84), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n833), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n833), .A2(new_n835), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n823), .A2(new_n828), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT34), .ZN(new_n839));
  INV_X1    g414(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n744), .A2(G25), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n662), .A2(G119), .ZN(new_n842));
  OAI21_X1  g417(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n843));
  INV_X1    g418(.A(G107), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n845), .B1(new_n468), .B2(G131), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(new_n847), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n841), .B1(new_n848), .B2(new_n744), .ZN(new_n849));
  XOR2_X1   g424(.A(KEYINPUT35), .B(G1991), .Z(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  NOR2_X1   g426(.A1(new_n824), .A2(G24), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n617), .A2(new_n621), .ZN(new_n853));
  AOI21_X1  g428(.A(new_n852), .B1(new_n853), .B2(new_n824), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(G1986), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n851), .A2(new_n855), .ZN(new_n856));
  OAI21_X1  g431(.A(new_n856), .B1(new_n838), .B2(KEYINPUT34), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT36), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT85), .ZN(new_n859));
  OR3_X1    g434(.A1(new_n840), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n858), .A2(KEYINPUT85), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n859), .B(new_n861), .C1(new_n840), .C2(new_n857), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n819), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(G311));
  INV_X1    g439(.A(KEYINPUT96), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n863), .B(new_n865), .ZN(G150));
  NAND2_X1  g441(.A1(G80), .A2(G543), .ZN(new_n867));
  INV_X1    g442(.A(G67), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n867), .B1(new_n561), .B2(new_n868), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n544), .A2(G55), .B1(new_n869), .B2(G651), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n530), .A2(new_n539), .A3(G93), .ZN(new_n871));
  AND2_X1   g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(G860), .ZN(new_n873));
  NOR2_X1   g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n874), .B(KEYINPUT37), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n634), .A2(G559), .ZN(new_n876));
  XOR2_X1   g451(.A(KEYINPUT97), .B(KEYINPUT38), .Z(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT98), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n876), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(new_n872), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n574), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g456(.A(new_n569), .B(new_n872), .C1(new_n572), .C2(new_n573), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n879), .B(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(new_n884), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n885), .A2(KEYINPUT39), .ZN(new_n886));
  OAI21_X1  g461(.A(new_n873), .B1(new_n885), .B2(KEYINPUT39), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n875), .B1(new_n886), .B2(new_n887), .ZN(G145));
  INV_X1    g463(.A(G37), .ZN(new_n889));
  OAI21_X1  g464(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n890));
  INV_X1    g465(.A(G118), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n890), .B1(new_n891), .B2(G2105), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n892), .B1(new_n468), .B2(G142), .ZN(new_n893));
  INV_X1    g468(.A(G130), .ZN(new_n894));
  OAI21_X1  g469(.A(new_n893), .B1(new_n491), .B2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n652), .B(new_n895), .ZN(new_n896));
  XNOR2_X1  g471(.A(new_n896), .B(new_n847), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT99), .ZN(new_n898));
  OR2_X1    g473(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n897), .A2(new_n898), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n777), .A2(new_n781), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n794), .B(G164), .ZN(new_n902));
  OR2_X1    g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NOR2_X1   g480(.A1(new_n905), .A2(new_n753), .ZN(new_n906));
  INV_X1    g481(.A(new_n753), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n907), .B1(new_n903), .B2(new_n904), .ZN(new_n908));
  OAI211_X1 g483(.A(new_n899), .B(new_n900), .C1(new_n906), .C2(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n663), .B(G160), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n910), .B(G162), .ZN(new_n911));
  INV_X1    g486(.A(new_n906), .ZN(new_n912));
  INV_X1    g487(.A(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g489(.A(new_n909), .B(new_n911), .C1(new_n914), .C2(new_n897), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n899), .A2(new_n900), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n912), .A2(new_n913), .A3(new_n916), .ZN(new_n917));
  AND2_X1   g492(.A1(new_n917), .A2(new_n909), .ZN(new_n918));
  OAI211_X1 g493(.A(new_n889), .B(new_n915), .C1(new_n918), .C2(new_n911), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n919), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g495(.A1(new_n570), .A2(new_n571), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT74), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n570), .A2(KEYINPUT74), .A3(new_n571), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n872), .B1(new_n925), .B2(new_n569), .ZN(new_n926));
  INV_X1    g501(.A(new_n882), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n648), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  OAI211_X1 g503(.A(new_n881), .B(new_n882), .C1(G559), .C2(new_n647), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n647), .A2(G299), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n596), .A2(new_n595), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n590), .B1(new_n589), .B2(new_n583), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n634), .A2(new_n934), .A3(new_n591), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n931), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n930), .A2(new_n936), .ZN(new_n937));
  AND3_X1   g512(.A1(new_n931), .A2(KEYINPUT41), .A3(new_n935), .ZN(new_n938));
  AOI21_X1  g513(.A(KEYINPUT41), .B1(new_n931), .B2(new_n935), .ZN(new_n939));
  NOR2_X1   g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  OAI211_X1 g516(.A(new_n937), .B(KEYINPUT100), .C1(new_n930), .C2(new_n941), .ZN(new_n942));
  INV_X1    g517(.A(KEYINPUT100), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n930), .A2(new_n943), .A3(new_n936), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n945), .A2(KEYINPUT42), .ZN(new_n946));
  INV_X1    g521(.A(new_n831), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n853), .B1(new_n947), .B2(new_n829), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n830), .A2(G290), .A3(new_n831), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  AND2_X1   g525(.A1(new_n540), .A2(new_n545), .ZN(new_n951));
  NAND3_X1  g526(.A1(G305), .A2(new_n951), .A3(new_n522), .ZN(new_n952));
  AOI22_X1  g527(.A1(new_n606), .A2(new_n609), .B1(G651), .B2(new_n614), .ZN(new_n953));
  NAND3_X1  g528(.A1(G303), .A2(new_n611), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  NAND4_X1  g531(.A1(new_n948), .A2(new_n949), .A3(new_n954), .A4(new_n952), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT42), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n942), .A2(new_n960), .A3(new_n944), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n946), .A2(new_n959), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n959), .B1(new_n946), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(G868), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n880), .A2(new_n643), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(G295));
  NAND2_X1  g541(.A1(new_n964), .A2(new_n965), .ZN(G331));
  NAND2_X1  g542(.A1(G301), .A2(KEYINPUT101), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n564), .A2(new_n565), .A3(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(G286), .A3(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(G168), .A2(new_n969), .A3(G171), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(new_n973), .B1(new_n926), .B2(new_n927), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n881), .A2(new_n882), .A3(new_n972), .A4(new_n971), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n936), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT102), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n974), .A2(new_n975), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n979), .A2(new_n940), .ZN(new_n980));
  NAND4_X1  g555(.A1(new_n974), .A2(new_n975), .A3(KEYINPUT102), .A4(new_n936), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n959), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n956), .A2(new_n957), .A3(KEYINPUT103), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT103), .B1(new_n956), .B2(new_n957), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AOI21_X1  g562(.A(G37), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  INV_X1    g563(.A(KEYINPUT104), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n983), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT103), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n958), .A2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n984), .ZN(new_n993));
  AOI22_X1  g568(.A1(new_n977), .A2(new_n976), .B1(new_n979), .B2(new_n940), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n993), .B1(new_n994), .B2(new_n981), .ZN(new_n995));
  OAI21_X1  g570(.A(KEYINPUT104), .B1(new_n995), .B2(G37), .ZN(new_n996));
  AOI21_X1  g571(.A(KEYINPUT43), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  OR2_X1    g572(.A1(new_n980), .A2(KEYINPUT105), .ZN(new_n998));
  INV_X1    g573(.A(new_n976), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n999), .B1(new_n980), .B2(KEYINPUT105), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n993), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n889), .B1(new_n982), .B2(new_n959), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  OAI21_X1  g579(.A(KEYINPUT44), .B1(new_n997), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n1003), .B1(new_n990), .B2(new_n996), .ZN(new_n1007));
  NOR3_X1   g582(.A1(new_n1001), .A2(new_n1002), .A3(KEYINPUT43), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1005), .A2(new_n1009), .ZN(G397));
  INV_X1    g585(.A(G1384), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n507), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT45), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n473), .B1(G2104), .B2(new_n474), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n471), .A2(KEYINPUT64), .A3(G2105), .ZN(new_n1016));
  OAI21_X1  g591(.A(G101), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1017), .A2(KEYINPUT65), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n476), .A2(new_n470), .A3(G101), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  NAND4_X1  g595(.A1(new_n1020), .A2(G40), .A3(new_n467), .A4(new_n469), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1014), .A2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g597(.A(new_n1022), .B(KEYINPUT106), .ZN(new_n1023));
  INV_X1    g598(.A(G1996), .ZN(new_n1024));
  XNOR2_X1  g599(.A(new_n901), .B(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(G2067), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n794), .B(new_n1026), .ZN(new_n1027));
  AND2_X1   g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n848), .A2(new_n850), .ZN(new_n1029));
  OR2_X1    g604(.A1(new_n848), .A2(new_n850), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .ZN(new_n1031));
  XNOR2_X1  g606(.A(G290), .B(G1986), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1023), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G40), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n480), .A2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1035), .A2(new_n1014), .A3(KEYINPUT112), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  AOI21_X1  g612(.A(KEYINPUT45), .B1(new_n507), .B2(new_n1011), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1037), .B1(new_n1021), .B2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1041), .A2(new_n734), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1012), .A2(KEYINPUT50), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT50), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n507), .A2(new_n1044), .A3(new_n1011), .ZN(new_n1045));
  XNOR2_X1  g620(.A(KEYINPUT113), .B(G2084), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1035), .A2(new_n1043), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1021), .B1(KEYINPUT50), .B2(new_n1012), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n1050), .A2(KEYINPUT114), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1042), .A2(G168), .A3(new_n1049), .A4(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1052), .A2(G8), .ZN(new_n1053));
  AND2_X1   g628(.A1(new_n1051), .A2(new_n1049), .ZN(new_n1054));
  AOI21_X1  g629(.A(G168), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT51), .B1(new_n1053), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT51), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n1052), .A2(new_n1057), .A3(G8), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1056), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT62), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT62), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1056), .A2(new_n1061), .A3(new_n1058), .ZN(new_n1062));
  INV_X1    g637(.A(G8), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1035), .A2(new_n1014), .A3(new_n1040), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1064), .A2(new_n827), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1035), .A2(new_n1043), .A3(new_n723), .A4(new_n1045), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1063), .B1(new_n1067), .B2(KEYINPUT107), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1063), .B1(new_n951), .B2(new_n522), .ZN(new_n1069));
  AOI21_X1  g644(.A(KEYINPUT108), .B1(new_n1069), .B2(KEYINPUT55), .ZN(new_n1070));
  NAND4_X1  g645(.A1(G303), .A2(KEYINPUT108), .A3(KEYINPUT55), .A4(G8), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(G303), .A2(G8), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT55), .ZN(new_n1074));
  AOI21_X1  g649(.A(KEYINPUT109), .B1(new_n1073), .B2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT109), .ZN(new_n1076));
  AOI211_X1 g651(.A(new_n1076), .B(KEYINPUT55), .C1(G303), .C2(G8), .ZN(new_n1077));
  OAI22_X1  g652(.A1(new_n1070), .A2(new_n1072), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT107), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1065), .A2(new_n1079), .A3(new_n1066), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1068), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT49), .ZN(new_n1082));
  NOR2_X1   g657(.A1(G305), .A2(G1981), .ZN(new_n1083));
  INV_X1    g658(.A(G1981), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n953), .B2(new_n611), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1082), .B1(new_n1083), .B2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(G305), .A2(G1981), .ZN(new_n1087));
  NAND3_X1  g662(.A1(new_n953), .A2(new_n1084), .A3(new_n611), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1087), .A2(KEYINPUT49), .A3(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1012), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1063), .B1(new_n1035), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1086), .A2(new_n1089), .A3(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n830), .A2(G1976), .A3(new_n831), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(new_n1091), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT52), .ZN(new_n1095));
  INV_X1    g670(.A(G1976), .ZN(new_n1096));
  AOI21_X1  g671(.A(KEYINPUT52), .B1(G288), .B2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1093), .A2(new_n1091), .A3(new_n1097), .ZN(new_n1098));
  AND3_X1   g673(.A1(new_n1092), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1076), .B1(new_n1069), .B2(KEYINPUT55), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1073), .A2(KEYINPUT109), .A3(new_n1074), .ZN(new_n1101));
  NAND3_X1  g676(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT108), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  AOI22_X1  g679(.A1(new_n1100), .A2(new_n1101), .B1(new_n1104), .B2(new_n1071), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n507), .A2(KEYINPUT45), .A3(new_n1011), .ZN(new_n1106));
  NOR3_X1   g681(.A1(new_n1106), .A2(new_n1021), .A3(new_n1038), .ZN(new_n1107));
  OAI211_X1 g682(.A(KEYINPUT111), .B(new_n1066), .C1(new_n1107), .C2(G1971), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1108), .A2(G8), .ZN(new_n1109));
  AOI21_X1  g684(.A(KEYINPUT111), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1081), .A2(new_n1099), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  NOR2_X1   g688(.A1(new_n1113), .A2(G2078), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .A4(new_n1114), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1035), .A2(new_n1014), .A3(new_n767), .A4(new_n1040), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1116), .A2(new_n1113), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1035), .A2(new_n1043), .A3(new_n1045), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1118), .A2(new_n799), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1120), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1121));
  AOI21_X1  g696(.A(KEYINPUT122), .B1(new_n1120), .B2(G171), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1112), .B1(new_n1121), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1060), .A2(new_n1062), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT119), .B1(G299), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n934), .A2(new_n1128), .A3(KEYINPUT57), .A4(new_n591), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(KEYINPUT117), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n932), .A2(new_n1131), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n596), .A2(KEYINPUT117), .A3(new_n595), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT116), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n582), .B2(new_n584), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n589), .A2(KEYINPUT116), .A3(new_n583), .ZN(new_n1136));
  NAND4_X1  g711(.A1(new_n1132), .A2(new_n1133), .A3(new_n1135), .A4(new_n1136), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1137), .A2(KEYINPUT118), .A3(new_n1126), .ZN(new_n1138));
  AOI21_X1  g713(.A(KEYINPUT118), .B1(new_n1137), .B2(new_n1126), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1130), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(KEYINPUT56), .B(G2072), .ZN(new_n1141));
  AOI22_X1  g716(.A1(new_n1107), .A2(new_n1141), .B1(new_n1118), .B2(new_n812), .ZN(new_n1142));
  AOI21_X1  g717(.A(KEYINPUT120), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(new_n1143), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1140), .A2(KEYINPUT120), .A3(new_n1142), .ZN(new_n1145));
  INV_X1    g720(.A(G1348), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1118), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1147), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT121), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1035), .A2(new_n1149), .A3(new_n1090), .ZN(new_n1150));
  OAI21_X1  g725(.A(KEYINPUT121), .B1(new_n1021), .B2(new_n1012), .ZN(new_n1151));
  AOI21_X1  g726(.A(G2067), .B1(new_n1150), .B2(new_n1151), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n634), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1142), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1154), .B(new_n1130), .C1(new_n1139), .C2(new_n1138), .ZN(new_n1155));
  AOI22_X1  g730(.A1(new_n1144), .A2(new_n1145), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  AND3_X1   g731(.A1(new_n1140), .A2(KEYINPUT120), .A3(new_n1142), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1155), .B1(new_n1157), .B2(new_n1143), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT61), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1161));
  AND3_X1   g736(.A1(new_n1161), .A2(KEYINPUT61), .A3(new_n1155), .ZN(new_n1162));
  INV_X1    g737(.A(new_n1152), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n1147), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT60), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1148), .B2(new_n1152), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n634), .A3(new_n1166), .ZN(new_n1167));
  NAND4_X1  g742(.A1(new_n1163), .A2(KEYINPUT60), .A3(new_n647), .A4(new_n1147), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1107), .A2(new_n1024), .ZN(new_n1169));
  XOR2_X1   g744(.A(KEYINPUT58), .B(G1341), .Z(new_n1170));
  NAND3_X1  g745(.A1(new_n1150), .A2(new_n1151), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n574), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g749(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1175));
  OAI211_X1 g750(.A(new_n1167), .B(new_n1168), .C1(new_n1174), .C2(new_n1175), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1162), .A2(new_n1176), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1156), .B1(new_n1160), .B2(new_n1177), .ZN(new_n1178));
  AND3_X1   g753(.A1(new_n1120), .A2(KEYINPUT122), .A3(G171), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n469), .B(new_n1180), .C1(new_n477), .C2(new_n479), .ZN(new_n1181));
  NOR3_X1   g756(.A1(new_n1113), .A2(new_n1034), .A3(G2078), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n467), .A3(new_n1182), .ZN(new_n1183));
  AOI21_X1  g758(.A(new_n1180), .B1(new_n1020), .B2(new_n469), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n1106), .A2(new_n1038), .ZN(new_n1186));
  AOI22_X1  g761(.A1(new_n1116), .A2(new_n1113), .B1(new_n1185), .B2(new_n1186), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT123), .ZN(new_n1188));
  AND3_X1   g763(.A1(new_n1118), .A2(new_n1188), .A3(new_n799), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1188), .B1(new_n1118), .B2(new_n799), .ZN(new_n1190));
  OAI211_X1 g765(.A(new_n1187), .B(G301), .C1(new_n1189), .C2(new_n1190), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1191), .ZN(new_n1192));
  NOR3_X1   g767(.A1(new_n1179), .A2(new_n1192), .A3(new_n1122), .ZN(new_n1193));
  OAI21_X1  g768(.A(KEYINPUT125), .B1(new_n1193), .B2(KEYINPUT54), .ZN(new_n1194));
  NAND3_X1  g769(.A1(new_n1123), .A2(new_n1121), .A3(new_n1191), .ZN(new_n1195));
  INV_X1    g770(.A(KEYINPUT125), .ZN(new_n1196));
  INV_X1    g771(.A(KEYINPUT54), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .ZN(new_n1198));
  NAND2_X1  g773(.A1(new_n1119), .A2(KEYINPUT123), .ZN(new_n1199));
  NAND3_X1  g774(.A1(new_n1118), .A2(new_n1188), .A3(new_n799), .ZN(new_n1200));
  NAND2_X1  g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  AOI21_X1  g776(.A(G301), .B1(new_n1201), .B2(new_n1187), .ZN(new_n1202));
  NOR2_X1   g777(.A1(new_n1120), .A2(G171), .ZN(new_n1203));
  NOR3_X1   g778(.A1(new_n1202), .A2(new_n1197), .A3(new_n1203), .ZN(new_n1204));
  NOR2_X1   g779(.A1(new_n1204), .A2(new_n1112), .ZN(new_n1205));
  NAND4_X1  g780(.A1(new_n1194), .A2(new_n1198), .A3(new_n1059), .A4(new_n1205), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1125), .B1(new_n1178), .B2(new_n1206), .ZN(new_n1207));
  INV_X1    g782(.A(KEYINPUT115), .ZN(new_n1208));
  INV_X1    g783(.A(KEYINPUT63), .ZN(new_n1209));
  NAND2_X1  g784(.A1(G168), .A2(G8), .ZN(new_n1210));
  AOI21_X1  g785(.A(new_n1210), .B1(new_n1054), .B2(new_n1042), .ZN(new_n1211));
  NAND4_X1  g786(.A1(new_n1081), .A2(new_n1099), .A3(new_n1211), .A4(new_n1111), .ZN(new_n1212));
  AOI21_X1  g787(.A(new_n1078), .B1(new_n1068), .B2(new_n1080), .ZN(new_n1213));
  INV_X1    g788(.A(new_n1210), .ZN(new_n1214));
  INV_X1    g789(.A(new_n1042), .ZN(new_n1215));
  NAND2_X1  g790(.A1(new_n1051), .A2(new_n1049), .ZN(new_n1216));
  OAI211_X1 g791(.A(KEYINPUT63), .B(new_n1214), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1213), .A2(new_n1217), .ZN(new_n1218));
  NAND3_X1  g793(.A1(new_n1092), .A2(new_n1095), .A3(new_n1098), .ZN(new_n1219));
  INV_X1    g794(.A(new_n1066), .ZN(new_n1220));
  NOR2_X1   g795(.A1(new_n1021), .A2(new_n1038), .ZN(new_n1221));
  AOI21_X1  g796(.A(G1971), .B1(new_n1221), .B2(new_n1040), .ZN(new_n1222));
  OAI21_X1  g797(.A(KEYINPUT107), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  AND3_X1   g798(.A1(new_n1223), .A2(G8), .A3(new_n1080), .ZN(new_n1224));
  AOI21_X1  g799(.A(new_n1219), .B1(new_n1224), .B2(new_n1078), .ZN(new_n1225));
  AOI22_X1  g800(.A1(new_n1209), .A2(new_n1212), .B1(new_n1218), .B2(new_n1225), .ZN(new_n1226));
  NOR2_X1   g801(.A1(G288), .A2(G1976), .ZN(new_n1227));
  AOI21_X1  g802(.A(new_n1083), .B1(new_n1092), .B2(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT110), .ZN(new_n1229));
  NAND2_X1  g804(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  INV_X1    g805(.A(new_n1230), .ZN(new_n1231));
  OAI21_X1  g806(.A(new_n1091), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1232));
  OAI22_X1  g807(.A1(new_n1231), .A2(new_n1232), .B1(new_n1081), .B2(new_n1219), .ZN(new_n1233));
  OAI21_X1  g808(.A(new_n1208), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g809(.A1(new_n1212), .A2(new_n1209), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1218), .A2(new_n1225), .ZN(new_n1236));
  NAND2_X1  g811(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g812(.A1(new_n1081), .A2(new_n1219), .ZN(new_n1238));
  INV_X1    g813(.A(new_n1232), .ZN(new_n1239));
  AOI21_X1  g814(.A(new_n1238), .B1(new_n1239), .B2(new_n1230), .ZN(new_n1240));
  NAND3_X1  g815(.A1(new_n1237), .A2(KEYINPUT115), .A3(new_n1240), .ZN(new_n1241));
  NAND2_X1  g816(.A1(new_n1234), .A2(new_n1241), .ZN(new_n1242));
  OAI21_X1  g817(.A(new_n1033), .B1(new_n1207), .B2(new_n1242), .ZN(new_n1243));
  NAND2_X1  g818(.A1(new_n1031), .A2(new_n1023), .ZN(new_n1244));
  INV_X1    g819(.A(G1986), .ZN(new_n1245));
  NAND3_X1  g820(.A1(new_n1023), .A2(new_n1245), .A3(new_n853), .ZN(new_n1246));
  INV_X1    g821(.A(KEYINPUT48), .ZN(new_n1247));
  NAND2_X1  g822(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1248));
  OR2_X1    g823(.A1(new_n1246), .A2(new_n1247), .ZN(new_n1249));
  NAND3_X1  g824(.A1(new_n1244), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  XOR2_X1   g825(.A(new_n1029), .B(KEYINPUT126), .Z(new_n1251));
  NAND2_X1  g826(.A1(new_n1028), .A2(new_n1251), .ZN(new_n1252));
  OAI21_X1  g827(.A(new_n1252), .B1(G2067), .B2(new_n794), .ZN(new_n1253));
  NAND2_X1  g828(.A1(new_n1253), .A2(new_n1023), .ZN(new_n1254));
  NAND2_X1  g829(.A1(new_n1250), .A2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g830(.A(KEYINPUT46), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1256));
  NAND3_X1  g831(.A1(new_n1023), .A2(KEYINPUT46), .A3(new_n1024), .ZN(new_n1257));
  XNOR2_X1  g832(.A(new_n1257), .B(KEYINPUT127), .ZN(new_n1258));
  NAND3_X1  g833(.A1(new_n1027), .A2(new_n777), .A3(new_n781), .ZN(new_n1259));
  AOI211_X1 g834(.A(new_n1256), .B(new_n1258), .C1(new_n1023), .C2(new_n1259), .ZN(new_n1260));
  INV_X1    g835(.A(KEYINPUT47), .ZN(new_n1261));
  OR2_X1    g836(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g837(.A1(new_n1260), .A2(new_n1261), .ZN(new_n1263));
  AOI21_X1  g838(.A(new_n1255), .B1(new_n1262), .B2(new_n1263), .ZN(new_n1264));
  NAND2_X1  g839(.A1(new_n1243), .A2(new_n1264), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g840(.A1(G229), .A2(new_n459), .A3(G401), .A4(G227), .ZN(new_n1267));
  OAI211_X1 g841(.A(new_n1267), .B(new_n919), .C1(new_n1007), .C2(new_n1008), .ZN(G225));
  INV_X1    g842(.A(G225), .ZN(G308));
endmodule


