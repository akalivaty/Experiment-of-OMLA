//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 0 1 0 1 0 1 0 1 0 1 1 1 1 1 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:39 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1262, new_n1263,
    new_n1264;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR3_X1   g0004(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n205));
  OAI211_X1 g0005(.A(new_n205), .B(G250), .C1(G257), .C2(G264), .ZN(new_n206));
  XOR2_X1   g0006(.A(new_n206), .B(KEYINPUT0), .Z(new_n207));
  AOI22_X1  g0007(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n208));
  INV_X1    g0008(.A(G116), .ZN(new_n209));
  INV_X1    g0009(.A(G270), .ZN(new_n210));
  OAI21_X1  g0010(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  INV_X1    g0014(.A(G97), .ZN(new_n215));
  INV_X1    g0015(.A(G257), .ZN(new_n216));
  OAI221_X1 g0016(.A(new_n212), .B1(new_n213), .B2(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  AOI211_X1 g0017(.A(new_n211), .B(new_n217), .C1(G58), .C2(G232), .ZN(new_n218));
  AOI21_X1  g0018(.A(new_n218), .B1(G1), .B2(G20), .ZN(new_n219));
  XOR2_X1   g0019(.A(new_n219), .B(KEYINPUT1), .Z(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n204), .ZN(new_n222));
  OAI21_X1  g0022(.A(G50), .B1(G58), .B2(G68), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  AOI211_X1 g0024(.A(new_n207), .B(new_n220), .C1(new_n222), .C2(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n226));
  XNOR2_X1  g0026(.A(G238), .B(G244), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G264), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(new_n210), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n230), .B(new_n233), .ZN(G358));
  XNOR2_X1  g0034(.A(G87), .B(G97), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT65), .ZN(new_n236));
  INV_X1    g0036(.A(G107), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n209), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G68), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G58), .ZN(new_n241));
  INV_X1    g0041(.A(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(new_n239), .B(new_n243), .Z(G351));
  OAI21_X1  g0044(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n245));
  INV_X1    g0045(.A(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G274), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n249), .A2(G226), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G97), .ZN(new_n252));
  AND2_X1   g0052(.A1(KEYINPUT3), .A2(G33), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT3), .A2(G33), .ZN(new_n254));
  OAI211_X1 g0054(.A(G232), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND3_X1  g0055(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  INV_X1    g0057(.A(G41), .ZN(new_n258));
  OAI211_X1 g0058(.A(G1), .B(G13), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  AOI21_X1  g0060(.A(new_n248), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT13), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n260), .A2(new_n246), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G238), .ZN(new_n264));
  AND3_X1   g0064(.A1(new_n261), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n262), .B1(new_n261), .B2(new_n264), .ZN(new_n266));
  OAI21_X1  g0066(.A(G169), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(KEYINPUT14), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n265), .A2(new_n266), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n269), .A2(G179), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT14), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n271), .B(G169), .C1(new_n265), .C2(new_n266), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n268), .A2(new_n270), .A3(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n221), .ZN(new_n276));
  INV_X1    g0076(.A(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(KEYINPUT67), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n278), .A2(new_n204), .A3(new_n257), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT67), .B1(G20), .B2(G33), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n257), .A2(G20), .ZN(new_n282));
  AOI22_X1  g0082(.A1(new_n281), .A2(G50), .B1(G77), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n213), .A2(G20), .ZN(new_n284));
  AOI21_X1  g0084(.A(new_n277), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n276), .B1(new_n203), .B2(G20), .ZN(new_n286));
  AOI22_X1  g0086(.A1(new_n285), .A2(KEYINPUT11), .B1(G68), .B2(new_n286), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n213), .ZN(new_n290));
  XNOR2_X1  g0090(.A(new_n290), .B(KEYINPUT12), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n287), .B(new_n291), .C1(KEYINPUT11), .C2(new_n285), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT72), .ZN(new_n293));
  OR2_X1    g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n292), .A2(new_n293), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT73), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n268), .A2(new_n270), .A3(new_n298), .A4(new_n272), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n274), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT8), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G58), .ZN(new_n302));
  INV_X1    g0102(.A(G58), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT8), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n281), .A2(new_n305), .B1(G20), .B2(G77), .ZN(new_n306));
  OR2_X1    g0106(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n306), .A2(KEYINPUT71), .ZN(new_n308));
  INV_X1    g0108(.A(new_n282), .ZN(new_n309));
  OR2_X1    g0109(.A1(KEYINPUT15), .A2(G87), .ZN(new_n310));
  NAND2_X1  g0110(.A1(KEYINPUT15), .A2(G87), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n307), .B(new_n308), .C1(new_n309), .C2(new_n312), .ZN(new_n313));
  AOI22_X1  g0113(.A1(new_n313), .A2(new_n276), .B1(new_n242), .B2(new_n289), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n286), .A2(G77), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n249), .A2(G232), .A3(new_n250), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n249), .A2(G1698), .ZN(new_n318));
  OAI221_X1 g0118(.A(new_n317), .B1(new_n237), .B2(new_n249), .C1(new_n318), .C2(new_n214), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT70), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n260), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n248), .B1(new_n263), .B2(G244), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT69), .B(G179), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  AND2_X1   g0125(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n322), .A2(new_n323), .ZN(new_n327));
  INV_X1    g0127(.A(G169), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n300), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n322), .A2(G190), .A3(new_n323), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n316), .B1(G200), .B2(new_n327), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n331), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n253), .A2(new_n254), .ZN(new_n335));
  AOI21_X1  g0135(.A(KEYINPUT7), .B1(new_n335), .B2(new_n204), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  NOR4_X1   g0137(.A1(new_n253), .A2(new_n254), .A3(new_n337), .A4(G20), .ZN(new_n338));
  OAI21_X1  g0138(.A(G68), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT74), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  OAI211_X1 g0141(.A(KEYINPUT74), .B(G68), .C1(new_n336), .C2(new_n338), .ZN(new_n342));
  XNOR2_X1  g0142(.A(G58), .B(G68), .ZN(new_n343));
  AOI22_X1  g0143(.A1(new_n281), .A2(G159), .B1(new_n343), .B2(G20), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n341), .A2(new_n342), .A3(KEYINPUT16), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n339), .A2(new_n344), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT16), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n345), .A2(new_n276), .A3(new_n348), .ZN(new_n349));
  XNOR2_X1  g0149(.A(KEYINPUT8), .B(G58), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(KEYINPUT66), .ZN(new_n351));
  OR2_X1    g0151(.A1(new_n302), .A2(KEYINPUT66), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n288), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n354), .B1(new_n286), .B2(new_n353), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(KEYINPUT75), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT75), .ZN(new_n357));
  OAI211_X1 g0157(.A(new_n354), .B(new_n357), .C1(new_n286), .C2(new_n353), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n349), .A2(new_n359), .ZN(new_n360));
  OAI211_X1 g0160(.A(G226), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n361));
  OAI211_X1 g0161(.A(G223), .B(new_n250), .C1(new_n253), .C2(new_n254), .ZN(new_n362));
  INV_X1    g0162(.A(G87), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n362), .C1(new_n257), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n364), .A2(new_n260), .ZN(new_n365));
  AND3_X1   g0165(.A1(new_n259), .A2(G232), .A3(new_n245), .ZN(new_n366));
  INV_X1    g0166(.A(new_n366), .ZN(new_n367));
  NAND4_X1  g0167(.A1(new_n365), .A2(new_n247), .A3(new_n324), .A4(new_n367), .ZN(new_n368));
  AOI211_X1 g0168(.A(new_n366), .B(new_n248), .C1(new_n364), .C2(new_n260), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n368), .B1(new_n369), .B2(G169), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT18), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n360), .A2(KEYINPUT18), .A3(new_n371), .ZN(new_n375));
  INV_X1    g0175(.A(G190), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n365), .A2(new_n376), .A3(new_n247), .A4(new_n367), .ZN(new_n377));
  OAI21_X1  g0177(.A(new_n377), .B1(new_n369), .B2(G200), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n349), .A2(new_n359), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT17), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT17), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n349), .A2(new_n381), .A3(new_n359), .A4(new_n378), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n374), .A2(new_n375), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n263), .A2(G226), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n335), .A2(G1698), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(G222), .B1(G77), .B2(new_n335), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n335), .A2(new_n250), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(G223), .ZN(new_n388));
  AND2_X1   g0188(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n247), .B(new_n384), .C1(new_n389), .C2(new_n259), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(new_n376), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n281), .A2(G150), .ZN(new_n392));
  OAI21_X1  g0192(.A(new_n392), .B1(new_n353), .B2(new_n309), .ZN(new_n393));
  NOR2_X1   g0193(.A1(G58), .A2(G68), .ZN(new_n394));
  INV_X1    g0194(.A(G50), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n204), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  XOR2_X1   g0196(.A(new_n396), .B(KEYINPUT68), .Z(new_n397));
  OAI21_X1  g0197(.A(new_n276), .B1(new_n393), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n289), .A2(new_n395), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n286), .A2(G50), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT9), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND4_X1  g0203(.A1(new_n398), .A2(KEYINPUT9), .A3(new_n399), .A4(new_n400), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n390), .A2(G200), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n391), .A2(new_n403), .A3(new_n404), .A4(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(new_n406), .B(KEYINPUT10), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n390), .A2(new_n328), .ZN(new_n408));
  INV_X1    g0208(.A(new_n324), .ZN(new_n409));
  OAI211_X1 g0209(.A(new_n408), .B(new_n401), .C1(new_n409), .C2(new_n390), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n269), .A2(G190), .ZN(new_n413));
  INV_X1    g0213(.A(G200), .ZN(new_n414));
  OAI211_X1 g0214(.A(new_n296), .B(new_n413), .C1(new_n414), .C2(new_n269), .ZN(new_n415));
  NAND4_X1  g0215(.A1(new_n334), .A2(new_n383), .A3(new_n412), .A4(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n203), .A2(G33), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n277), .A2(new_n288), .A3(new_n417), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n418), .A2(new_n237), .ZN(new_n419));
  NAND2_X1  g0219(.A1(G33), .A2(G116), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n420), .A2(G20), .ZN(new_n421));
  OAI211_X1 g0221(.A(new_n204), .B(G87), .C1(new_n253), .C2(new_n254), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT22), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT22), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n249), .A2(new_n424), .A3(new_n204), .A4(G87), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n421), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(new_n204), .A2(G107), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT23), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(KEYINPUT24), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT24), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n426), .A2(new_n431), .A3(new_n428), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(new_n419), .B1(new_n433), .B2(new_n276), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n387), .A2(G257), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n385), .A2(G250), .ZN(new_n436));
  XOR2_X1   g0236(.A(KEYINPUT80), .B(G294), .Z(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(G33), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G45), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n440), .A2(G1), .ZN(new_n441));
  NAND2_X1  g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g0243(.A1(KEYINPUT5), .A2(G41), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(new_n259), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n439), .A2(new_n260), .B1(G264), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n203), .A2(G45), .ZN(new_n449));
  OR2_X1    g0249(.A1(KEYINPUT5), .A2(G41), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(new_n442), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n451), .A2(G274), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(G200), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n448), .A2(G190), .A3(new_n452), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n288), .A2(G107), .ZN(new_n456));
  XNOR2_X1  g0256(.A(new_n456), .B(KEYINPUT25), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n434), .A2(new_n454), .A3(new_n455), .A4(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(G244), .B(new_n250), .C1(new_n253), .C2(new_n254), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT4), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n250), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n249), .A2(G250), .A3(G1698), .ZN(new_n463));
  NAND2_X1  g0263(.A1(G33), .A2(G283), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n260), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n452), .B1(new_n446), .B2(new_n216), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(G190), .A3(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n288), .A2(G97), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n418), .A2(new_n215), .ZN(new_n471));
  OAI21_X1  g0271(.A(G107), .B1(new_n336), .B2(new_n338), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT6), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n215), .A2(new_n237), .ZN(new_n474));
  NOR2_X1   g0274(.A1(G97), .A2(G107), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n237), .A2(KEYINPUT6), .A3(G97), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G20), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n281), .A2(G77), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n472), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI211_X1 g0281(.A(new_n470), .B(new_n471), .C1(new_n481), .C2(new_n276), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT76), .ZN(new_n483));
  AND3_X1   g0283(.A1(new_n465), .A2(new_n483), .A3(new_n260), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n483), .B1(new_n465), .B2(new_n260), .ZN(new_n485));
  NOR3_X1   g0285(.A1(new_n484), .A2(new_n485), .A3(new_n467), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n469), .B(new_n482), .C1(new_n486), .C2(new_n414), .ZN(new_n487));
  INV_X1    g0287(.A(new_n485), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n465), .A2(new_n483), .A3(new_n260), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n488), .A2(new_n324), .A3(new_n468), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n470), .B1(new_n481), .B2(new_n276), .ZN(new_n491));
  INV_X1    g0291(.A(new_n471), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n466), .A2(new_n468), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n328), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n490), .A2(new_n493), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n289), .A2(new_n209), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n275), .A2(new_n221), .B1(G20), .B2(new_n209), .ZN(new_n498));
  OAI211_X1 g0298(.A(new_n464), .B(new_n204), .C1(G33), .C2(new_n215), .ZN(new_n499));
  AND3_X1   g0299(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(KEYINPUT20), .B1(new_n498), .B2(new_n499), .ZN(new_n501));
  OAI221_X1 g0301(.A(new_n497), .B1(new_n418), .B2(new_n209), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n445), .A2(G270), .A3(new_n259), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n452), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n504), .A2(KEYINPUT79), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n249), .A2(G257), .A3(new_n250), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n249), .A2(G264), .A3(G1698), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n335), .A2(G303), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n509), .A2(new_n260), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT79), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n503), .A2(new_n452), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n505), .A2(new_n510), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g0313(.A(new_n502), .B1(new_n513), .B2(G200), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n376), .B2(new_n513), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n458), .A2(new_n487), .A3(new_n496), .A4(new_n515), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n503), .A2(new_n452), .A3(new_n511), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n511), .B1(new_n503), .B2(new_n452), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n328), .B1(new_n519), .B2(new_n510), .ZN(new_n520));
  AOI21_X1  g0320(.A(KEYINPUT21), .B1(new_n520), .B2(new_n502), .ZN(new_n521));
  NAND4_X1  g0321(.A1(new_n513), .A2(KEYINPUT21), .A3(G169), .A4(new_n502), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n519), .A2(new_n502), .A3(G179), .A4(new_n510), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  AND3_X1   g0325(.A1(new_n426), .A2(new_n431), .A3(new_n428), .ZN(new_n526));
  AOI21_X1  g0326(.A(new_n431), .B1(new_n426), .B2(new_n428), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n276), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n419), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n528), .A2(new_n529), .A3(new_n457), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n453), .A2(new_n328), .ZN(new_n531));
  INV_X1    g0331(.A(G179), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n448), .A2(new_n532), .A3(new_n452), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  AND3_X1   g0334(.A1(new_n277), .A2(new_n288), .A3(new_n417), .ZN(new_n535));
  INV_X1    g0335(.A(new_n312), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT78), .ZN(new_n538));
  NAND3_X1  g0338(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n204), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n363), .A2(new_n215), .A3(new_n237), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n204), .B(G68), .C1(new_n253), .C2(new_n254), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n204), .A2(G33), .A3(G97), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT19), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n276), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n288), .B1(new_n310), .B2(new_n311), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n538), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  AOI211_X1 g0351(.A(KEYINPUT78), .B(new_n549), .C1(new_n547), .C2(new_n276), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n537), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(G244), .B(G1698), .C1(new_n253), .C2(new_n254), .ZN(new_n554));
  OAI211_X1 g0354(.A(G238), .B(new_n250), .C1(new_n253), .C2(new_n254), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n554), .A2(new_n555), .A3(new_n420), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n556), .A2(new_n260), .B1(G274), .B2(new_n441), .ZN(new_n557));
  AND2_X1   g0357(.A1(G33), .A2(G41), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n449), .B(G250), .C1(new_n558), .C2(new_n221), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT77), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n259), .A2(KEYINPUT77), .A3(G250), .A4(new_n449), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n557), .A2(new_n324), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n556), .A2(new_n260), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n441), .A2(G274), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n565), .A2(new_n566), .A3(new_n563), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n328), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n553), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n548), .A2(new_n538), .A3(new_n550), .ZN(new_n570));
  AOI22_X1  g0370(.A1(new_n540), .A2(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n277), .B1(new_n571), .B2(new_n543), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT78), .B1(new_n572), .B2(new_n549), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n535), .A2(G87), .ZN(new_n575));
  AND4_X1   g0375(.A1(new_n376), .A2(new_n565), .A3(new_n566), .A4(new_n563), .ZN(new_n576));
  AOI21_X1  g0376(.A(G200), .B1(new_n557), .B2(new_n563), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n574), .B(new_n575), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n569), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n525), .A2(new_n534), .A3(new_n579), .ZN(new_n580));
  NOR3_X1   g0380(.A1(new_n416), .A2(new_n516), .A3(new_n580), .ZN(G372));
  NAND2_X1  g0381(.A1(new_n380), .A2(new_n382), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n331), .A2(new_n582), .A3(new_n415), .ZN(new_n583));
  INV_X1    g0383(.A(new_n375), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT18), .B1(new_n360), .B2(new_n371), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n407), .B1(new_n583), .B2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n587), .A2(new_n410), .ZN(new_n588));
  AND4_X1   g0388(.A1(new_n334), .A2(new_n383), .A3(new_n412), .A4(new_n415), .ZN(new_n589));
  INV_X1    g0389(.A(new_n569), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT82), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n525), .A2(new_n534), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n591), .B1(new_n525), .B2(new_n534), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  AND3_X1   g0394(.A1(new_n569), .A2(KEYINPUT81), .A3(new_n578), .ZN(new_n595));
  AOI21_X1  g0395(.A(KEYINPUT81), .B1(new_n569), .B2(new_n578), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n458), .A2(new_n487), .A3(new_n496), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n590), .B1(new_n594), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n576), .A2(new_n577), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n574), .A2(new_n575), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n568), .A2(new_n564), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n570), .A2(new_n573), .B1(new_n536), .B2(new_n535), .ZN(new_n604));
  OAI22_X1  g0404(.A1(new_n601), .A2(new_n602), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT81), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n569), .A2(KEYINPUT81), .A3(new_n578), .ZN(new_n608));
  AOI21_X1  g0408(.A(new_n496), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(KEYINPUT83), .B1(new_n609), .B2(KEYINPUT26), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n605), .A2(new_n496), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(KEYINPUT26), .ZN(new_n612));
  INV_X1    g0412(.A(new_n496), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n613), .B1(new_n595), .B2(new_n596), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT83), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT26), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n614), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n610), .A2(new_n612), .A3(new_n617), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n600), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n589), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n588), .A2(new_n620), .ZN(G369));
  INV_X1    g0421(.A(new_n458), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n203), .A2(new_n204), .A3(G13), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g0426(.A(new_n626), .B(KEYINPUT84), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(G343), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  AND2_X1   g0430(.A1(new_n530), .A2(new_n630), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n534), .B1(new_n622), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT85), .ZN(new_n633));
  OR2_X1    g0433(.A1(new_n534), .A2(new_n630), .ZN(new_n634));
  AND3_X1   g0434(.A1(new_n632), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n633), .B1(new_n632), .B2(new_n634), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n525), .A2(new_n630), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n640), .A2(new_n634), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n630), .A2(new_n502), .ZN(new_n642));
  XNOR2_X1  g0442(.A(new_n525), .B(new_n642), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n643), .A2(new_n515), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(G330), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n637), .A2(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n641), .A2(new_n647), .ZN(G399));
  INV_X1    g0448(.A(new_n205), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n649), .A2(G41), .ZN(new_n650));
  INV_X1    g0450(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n541), .A2(G116), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n651), .A2(G1), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n653), .B1(new_n223), .B2(new_n651), .ZN(new_n654));
  XNOR2_X1  g0454(.A(new_n654), .B(KEYINPUT28), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n607), .A2(new_n608), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n525), .A2(new_n534), .ZN(new_n657));
  AND2_X1   g0457(.A1(new_n487), .A2(new_n496), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(new_n458), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n614), .A2(KEYINPUT26), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n590), .B1(new_n611), .B2(new_n616), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n630), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT87), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(KEYINPUT87), .A3(new_n663), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(KEYINPUT29), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n630), .B1(new_n600), .B2(new_n618), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT29), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G330), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n494), .A2(new_n567), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n513), .A2(new_n532), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n674), .A2(new_n675), .A3(new_n448), .ZN(new_n676));
  INV_X1    g0476(.A(KEYINPUT30), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n674), .A2(new_n675), .A3(KEYINPUT30), .A4(new_n448), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n488), .A2(new_n468), .A3(new_n489), .ZN(new_n680));
  AOI21_X1  g0480(.A(new_n409), .B1(new_n557), .B2(new_n563), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n680), .A2(new_n453), .A3(new_n513), .A4(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n678), .A2(new_n679), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n683), .A2(new_n630), .ZN(new_n684));
  NOR3_X1   g0484(.A1(new_n516), .A2(new_n580), .A3(new_n630), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT31), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n684), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n683), .A2(KEYINPUT31), .A3(new_n630), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT86), .ZN(new_n689));
  XNOR2_X1  g0489(.A(new_n688), .B(new_n689), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n673), .B1(new_n687), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n672), .A2(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n655), .B1(new_n692), .B2(G1), .ZN(new_n693));
  XOR2_X1   g0493(.A(new_n693), .B(KEYINPUT88), .Z(G364));
  NAND2_X1  g0494(.A1(new_n204), .A2(G13), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT89), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G45), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n697), .A2(G1), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(new_n650), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n645), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n644), .A2(G330), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n700), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n204), .A2(G179), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n704), .A2(G190), .A3(G200), .ZN(new_n705));
  INV_X1    g0505(.A(G303), .ZN(new_n706));
  INV_X1    g0506(.A(G283), .ZN(new_n707));
  NAND3_X1  g0507(.A1(new_n704), .A2(new_n376), .A3(G200), .ZN(new_n708));
  OAI221_X1 g0508(.A(new_n335), .B1(new_n705), .B2(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n324), .A2(new_n204), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT91), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(G190), .A3(G200), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  XOR2_X1   g0513(.A(KEYINPUT94), .B(G326), .Z(new_n714));
  NOR3_X1   g0514(.A1(new_n376), .A2(G179), .A3(G200), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n715), .A2(new_n204), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  AOI22_X1  g0517(.A1(new_n713), .A2(new_n714), .B1(new_n437), .B2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n719));
  AND3_X1   g0519(.A1(new_n711), .A2(new_n376), .A3(new_n414), .ZN(new_n720));
  AOI211_X1 g0520(.A(new_n709), .B(new_n719), .C1(G311), .C2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n704), .A2(new_n376), .A3(new_n414), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G329), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n711), .A2(G190), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n725), .A2(G200), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n711), .A2(new_n376), .A3(G200), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT33), .B(G317), .ZN(new_n729));
  AOI22_X1  g0529(.A1(G322), .A2(new_n726), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT96), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n718), .A2(KEYINPUT95), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n721), .A2(new_n724), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  OAI22_X1  g0533(.A1(new_n727), .A2(new_n213), .B1(new_n215), .B2(new_n716), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT93), .ZN(new_n735));
  AOI22_X1  g0535(.A1(new_n726), .A2(G58), .B1(new_n720), .B2(G77), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n249), .B1(new_n705), .B2(new_n363), .C1(new_n237), .C2(new_n708), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n713), .B2(G50), .ZN(new_n738));
  NAND3_X1  g0538(.A1(new_n735), .A2(new_n736), .A3(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(G159), .ZN(new_n740));
  NOR2_X1   g0540(.A1(new_n722), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g0541(.A(KEYINPUT92), .B(KEYINPUT32), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n741), .B(new_n742), .Z(new_n743));
  OAI21_X1  g0543(.A(new_n733), .B1(new_n739), .B2(new_n743), .ZN(new_n744));
  AOI21_X1  g0544(.A(new_n221), .B1(G20), .B2(new_n328), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n649), .A2(new_n249), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n224), .A2(new_n440), .ZN(new_n748));
  OAI211_X1 g0548(.A(new_n747), .B(new_n748), .C1(new_n243), .C2(new_n440), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n249), .A2(new_n205), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT90), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n751), .A2(G355), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n749), .B(new_n752), .C1(G116), .C2(new_n205), .ZN(new_n753));
  NOR2_X1   g0553(.A1(G13), .A2(G33), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G20), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n756), .A2(new_n745), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n756), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n746), .B(new_n758), .C1(new_n644), .C2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n703), .B1(new_n761), .B2(new_n700), .ZN(new_n762));
  XOR2_X1   g0562(.A(new_n762), .B(KEYINPUT97), .Z(G396));
  NAND3_X1  g0563(.A1(new_n326), .A2(new_n329), .A3(new_n630), .ZN(new_n764));
  INV_X1    g0564(.A(KEYINPUT98), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n326), .A2(KEYINPUT98), .A3(new_n329), .A4(new_n630), .ZN(new_n767));
  AOI22_X1  g0567(.A1(new_n333), .A2(new_n332), .B1(new_n316), .B2(new_n630), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(new_n767), .B1(new_n768), .B2(new_n330), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n669), .B(new_n770), .ZN(new_n771));
  XNOR2_X1  g0571(.A(new_n771), .B(new_n691), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(new_n700), .ZN(new_n773));
  AOI22_X1  g0573(.A1(G137), .A2(new_n713), .B1(new_n728), .B2(G150), .ZN(new_n774));
  INV_X1    g0574(.A(new_n720), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n774), .B1(new_n740), .B2(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n776), .B1(G143), .B2(new_n726), .ZN(new_n777));
  XOR2_X1   g0577(.A(new_n777), .B(KEYINPUT34), .Z(new_n778));
  NOR2_X1   g0578(.A1(new_n708), .A2(new_n213), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n249), .B1(new_n716), .B2(new_n303), .ZN(new_n780));
  INV_X1    g0580(.A(new_n705), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n779), .B(new_n780), .C1(G50), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(G132), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n778), .B(new_n782), .C1(new_n783), .C2(new_n722), .ZN(new_n784));
  INV_X1    g0584(.A(new_n708), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n785), .A2(G87), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n786), .B1(new_n215), .B2(new_n716), .C1(new_n237), .C2(new_n705), .ZN(new_n787));
  INV_X1    g0587(.A(G311), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n335), .B1(new_n722), .B2(new_n788), .ZN(new_n789));
  AOI211_X1 g0589(.A(new_n787), .B(new_n789), .C1(new_n728), .C2(G283), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n726), .A2(G294), .B1(new_n720), .B2(G116), .ZN(new_n791));
  OAI211_X1 g0591(.A(new_n790), .B(new_n791), .C1(new_n706), .C2(new_n712), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n745), .A2(new_n754), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n793), .A2(new_n745), .B1(new_n242), .B2(new_n794), .ZN(new_n795));
  OAI211_X1 g0595(.A(new_n795), .B(new_n699), .C1(new_n755), .C2(new_n770), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n773), .A2(new_n796), .ZN(G384));
  AOI21_X1  g0597(.A(new_n769), .B1(new_n687), .B2(new_n688), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n300), .A2(new_n415), .ZN(new_n799));
  NAND3_X1  g0599(.A1(new_n294), .A2(new_n295), .A3(new_n630), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n800), .B(KEYINPUT100), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n803));
  OR2_X1    g0603(.A1(new_n800), .A2(KEYINPUT100), .ZN(new_n804));
  NAND4_X1  g0604(.A1(new_n300), .A2(new_n415), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g0606(.A1(new_n798), .A2(KEYINPUT40), .A3(new_n806), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n360), .A2(new_n627), .ZN(new_n808));
  OAI21_X1  g0608(.A(KEYINPUT103), .B1(new_n383), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n582), .B1(new_n584), .B2(new_n585), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT103), .ZN(new_n811));
  INV_X1    g0611(.A(new_n808), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n810), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n349), .A2(new_n359), .B1(new_n370), .B2(new_n628), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT37), .ZN(new_n816));
  NAND3_X1  g0616(.A1(new_n815), .A2(new_n816), .A3(new_n379), .ZN(new_n817));
  INV_X1    g0617(.A(new_n379), .ZN(new_n818));
  OAI21_X1  g0618(.A(KEYINPUT37), .B1(new_n818), .B2(new_n814), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT102), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n815), .A2(KEYINPUT102), .A3(new_n816), .A4(new_n379), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n809), .A2(new_n813), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT38), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n341), .A2(new_n344), .A3(new_n342), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n347), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n827), .A2(new_n276), .A3(new_n345), .ZN(new_n828));
  AOI22_X1  g0628(.A1(new_n828), .A2(new_n359), .B1(new_n370), .B2(new_n628), .ZN(new_n829));
  OAI21_X1  g0629(.A(KEYINPUT37), .B1(new_n829), .B2(new_n818), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n830), .A2(KEYINPUT101), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT101), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n832), .B(KEYINPUT37), .C1(new_n829), .C2(new_n818), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n831), .A2(new_n817), .A3(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n828), .A2(new_n359), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n810), .A2(new_n627), .A3(new_n835), .ZN(new_n836));
  NAND3_X1  g0636(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n825), .A2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(KEYINPUT106), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n825), .A2(KEYINPUT106), .A3(new_n837), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n807), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n798), .A2(new_n806), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n834), .A2(new_n836), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n824), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n845), .A2(new_n837), .ZN(new_n846));
  AOI21_X1  g0646(.A(KEYINPUT40), .B1(new_n843), .B2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n842), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(new_n416), .B1(new_n687), .B2(new_n688), .ZN(new_n849));
  XOR2_X1   g0649(.A(new_n848), .B(new_n849), .Z(new_n850));
  NAND2_X1  g0650(.A1(new_n850), .A2(G330), .ZN(new_n851));
  AND3_X1   g0651(.A1(new_n662), .A2(KEYINPUT87), .A3(new_n663), .ZN(new_n852));
  AOI21_X1  g0652(.A(KEYINPUT87), .B1(new_n662), .B2(new_n663), .ZN(new_n853));
  NOR3_X1   g0653(.A1(new_n852), .A2(new_n853), .A3(new_n670), .ZN(new_n854));
  AOI211_X1 g0654(.A(KEYINPUT29), .B(new_n630), .C1(new_n600), .C2(new_n618), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n589), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT105), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT105), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n672), .A2(new_n858), .A3(new_n589), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n588), .ZN(new_n861));
  XNOR2_X1  g0661(.A(new_n851), .B(new_n861), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n300), .A2(new_n630), .ZN(new_n863));
  INV_X1    g0663(.A(new_n863), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n825), .A2(new_n865), .A3(new_n837), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(new_n845), .B2(new_n837), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AND3_X1   g0669(.A1(new_n834), .A2(KEYINPUT38), .A3(new_n836), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n824), .B2(new_n823), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT104), .A3(new_n865), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n864), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  AND3_X1   g0673(.A1(new_n619), .A2(new_n663), .A3(new_n770), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n330), .A2(new_n630), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n846), .B(new_n806), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n586), .A2(new_n628), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NOR2_X1   g0678(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g0679(.A(new_n862), .B(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n880), .B1(new_n203), .B2(new_n696), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n209), .B1(new_n478), .B2(KEYINPUT35), .ZN(new_n882));
  OAI211_X1 g0682(.A(new_n882), .B(new_n222), .C1(KEYINPUT35), .C2(new_n478), .ZN(new_n883));
  XNOR2_X1  g0683(.A(new_n883), .B(KEYINPUT36), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT99), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n213), .B2(G50), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n395), .A2(KEYINPUT99), .A3(G68), .ZN(new_n887));
  OAI21_X1  g0687(.A(G77), .B1(new_n303), .B2(new_n213), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n886), .B(new_n887), .C1(new_n888), .C2(new_n223), .ZN(new_n889));
  INV_X1    g0689(.A(G13), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(G1), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n881), .A2(new_n884), .A3(new_n891), .ZN(G367));
  INV_X1    g0692(.A(new_n726), .ZN(new_n893));
  INV_X1    g0693(.A(G150), .ZN(new_n894));
  OAI22_X1  g0694(.A1(new_n893), .A2(new_n894), .B1(new_n775), .B2(new_n395), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n249), .B1(new_n708), .B2(new_n242), .ZN(new_n896));
  OR2_X1    g0696(.A1(new_n896), .A2(KEYINPUT111), .ZN(new_n897));
  OAI221_X1 g0697(.A(new_n897), .B1(new_n303), .B2(new_n705), .C1(new_n213), .C2(new_n716), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n898), .B1(KEYINPUT111), .B2(new_n896), .ZN(new_n899));
  INV_X1    g0699(.A(G137), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n899), .B1(new_n900), .B2(new_n722), .C1(new_n740), .C2(new_n727), .ZN(new_n901));
  AOI211_X1 g0701(.A(new_n895), .B(new_n901), .C1(G143), .C2(new_n713), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n785), .A2(G97), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n903), .B1(new_n237), .B2(new_n716), .ZN(new_n904));
  AOI211_X1 g0704(.A(new_n249), .B(new_n904), .C1(G317), .C2(new_n723), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n781), .A2(G116), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n906), .B(KEYINPUT46), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n905), .B(new_n907), .C1(new_n712), .C2(new_n788), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n728), .A2(new_n437), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n893), .B2(new_n706), .ZN(new_n910));
  AOI211_X1 g0710(.A(new_n908), .B(new_n910), .C1(G283), .C2(new_n720), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n902), .A2(new_n911), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT47), .Z(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n745), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n630), .A2(new_n602), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n915), .A2(new_n569), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n916), .B1(new_n656), .B2(new_n915), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n756), .ZN(new_n918));
  INV_X1    g0718(.A(new_n747), .ZN(new_n919));
  OAI221_X1 g0719(.A(new_n757), .B1(new_n205), .B2(new_n312), .C1(new_n233), .C2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n920), .A2(new_n699), .ZN(new_n921));
  XNOR2_X1  g0721(.A(new_n921), .B(KEYINPUT110), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n914), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n698), .ZN(new_n925));
  INV_X1    g0725(.A(new_n692), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT44), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n658), .B1(new_n482), .B2(new_n663), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n613), .A2(new_n630), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n927), .B1(new_n641), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n640), .A2(new_n634), .ZN(new_n932));
  NAND4_X1  g0732(.A1(new_n932), .A2(KEYINPUT44), .A3(new_n928), .A4(new_n929), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n640), .A2(new_n634), .A3(new_n930), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT45), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n935), .B(new_n936), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n934), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n938), .A2(KEYINPUT109), .A3(new_n647), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n647), .A2(KEYINPUT109), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n647), .A2(KEYINPUT109), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n934), .A2(new_n937), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n939), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n637), .B1(new_n525), .B2(new_n630), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n640), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n945), .B(new_n701), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n692), .ZN(new_n947));
  INV_X1    g0747(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n926), .B1(new_n943), .B2(new_n948), .ZN(new_n949));
  XOR2_X1   g0749(.A(new_n650), .B(KEYINPUT41), .Z(new_n950));
  OAI21_X1  g0750(.A(new_n925), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n638), .A2(new_n639), .A3(new_n930), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT42), .Z(new_n953));
  INV_X1    g0753(.A(new_n487), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n496), .B1(new_n954), .B2(new_n534), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n663), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT43), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n917), .B(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OR2_X1    g0760(.A1(new_n917), .A2(new_n958), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n959), .A2(new_n958), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n953), .A2(new_n962), .A3(new_n956), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n646), .A2(KEYINPUT108), .A3(new_n930), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n960), .A2(new_n961), .A3(new_n963), .A4(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(KEYINPUT108), .B1(new_n646), .B2(new_n930), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n965), .B(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n924), .B1(new_n951), .B2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n968), .ZN(G387));
  OR2_X1    g0769(.A1(new_n946), .A2(new_n692), .ZN(new_n970));
  NAND3_X1  g0770(.A1(new_n970), .A2(new_n650), .A3(new_n947), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n638), .A2(new_n759), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n350), .A2(G50), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT50), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n652), .B1(new_n213), .B2(new_n242), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  AOI211_X1 g0775(.A(G45), .B(new_n975), .C1(new_n974), .C2(new_n973), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n747), .B1(new_n230), .B2(new_n440), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n751), .B1(G116), .B2(new_n541), .ZN(new_n978));
  AOI21_X1  g0778(.A(new_n976), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  NOR2_X1   g0779(.A1(new_n205), .A2(G107), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR3_X1   g0781(.A1(new_n981), .A2(new_n756), .A3(new_n745), .ZN(new_n982));
  AOI22_X1  g0782(.A1(new_n726), .A2(G317), .B1(new_n720), .B2(G303), .ZN(new_n983));
  INV_X1    g0783(.A(G322), .ZN(new_n984));
  OAI221_X1 g0784(.A(new_n983), .B1(new_n788), .B2(new_n727), .C1(new_n984), .C2(new_n712), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n985), .B(KEYINPUT48), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n781), .A2(new_n437), .ZN(new_n987));
  OAI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(new_n707), .C2(new_n716), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT49), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n723), .A2(new_n714), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n988), .A2(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n249), .B1(new_n785), .B2(G116), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n990), .A2(new_n991), .A3(new_n992), .A4(new_n993), .ZN(new_n994));
  OAI22_X1  g0794(.A1(new_n775), .A2(new_n213), .B1(new_n353), .B2(new_n727), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT112), .ZN(new_n996));
  NOR2_X1   g0796(.A1(new_n716), .A2(new_n312), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n705), .A2(new_n242), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n894), .B2(new_n722), .ZN(new_n1000));
  NOR2_X1   g0800(.A1(new_n712), .A2(new_n740), .ZN(new_n1001));
  AOI211_X1 g0801(.A(new_n1000), .B(new_n1001), .C1(G50), .C2(new_n726), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n996), .A2(new_n249), .A3(new_n903), .A4(new_n1002), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n994), .A2(new_n1003), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n972), .B(new_n982), .C1(new_n1004), .C2(new_n745), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n1005), .A2(new_n699), .B1(new_n698), .B2(new_n946), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n971), .A2(new_n1006), .ZN(G393));
  NAND2_X1  g0807(.A1(new_n943), .A2(new_n698), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G50), .A2(new_n728), .B1(new_n720), .B2(new_n305), .ZN(new_n1009));
  INV_X1    g0809(.A(new_n1009), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT113), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n705), .A2(new_n213), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n716), .A2(new_n242), .ZN(new_n1013));
  AOI211_X1 g0813(.A(new_n1012), .B(new_n1013), .C1(G143), .C2(new_n723), .ZN(new_n1014));
  AND4_X1   g0814(.A1(new_n249), .A2(new_n1011), .A3(new_n786), .A4(new_n1014), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n893), .A2(new_n740), .B1(new_n894), .B2(new_n712), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT51), .ZN(new_n1017));
  AOI22_X1  g0817(.A1(KEYINPUT113), .A2(new_n1010), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OAI211_X1 g0818(.A(new_n1015), .B(new_n1018), .C1(new_n1017), .C2(new_n1016), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(G311), .A2(new_n726), .B1(new_n713), .B2(G317), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT52), .Z(new_n1021));
  INV_X1    g0821(.A(G294), .ZN(new_n1022));
  OAI221_X1 g0822(.A(new_n335), .B1(new_n984), .B2(new_n722), .C1(new_n775), .C2(new_n1022), .ZN(new_n1023));
  AOI22_X1  g0823(.A1(new_n728), .A2(G303), .B1(G116), .B2(new_n717), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n1023), .B1(new_n1024), .B2(KEYINPUT114), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n1024), .A2(KEYINPUT114), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n781), .A2(G283), .B1(new_n785), .B2(G107), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1019), .A2(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n700), .B1(new_n1029), .B2(new_n745), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n239), .A2(new_n747), .B1(G97), .B2(new_n649), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n757), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n928), .A2(new_n756), .A3(new_n929), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1030), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1008), .A2(KEYINPUT115), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(KEYINPUT115), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n925), .B1(new_n939), .B2(new_n942), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1034), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1035), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n943), .A2(new_n948), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n939), .A2(new_n947), .A3(new_n942), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1041), .A2(new_n650), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1040), .A2(new_n1043), .ZN(G390));
  INV_X1    g0844(.A(new_n806), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n669), .A2(new_n770), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n875), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1045), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n869), .B(new_n872), .C1(new_n863), .C2(new_n1048), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n840), .A2(new_n841), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n769), .B1(new_n666), .B2(new_n667), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n806), .B1(new_n1051), .B2(new_n875), .ZN(new_n1052));
  NAND3_X1  g0852(.A1(new_n1050), .A2(new_n864), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1049), .A2(new_n1053), .ZN(new_n1054));
  AND3_X1   g0854(.A1(new_n798), .A2(G330), .A3(new_n806), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  NAND3_X1  g0857(.A1(new_n691), .A2(new_n770), .A3(new_n806), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n1058), .ZN(new_n1059));
  NAND3_X1  g0859(.A1(new_n1049), .A2(new_n1053), .A3(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1057), .A2(new_n1060), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n849), .A2(G330), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n806), .B1(new_n691), .B2(new_n770), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1063), .B1(new_n1055), .B2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n684), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n516), .A2(new_n580), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1067), .A2(new_n663), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1066), .B1(new_n1068), .B2(KEYINPUT31), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n688), .ZN(new_n1070));
  OAI211_X1 g0870(.A(G330), .B(new_n770), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1071), .A2(new_n1045), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n770), .B1(new_n852), .B2(new_n853), .ZN(new_n1073));
  NAND4_X1  g0873(.A1(new_n1072), .A2(new_n1047), .A3(new_n1058), .A4(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1065), .A2(new_n1074), .ZN(new_n1075));
  NAND4_X1  g0875(.A1(new_n860), .A2(new_n588), .A3(new_n1062), .A4(new_n1075), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1061), .A2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n1057), .A2(new_n1076), .A3(new_n1060), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n650), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n869), .A2(new_n754), .A3(new_n872), .ZN(new_n1081));
  XOR2_X1   g0881(.A(KEYINPUT54), .B(G143), .Z(new_n1082));
  AOI22_X1  g0882(.A1(G137), .A2(new_n728), .B1(new_n720), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1083), .B1(new_n740), .B2(new_n716), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT116), .Z(new_n1085));
  NOR2_X1   g0885(.A1(new_n705), .A2(new_n894), .ZN(new_n1086));
  XOR2_X1   g0886(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1087));
  OAI221_X1 g0887(.A(new_n249), .B1(new_n395), .B2(new_n708), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1089), .B1(new_n893), .B2(new_n783), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1090), .B1(G128), .B2(new_n713), .ZN(new_n1091));
  INV_X1    g0891(.A(G125), .ZN(new_n1092));
  OAI211_X1 g0892(.A(new_n1085), .B(new_n1091), .C1(new_n1092), .C2(new_n722), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n335), .B1(new_n1022), .B2(new_n722), .C1(new_n727), .C2(new_n237), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n705), .A2(new_n363), .ZN(new_n1095));
  NOR4_X1   g0895(.A1(new_n1094), .A2(new_n1095), .A3(new_n779), .A4(new_n1013), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n726), .A2(G116), .B1(new_n720), .B2(G97), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1096), .B(new_n1097), .C1(new_n707), .C2(new_n712), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1093), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n1099), .A2(new_n745), .B1(new_n353), .B2(new_n794), .ZN(new_n1100));
  AND2_X1   g0900(.A1(new_n1081), .A2(new_n1100), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n1061), .A2(new_n698), .B1(new_n699), .B2(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1080), .A2(new_n1102), .ZN(G378));
  AOI21_X1  g0903(.A(new_n1076), .B1(new_n1057), .B2(new_n1060), .ZN(new_n1104));
  AOI211_X1 g0904(.A(KEYINPUT105), .B(new_n416), .C1(new_n668), .C2(new_n671), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n858), .B1(new_n672), .B2(new_n589), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n588), .B(new_n1062), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  INV_X1    g0907(.A(KEYINPUT121), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n860), .A2(KEYINPUT121), .A3(new_n588), .A4(new_n1062), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(KEYINPUT38), .B1(new_n834), .B2(new_n836), .ZN(new_n1112));
  OAI21_X1  g0912(.A(KEYINPUT39), .B1(new_n870), .B2(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(new_n871), .A2(new_n865), .B1(new_n1113), .B2(KEYINPUT104), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n866), .A2(new_n868), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n863), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n876), .A2(new_n877), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n401), .A2(new_n627), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n412), .A2(new_n1118), .ZN(new_n1119));
  INV_X1    g0919(.A(KEYINPUT55), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1118), .B1(new_n407), .B2(new_n410), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1119), .A2(new_n1120), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1118), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n411), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT55), .B1(new_n1125), .B2(new_n1121), .ZN(new_n1126));
  AND3_X1   g0926(.A1(new_n1123), .A2(new_n1126), .A3(KEYINPUT56), .ZN(new_n1127));
  AOI21_X1  g0927(.A(KEYINPUT56), .B1(new_n1123), .B2(new_n1126), .ZN(new_n1128));
  OR2_X1    g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1116), .A2(new_n1117), .A3(new_n1129), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1131), .B1(new_n873), .B2(new_n878), .ZN(new_n1132));
  NOR3_X1   g0932(.A1(new_n842), .A2(new_n847), .A3(new_n673), .ZN(new_n1133));
  AND3_X1   g0933(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1133), .B1(new_n1130), .B2(new_n1132), .ZN(new_n1135));
  OAI22_X1  g0935(.A1(new_n1104), .A2(new_n1111), .B1(new_n1134), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(KEYINPUT57), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1133), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1129), .B1(new_n1116), .B2(new_n1117), .ZN(new_n1140));
  NOR3_X1   g0940(.A1(new_n873), .A2(new_n878), .A3(new_n1131), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1139), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1130), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(KEYINPUT57), .C1(new_n1104), .C2(new_n1111), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1138), .A2(new_n650), .A3(new_n1145), .ZN(new_n1146));
  OAI22_X1  g0946(.A1(new_n1092), .A2(new_n712), .B1(new_n727), .B2(new_n783), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n781), .A2(new_n1082), .ZN(new_n1148));
  OAI221_X1 g0948(.A(new_n1148), .B1(new_n894), .B2(new_n716), .C1(new_n775), .C2(new_n900), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1147), .B(new_n1149), .C1(G128), .C2(new_n726), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT59), .ZN(new_n1151));
  AOI21_X1  g0951(.A(G41), .B1(new_n785), .B2(G159), .ZN(new_n1152));
  AOI21_X1  g0952(.A(G33), .B1(new_n723), .B2(G124), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n395), .B1(new_n253), .B2(G41), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1156), .A2(KEYINPUT118), .ZN(new_n1157));
  AOI211_X1 g0957(.A(G41), .B(new_n998), .C1(G68), .C2(new_n717), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n893), .B2(new_n237), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n775), .A2(new_n312), .B1(new_n215), .B2(new_n727), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n708), .A2(new_n303), .ZN(new_n1161));
  XNOR2_X1  g0961(.A(new_n1161), .B(KEYINPUT119), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n335), .B1(new_n722), .B2(new_n707), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1162), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1164), .B1(new_n209), .B2(new_n712), .ZN(new_n1165));
  INV_X1    g0965(.A(KEYINPUT58), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1157), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1154), .B(new_n1168), .C1(KEYINPUT118), .C2(new_n1156), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n1169), .A2(new_n745), .B1(new_n395), .B2(new_n794), .ZN(new_n1170));
  OAI211_X1 g0970(.A(new_n699), .B(new_n1170), .C1(new_n1129), .C2(new_n755), .ZN(new_n1171));
  XOR2_X1   g0971(.A(new_n1171), .B(KEYINPUT120), .Z(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n698), .B2(new_n1144), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1146), .A2(new_n1173), .ZN(G375));
  NAND2_X1  g0974(.A1(new_n1045), .A2(new_n754), .ZN(new_n1175));
  OAI22_X1  g0975(.A1(new_n722), .A2(new_n706), .B1(new_n705), .B2(new_n215), .ZN(new_n1176));
  XOR2_X1   g0976(.A(new_n1176), .B(KEYINPUT123), .Z(new_n1177));
  OAI211_X1 g0977(.A(new_n335), .B(new_n1177), .C1(new_n893), .C2(new_n707), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n997), .B(new_n1178), .C1(G77), .C2(new_n785), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(G116), .A2(new_n728), .B1(new_n713), .B2(G294), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n237), .C2(new_n775), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n1162), .A2(new_n335), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n1182), .A2(KEYINPUT124), .B1(new_n712), .B2(new_n783), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G150), .B2(new_n720), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n728), .A2(new_n1082), .B1(new_n1182), .B2(KEYINPUT124), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n726), .A2(G137), .B1(G50), .B2(new_n717), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1184), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(G128), .A2(new_n723), .B1(new_n781), .B2(G159), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT125), .Z(new_n1189));
  OAI21_X1  g0989(.A(new_n1181), .B1(new_n1187), .B2(new_n1189), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n1190), .A2(new_n745), .B1(new_n213), .B2(new_n794), .ZN(new_n1191));
  AND3_X1   g0991(.A1(new_n1175), .A2(new_n699), .A3(new_n1191), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(new_n1075), .B2(new_n698), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n950), .B(KEYINPUT122), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1077), .A2(new_n1194), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n1075), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1107), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1193), .B1(new_n1195), .B2(new_n1198), .ZN(G381));
  NOR2_X1   g0999(.A1(G387), .A2(G381), .ZN(new_n1200));
  INV_X1    g1000(.A(G378), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1146), .A2(new_n1201), .A3(new_n1173), .ZN(new_n1202));
  INV_X1    g1002(.A(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(G396), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1204), .A2(new_n1006), .A3(new_n971), .ZN(new_n1205));
  NOR3_X1   g1005(.A1(G390), .A2(G384), .A3(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(new_n1203), .A3(new_n1206), .ZN(G407));
  OAI211_X1 g1007(.A(G407), .B(G213), .C1(G343), .C2(new_n1202), .ZN(G409));
  NAND2_X1  g1008(.A1(G375), .A2(G378), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n629), .A2(G213), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1144), .A2(new_n698), .ZN(new_n1211));
  NAND4_X1  g1011(.A1(new_n1080), .A2(new_n1211), .A3(new_n1102), .A4(new_n1171), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1136), .A2(new_n1194), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1210), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n651), .B1(new_n1197), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1107), .A2(KEYINPUT60), .A3(new_n1196), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1076), .A3(new_n1218), .ZN(new_n1219));
  AND3_X1   g1019(.A1(new_n1219), .A2(G384), .A3(new_n1193), .ZN(new_n1220));
  AOI21_X1  g1020(.A(G384), .B1(new_n1219), .B2(new_n1193), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1220), .A2(new_n1221), .ZN(new_n1222));
  NAND3_X1  g1022(.A1(new_n1209), .A2(new_n1215), .A3(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(KEYINPUT62), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT61), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1219), .A2(new_n1193), .ZN(new_n1226));
  INV_X1    g1026(.A(G384), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1219), .A2(G384), .A3(new_n1193), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n629), .A2(G213), .A3(G2897), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1228), .A2(new_n1229), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1230), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n1232), .B1(new_n1220), .B2(new_n1221), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n1201), .B1(new_n1146), .B2(new_n1173), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1231), .B(new_n1233), .C1(new_n1234), .C2(new_n1214), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT62), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1209), .A2(new_n1236), .A3(new_n1215), .A4(new_n1222), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1224), .A2(new_n1225), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1205), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1040), .A2(new_n1043), .A3(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1240), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1243));
  OAI21_X1  g1043(.A(G387), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1240), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(G390), .A2(new_n1245), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n968), .A3(new_n1241), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1238), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1233), .A2(new_n1231), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1209), .B2(new_n1215), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1223), .B1(new_n1251), .B2(new_n1252), .ZN(new_n1253));
  AND3_X1   g1053(.A1(new_n1244), .A2(new_n1225), .A3(new_n1247), .ZN(new_n1254));
  INV_X1    g1054(.A(KEYINPUT126), .ZN(new_n1255));
  OAI21_X1  g1055(.A(new_n1255), .B1(new_n1223), .B2(new_n1252), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1222), .ZN(new_n1257));
  NOR3_X1   g1057(.A1(new_n1234), .A2(new_n1257), .A3(new_n1214), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1258), .A2(KEYINPUT126), .A3(KEYINPUT63), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .A4(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1249), .A2(new_n1260), .ZN(G405));
  OAI21_X1  g1061(.A(new_n1222), .B1(new_n1203), .B2(new_n1234), .ZN(new_n1262));
  NAND3_X1  g1062(.A1(new_n1209), .A2(new_n1202), .A3(new_n1257), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1262), .A2(new_n1263), .ZN(new_n1264));
  XOR2_X1   g1064(.A(new_n1264), .B(new_n1248), .Z(G402));
endmodule


