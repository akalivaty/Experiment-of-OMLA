

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NAND2_X2 U553 ( .A1(n613), .A2(n612), .ZN(n997) );
  NOR2_X1 U554 ( .A1(n737), .A2(n736), .ZN(n756) );
  NOR2_X2 U555 ( .A1(n599), .A2(n598), .ZN(G160) );
  AND2_X1 U556 ( .A1(n534), .A2(n533), .ZN(G164) );
  AND2_X1 U557 ( .A1(n899), .A2(G126), .ZN(n520) );
  XOR2_X1 U558 ( .A(n626), .B(KEYINPUT102), .Z(n521) );
  NAND2_X1 U559 ( .A1(n982), .A2(G29), .ZN(n522) );
  NOR2_X1 U560 ( .A1(n749), .A2(n691), .ZN(n523) );
  XOR2_X1 U561 ( .A(n669), .B(KEYINPUT31), .Z(n524) );
  OR2_X1 U562 ( .A1(n661), .A2(G168), .ZN(n659) );
  INV_X1 U563 ( .A(n652), .ZN(n670) );
  NAND2_X1 U564 ( .A1(n670), .A2(n524), .ZN(n675) );
  XNOR2_X1 U565 ( .A(KEYINPUT106), .B(KEYINPUT32), .ZN(n683) );
  XNOR2_X1 U566 ( .A(n688), .B(n687), .ZN(n738) );
  NOR2_X1 U567 ( .A1(n575), .A2(G651), .ZN(n807) );
  NOR2_X1 U568 ( .A1(n532), .A2(n520), .ZN(n533) );
  NOR2_X1 U569 ( .A1(G2105), .A2(G2104), .ZN(n525) );
  XOR2_X1 U570 ( .A(KEYINPUT17), .B(n525), .Z(n526) );
  XNOR2_X2 U571 ( .A(KEYINPUT66), .B(n526), .ZN(n906) );
  NAND2_X1 U572 ( .A1(G138), .A2(n906), .ZN(n534) );
  NAND2_X1 U573 ( .A1(n531), .A2(G2104), .ZN(n527) );
  XNOR2_X2 U574 ( .A(n527), .B(KEYINPUT65), .ZN(n903) );
  NAND2_X1 U575 ( .A1(n903), .A2(G102), .ZN(n530) );
  AND2_X1 U576 ( .A1(G2105), .A2(G2104), .ZN(n898) );
  NAND2_X1 U577 ( .A1(G114), .A2(n898), .ZN(n528) );
  XOR2_X1 U578 ( .A(KEYINPUT89), .B(n528), .Z(n529) );
  NAND2_X1 U579 ( .A1(n530), .A2(n529), .ZN(n532) );
  INV_X1 U580 ( .A(G2105), .ZN(n531) );
  NOR2_X1 U581 ( .A1(G2104), .A2(n531), .ZN(n899) );
  NOR2_X1 U582 ( .A1(G543), .A2(G651), .ZN(n802) );
  NAND2_X1 U583 ( .A1(n802), .A2(G89), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n535), .B(KEYINPUT4), .ZN(n537) );
  XOR2_X1 U585 ( .A(KEYINPUT0), .B(G543), .Z(n575) );
  INV_X1 U586 ( .A(G651), .ZN(n539) );
  NOR2_X1 U587 ( .A1(n575), .A2(n539), .ZN(n803) );
  NAND2_X1 U588 ( .A1(G76), .A2(n803), .ZN(n536) );
  NAND2_X1 U589 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U590 ( .A(KEYINPUT5), .B(n538), .ZN(n546) );
  NOR2_X1 U591 ( .A1(G543), .A2(n539), .ZN(n540) );
  XOR2_X1 U592 ( .A(KEYINPUT1), .B(n540), .Z(n806) );
  NAND2_X1 U593 ( .A1(G63), .A2(n806), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G51), .A2(n807), .ZN(n541) );
  NAND2_X1 U595 ( .A1(n542), .A2(n541), .ZN(n544) );
  XOR2_X1 U596 ( .A(KEYINPUT76), .B(KEYINPUT6), .Z(n543) );
  XNOR2_X1 U597 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U599 ( .A(KEYINPUT7), .B(n547), .ZN(G168) );
  NAND2_X1 U600 ( .A1(G91), .A2(n802), .ZN(n549) );
  NAND2_X1 U601 ( .A1(G78), .A2(n803), .ZN(n548) );
  NAND2_X1 U602 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U603 ( .A(KEYINPUT71), .B(n550), .ZN(n554) );
  NAND2_X1 U604 ( .A1(G65), .A2(n806), .ZN(n552) );
  NAND2_X1 U605 ( .A1(G53), .A2(n807), .ZN(n551) );
  AND2_X1 U606 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U607 ( .A1(n554), .A2(n553), .ZN(G299) );
  NAND2_X1 U608 ( .A1(G64), .A2(n806), .ZN(n555) );
  XNOR2_X1 U609 ( .A(n555), .B(KEYINPUT68), .ZN(n558) );
  NAND2_X1 U610 ( .A1(G52), .A2(n807), .ZN(n556) );
  XOR2_X1 U611 ( .A(KEYINPUT69), .B(n556), .Z(n557) );
  NAND2_X1 U612 ( .A1(n558), .A2(n557), .ZN(n563) );
  NAND2_X1 U613 ( .A1(G90), .A2(n802), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G77), .A2(n803), .ZN(n559) );
  NAND2_X1 U615 ( .A1(n560), .A2(n559), .ZN(n561) );
  XOR2_X1 U616 ( .A(KEYINPUT9), .B(n561), .Z(n562) );
  NOR2_X1 U617 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U618 ( .A(KEYINPUT70), .B(n564), .ZN(G171) );
  INV_X1 U619 ( .A(G171), .ZN(G301) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G75), .A2(n803), .ZN(n565) );
  XNOR2_X1 U622 ( .A(n565), .B(KEYINPUT84), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n802), .A2(G88), .ZN(n566) );
  NAND2_X1 U624 ( .A1(n567), .A2(n566), .ZN(n571) );
  NAND2_X1 U625 ( .A1(G62), .A2(n806), .ZN(n569) );
  NAND2_X1 U626 ( .A1(G50), .A2(n807), .ZN(n568) );
  NAND2_X1 U627 ( .A1(n569), .A2(n568), .ZN(n570) );
  NOR2_X1 U628 ( .A1(n571), .A2(n570), .ZN(G166) );
  INV_X1 U629 ( .A(G166), .ZN(G303) );
  NAND2_X1 U630 ( .A1(G49), .A2(n807), .ZN(n573) );
  NAND2_X1 U631 ( .A1(G74), .A2(G651), .ZN(n572) );
  NAND2_X1 U632 ( .A1(n573), .A2(n572), .ZN(n574) );
  NOR2_X1 U633 ( .A1(n806), .A2(n574), .ZN(n577) );
  NAND2_X1 U634 ( .A1(n575), .A2(G87), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n577), .A2(n576), .ZN(G288) );
  NAND2_X1 U636 ( .A1(G86), .A2(n802), .ZN(n579) );
  NAND2_X1 U637 ( .A1(G61), .A2(n806), .ZN(n578) );
  NAND2_X1 U638 ( .A1(n579), .A2(n578), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n803), .A2(G73), .ZN(n580) );
  XOR2_X1 U640 ( .A(KEYINPUT2), .B(n580), .Z(n581) );
  NOR2_X1 U641 ( .A1(n582), .A2(n581), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n807), .A2(G48), .ZN(n583) );
  NAND2_X1 U643 ( .A1(n584), .A2(n583), .ZN(G305) );
  NAND2_X1 U644 ( .A1(G85), .A2(n802), .ZN(n586) );
  NAND2_X1 U645 ( .A1(G72), .A2(n803), .ZN(n585) );
  NAND2_X1 U646 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U647 ( .A(KEYINPUT67), .B(n587), .ZN(n591) );
  NAND2_X1 U648 ( .A1(G60), .A2(n806), .ZN(n589) );
  NAND2_X1 U649 ( .A1(G47), .A2(n807), .ZN(n588) );
  AND2_X1 U650 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U651 ( .A1(n591), .A2(n590), .ZN(G290) );
  INV_X1 U652 ( .A(KEYINPUT107), .ZN(n688) );
  NAND2_X1 U653 ( .A1(G125), .A2(n899), .ZN(n592) );
  XNOR2_X1 U654 ( .A(n592), .B(KEYINPUT64), .ZN(n595) );
  NAND2_X1 U655 ( .A1(G101), .A2(n903), .ZN(n593) );
  XOR2_X1 U656 ( .A(KEYINPUT23), .B(n593), .Z(n594) );
  NAND2_X1 U657 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U658 ( .A1(G113), .A2(n898), .ZN(n597) );
  NAND2_X1 U659 ( .A1(G137), .A2(n906), .ZN(n596) );
  NAND2_X1 U660 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U661 ( .A1(G160), .A2(G40), .ZN(n711) );
  INV_X1 U662 ( .A(n711), .ZN(n600) );
  NOR2_X1 U663 ( .A1(G164), .A2(G1384), .ZN(n712) );
  NAND2_X1 U664 ( .A1(n600), .A2(n712), .ZN(n614) );
  NOR2_X1 U665 ( .A1(G2084), .A2(n614), .ZN(n653) );
  NAND2_X1 U666 ( .A1(n653), .A2(G8), .ZN(n674) );
  NAND2_X1 U667 ( .A1(G8), .A2(n614), .ZN(n749) );
  NOR2_X1 U668 ( .A1(G1966), .A2(n749), .ZN(n672) );
  INV_X1 U669 ( .A(n614), .ZN(n647) );
  AND2_X1 U670 ( .A1(n647), .A2(G1996), .ZN(n602) );
  INV_X1 U671 ( .A(KEYINPUT26), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(n617) );
  NAND2_X1 U673 ( .A1(n802), .A2(G81), .ZN(n603) );
  XNOR2_X1 U674 ( .A(n603), .B(KEYINPUT12), .ZN(n605) );
  NAND2_X1 U675 ( .A1(G68), .A2(n803), .ZN(n604) );
  NAND2_X1 U676 ( .A1(n605), .A2(n604), .ZN(n606) );
  XNOR2_X1 U677 ( .A(n606), .B(KEYINPUT13), .ZN(n610) );
  NAND2_X1 U678 ( .A1(G56), .A2(n806), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n607), .B(KEYINPUT72), .ZN(n608) );
  XNOR2_X1 U680 ( .A(KEYINPUT14), .B(n608), .ZN(n609) );
  NAND2_X1 U681 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U682 ( .A(n611), .B(KEYINPUT73), .ZN(n613) );
  NAND2_X1 U683 ( .A1(G43), .A2(n807), .ZN(n612) );
  AND2_X1 U684 ( .A1(n614), .A2(G1341), .ZN(n615) );
  NOR2_X1 U685 ( .A1(n997), .A2(n615), .ZN(n616) );
  AND2_X1 U686 ( .A1(n617), .A2(n616), .ZN(n627) );
  NAND2_X1 U687 ( .A1(G54), .A2(n807), .ZN(n624) );
  NAND2_X1 U688 ( .A1(G92), .A2(n802), .ZN(n619) );
  NAND2_X1 U689 ( .A1(G79), .A2(n803), .ZN(n618) );
  NAND2_X1 U690 ( .A1(n619), .A2(n618), .ZN(n622) );
  NAND2_X1 U691 ( .A1(G66), .A2(n806), .ZN(n620) );
  XNOR2_X1 U692 ( .A(KEYINPUT75), .B(n620), .ZN(n621) );
  NOR2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT15), .ZN(n988) );
  NOR2_X1 U696 ( .A1(n627), .A2(n988), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n627), .A2(n988), .ZN(n631) );
  NOR2_X1 U698 ( .A1(n647), .A2(G1348), .ZN(n629) );
  NOR2_X1 U699 ( .A1(G2067), .A2(n614), .ZN(n628) );
  NOR2_X1 U700 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U701 ( .A1(n631), .A2(n630), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n521), .A2(n632), .ZN(n639) );
  INV_X1 U703 ( .A(G299), .ZN(n816) );
  INV_X1 U704 ( .A(KEYINPUT101), .ZN(n634) );
  NAND2_X1 U705 ( .A1(G2072), .A2(n647), .ZN(n633) );
  XNOR2_X1 U706 ( .A(n634), .B(n633), .ZN(n635) );
  XNOR2_X1 U707 ( .A(n635), .B(KEYINPUT27), .ZN(n637) );
  INV_X1 U708 ( .A(G1956), .ZN(n1011) );
  NOR2_X1 U709 ( .A1(n647), .A2(n1011), .ZN(n636) );
  NOR2_X1 U710 ( .A1(n637), .A2(n636), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n816), .A2(n640), .ZN(n638) );
  NAND2_X1 U712 ( .A1(n639), .A2(n638), .ZN(n644) );
  NOR2_X1 U713 ( .A1(n816), .A2(n640), .ZN(n642) );
  INV_X1 U714 ( .A(KEYINPUT28), .ZN(n641) );
  XNOR2_X1 U715 ( .A(n642), .B(n641), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U717 ( .A(n645), .B(KEYINPUT29), .ZN(n651) );
  XOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .Z(n946) );
  NOR2_X1 U719 ( .A1(n946), .A2(n614), .ZN(n646) );
  XNOR2_X1 U720 ( .A(n646), .B(KEYINPUT100), .ZN(n649) );
  NOR2_X1 U721 ( .A1(n647), .A2(G1961), .ZN(n648) );
  NOR2_X1 U722 ( .A1(n649), .A2(n648), .ZN(n664) );
  NOR2_X1 U723 ( .A1(G301), .A2(n664), .ZN(n650) );
  NOR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n652) );
  INV_X1 U725 ( .A(n653), .ZN(n654) );
  NAND2_X1 U726 ( .A1(G8), .A2(n654), .ZN(n655) );
  NOR2_X1 U727 ( .A1(n672), .A2(n655), .ZN(n657) );
  INV_X1 U728 ( .A(KEYINPUT30), .ZN(n656) );
  XNOR2_X1 U729 ( .A(n657), .B(n656), .ZN(n661) );
  INV_X1 U730 ( .A(KEYINPUT103), .ZN(n658) );
  NAND2_X1 U731 ( .A1(n659), .A2(n658), .ZN(n663) );
  OR2_X1 U732 ( .A1(G168), .A2(n658), .ZN(n660) );
  OR2_X1 U733 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U734 ( .A1(n663), .A2(n662), .ZN(n667) );
  NAND2_X1 U735 ( .A1(G301), .A2(n664), .ZN(n665) );
  XNOR2_X1 U736 ( .A(KEYINPUT104), .B(n665), .ZN(n666) );
  NAND2_X1 U737 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U738 ( .A(n668), .B(KEYINPUT105), .ZN(n669) );
  INV_X1 U739 ( .A(n675), .ZN(n671) );
  NOR2_X1 U740 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U741 ( .A1(n674), .A2(n673), .ZN(n686) );
  NAND2_X1 U742 ( .A1(n675), .A2(G286), .ZN(n682) );
  INV_X1 U743 ( .A(G8), .ZN(n680) );
  NOR2_X1 U744 ( .A1(G1971), .A2(n749), .ZN(n677) );
  NOR2_X1 U745 ( .A1(G2090), .A2(n614), .ZN(n676) );
  NOR2_X1 U746 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U747 ( .A1(n678), .A2(G303), .ZN(n679) );
  OR2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  AND2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U751 ( .A1(n686), .A2(n685), .ZN(n687) );
  NOR2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n729) );
  NOR2_X1 U753 ( .A1(G1971), .A2(G303), .ZN(n689) );
  NOR2_X1 U754 ( .A1(n729), .A2(n689), .ZN(n992) );
  NAND2_X1 U755 ( .A1(n738), .A2(n992), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n690), .B(KEYINPUT108), .ZN(n734) );
  NAND2_X1 U757 ( .A1(G1976), .A2(G288), .ZN(n987) );
  INV_X1 U758 ( .A(n987), .ZN(n691) );
  XOR2_X1 U759 ( .A(G1981), .B(G305), .Z(n1000) );
  NAND2_X1 U760 ( .A1(G95), .A2(n903), .ZN(n693) );
  NAND2_X1 U761 ( .A1(G131), .A2(n906), .ZN(n692) );
  NAND2_X1 U762 ( .A1(n693), .A2(n692), .ZN(n694) );
  XOR2_X1 U763 ( .A(KEYINPUT96), .B(n694), .Z(n696) );
  NAND2_X1 U764 ( .A1(n899), .A2(G119), .ZN(n695) );
  NAND2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U766 ( .A1(G107), .A2(n898), .ZN(n697) );
  XNOR2_X1 U767 ( .A(KEYINPUT95), .B(n697), .ZN(n698) );
  NOR2_X1 U768 ( .A1(n699), .A2(n698), .ZN(n890) );
  INV_X1 U769 ( .A(G1991), .ZN(n940) );
  NOR2_X1 U770 ( .A1(n890), .A2(n940), .ZN(n710) );
  NAND2_X1 U771 ( .A1(G117), .A2(n898), .ZN(n701) );
  NAND2_X1 U772 ( .A1(G129), .A2(n899), .ZN(n700) );
  NAND2_X1 U773 ( .A1(n701), .A2(n700), .ZN(n702) );
  XNOR2_X1 U774 ( .A(KEYINPUT97), .B(n702), .ZN(n708) );
  NAND2_X1 U775 ( .A1(G105), .A2(n903), .ZN(n703) );
  XOR2_X1 U776 ( .A(KEYINPUT38), .B(n703), .Z(n706) );
  NAND2_X1 U777 ( .A1(n906), .A2(G141), .ZN(n704) );
  XOR2_X1 U778 ( .A(KEYINPUT98), .B(n704), .Z(n705) );
  NOR2_X1 U779 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U780 ( .A1(n708), .A2(n707), .ZN(n894) );
  AND2_X1 U781 ( .A1(n894), .A2(G1996), .ZN(n709) );
  NOR2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n968) );
  NOR2_X1 U783 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U784 ( .A(KEYINPUT91), .B(n713), .ZN(n715) );
  NOR2_X1 U785 ( .A1(n968), .A2(n715), .ZN(n763) );
  INV_X1 U786 ( .A(n763), .ZN(n714) );
  AND2_X1 U787 ( .A1(n1000), .A2(n714), .ZN(n728) );
  INV_X1 U788 ( .A(n715), .ZN(n770) );
  NAND2_X1 U789 ( .A1(G140), .A2(n906), .ZN(n716) );
  XNOR2_X1 U790 ( .A(KEYINPUT93), .B(n716), .ZN(n719) );
  NAND2_X1 U791 ( .A1(n903), .A2(G104), .ZN(n717) );
  XOR2_X1 U792 ( .A(KEYINPUT92), .B(n717), .Z(n718) );
  NOR2_X1 U793 ( .A1(n719), .A2(n718), .ZN(n720) );
  XNOR2_X1 U794 ( .A(KEYINPUT34), .B(n720), .ZN(n725) );
  NAND2_X1 U795 ( .A1(G116), .A2(n898), .ZN(n722) );
  NAND2_X1 U796 ( .A1(G128), .A2(n899), .ZN(n721) );
  NAND2_X1 U797 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U798 ( .A(KEYINPUT35), .B(n723), .ZN(n724) );
  NAND2_X1 U799 ( .A1(n725), .A2(n724), .ZN(n726) );
  XNOR2_X1 U800 ( .A(n726), .B(KEYINPUT36), .ZN(n727) );
  XOR2_X1 U801 ( .A(KEYINPUT94), .B(n727), .Z(n895) );
  XNOR2_X1 U802 ( .A(KEYINPUT37), .B(G2067), .ZN(n768) );
  NOR2_X1 U803 ( .A1(n895), .A2(n768), .ZN(n978) );
  NAND2_X1 U804 ( .A1(n770), .A2(n978), .ZN(n766) );
  NAND2_X1 U805 ( .A1(n728), .A2(n766), .ZN(n732) );
  NAND2_X1 U806 ( .A1(n729), .A2(KEYINPUT33), .ZN(n730) );
  NOR2_X1 U807 ( .A1(n749), .A2(n730), .ZN(n731) );
  NOR2_X1 U808 ( .A1(n732), .A2(n731), .ZN(n735) );
  AND2_X1 U809 ( .A1(n523), .A2(n735), .ZN(n733) );
  AND2_X1 U810 ( .A1(n734), .A2(n733), .ZN(n737) );
  AND2_X1 U811 ( .A1(n735), .A2(KEYINPUT33), .ZN(n736) );
  INV_X1 U812 ( .A(n738), .ZN(n741) );
  NAND2_X1 U813 ( .A1(G8), .A2(G166), .ZN(n739) );
  NOR2_X1 U814 ( .A1(G2090), .A2(n739), .ZN(n740) );
  NOR2_X1 U815 ( .A1(n741), .A2(n740), .ZN(n745) );
  INV_X1 U816 ( .A(n749), .ZN(n743) );
  INV_X1 U817 ( .A(n766), .ZN(n742) );
  OR2_X1 U818 ( .A1(n742), .A2(n763), .ZN(n746) );
  OR2_X1 U819 ( .A1(n743), .A2(n746), .ZN(n744) );
  NOR2_X1 U820 ( .A1(n745), .A2(n744), .ZN(n754) );
  INV_X1 U821 ( .A(n746), .ZN(n752) );
  NOR2_X1 U822 ( .A1(G1981), .A2(G305), .ZN(n747) );
  XNOR2_X1 U823 ( .A(n747), .B(KEYINPUT99), .ZN(n748) );
  XNOR2_X1 U824 ( .A(n748), .B(KEYINPUT24), .ZN(n750) );
  NOR2_X1 U825 ( .A1(n750), .A2(n749), .ZN(n751) );
  AND2_X1 U826 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U827 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n759) );
  XNOR2_X1 U829 ( .A(G1986), .B(KEYINPUT90), .ZN(n757) );
  XNOR2_X1 U830 ( .A(n757), .B(G290), .ZN(n985) );
  NAND2_X1 U831 ( .A1(n985), .A2(n770), .ZN(n758) );
  NAND2_X1 U832 ( .A1(n759), .A2(n758), .ZN(n773) );
  NOR2_X1 U833 ( .A1(G1996), .A2(n894), .ZN(n760) );
  XOR2_X1 U834 ( .A(KEYINPUT109), .B(n760), .Z(n973) );
  AND2_X1 U835 ( .A1(n940), .A2(n890), .ZN(n970) );
  NOR2_X1 U836 ( .A1(G1986), .A2(G290), .ZN(n761) );
  NOR2_X1 U837 ( .A1(n970), .A2(n761), .ZN(n762) );
  NOR2_X1 U838 ( .A1(n763), .A2(n762), .ZN(n764) );
  NOR2_X1 U839 ( .A1(n973), .A2(n764), .ZN(n765) );
  XNOR2_X1 U840 ( .A(n765), .B(KEYINPUT39), .ZN(n767) );
  NAND2_X1 U841 ( .A1(n767), .A2(n766), .ZN(n769) );
  NAND2_X1 U842 ( .A1(n895), .A2(n768), .ZN(n979) );
  NAND2_X1 U843 ( .A1(n769), .A2(n979), .ZN(n771) );
  NAND2_X1 U844 ( .A1(n771), .A2(n770), .ZN(n772) );
  NAND2_X1 U845 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U846 ( .A(n774), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U847 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U848 ( .A1(G99), .A2(n903), .ZN(n775) );
  XNOR2_X1 U849 ( .A(n775), .B(KEYINPUT80), .ZN(n782) );
  NAND2_X1 U850 ( .A1(G111), .A2(n898), .ZN(n777) );
  NAND2_X1 U851 ( .A1(G135), .A2(n906), .ZN(n776) );
  NAND2_X1 U852 ( .A1(n777), .A2(n776), .ZN(n780) );
  NAND2_X1 U853 ( .A1(n899), .A2(G123), .ZN(n778) );
  XOR2_X1 U854 ( .A(KEYINPUT18), .B(n778), .Z(n779) );
  NOR2_X1 U855 ( .A1(n780), .A2(n779), .ZN(n781) );
  NAND2_X1 U856 ( .A1(n782), .A2(n781), .ZN(n958) );
  XNOR2_X1 U857 ( .A(G2096), .B(n958), .ZN(n783) );
  OR2_X1 U858 ( .A1(G2100), .A2(n783), .ZN(G156) );
  INV_X1 U859 ( .A(G57), .ZN(G237) );
  NAND2_X1 U860 ( .A1(G7), .A2(G661), .ZN(n785) );
  XNOR2_X1 U861 ( .A(n785), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U862 ( .A(G223), .ZN(n839) );
  NAND2_X1 U863 ( .A1(n839), .A2(G567), .ZN(n786) );
  XOR2_X1 U864 ( .A(KEYINPUT11), .B(n786), .Z(G234) );
  INV_X1 U865 ( .A(G860), .ZN(n846) );
  OR2_X1 U866 ( .A1(n997), .A2(n846), .ZN(G153) );
  INV_X1 U867 ( .A(G868), .ZN(n821) );
  NOR2_X1 U868 ( .A1(n821), .A2(G171), .ZN(n787) );
  XOR2_X1 U869 ( .A(n787), .B(KEYINPUT74), .Z(n789) );
  OR2_X1 U870 ( .A1(G868), .A2(n988), .ZN(n788) );
  NAND2_X1 U871 ( .A1(n789), .A2(n788), .ZN(G284) );
  NAND2_X1 U872 ( .A1(n816), .A2(n821), .ZN(n790) );
  XNOR2_X1 U873 ( .A(n790), .B(KEYINPUT77), .ZN(n792) );
  NOR2_X1 U874 ( .A1(n821), .A2(G286), .ZN(n791) );
  NOR2_X1 U875 ( .A1(n792), .A2(n791), .ZN(G297) );
  NAND2_X1 U876 ( .A1(n846), .A2(G559), .ZN(n793) );
  NAND2_X1 U877 ( .A1(n793), .A2(n988), .ZN(n794) );
  XNOR2_X1 U878 ( .A(n794), .B(KEYINPUT78), .ZN(n795) );
  XNOR2_X1 U879 ( .A(KEYINPUT16), .B(n795), .ZN(G148) );
  NOR2_X1 U880 ( .A1(G868), .A2(n997), .ZN(n796) );
  XOR2_X1 U881 ( .A(KEYINPUT79), .B(n796), .Z(n799) );
  NAND2_X1 U882 ( .A1(G868), .A2(n988), .ZN(n797) );
  NOR2_X1 U883 ( .A1(G559), .A2(n797), .ZN(n798) );
  NOR2_X1 U884 ( .A1(n799), .A2(n798), .ZN(G282) );
  XNOR2_X1 U885 ( .A(n997), .B(KEYINPUT81), .ZN(n801) );
  NAND2_X1 U886 ( .A1(n988), .A2(G559), .ZN(n800) );
  XNOR2_X1 U887 ( .A(n801), .B(n800), .ZN(n847) );
  XNOR2_X1 U888 ( .A(KEYINPUT19), .B(KEYINPUT85), .ZN(n814) );
  NAND2_X1 U889 ( .A1(G93), .A2(n802), .ZN(n805) );
  NAND2_X1 U890 ( .A1(G80), .A2(n803), .ZN(n804) );
  NAND2_X1 U891 ( .A1(n805), .A2(n804), .ZN(n811) );
  NAND2_X1 U892 ( .A1(G67), .A2(n806), .ZN(n809) );
  NAND2_X1 U893 ( .A1(G55), .A2(n807), .ZN(n808) );
  NAND2_X1 U894 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U895 ( .A1(n811), .A2(n810), .ZN(n812) );
  XNOR2_X1 U896 ( .A(KEYINPUT83), .B(n812), .ZN(n845) );
  XOR2_X1 U897 ( .A(G288), .B(n845), .Z(n813) );
  XNOR2_X1 U898 ( .A(n814), .B(n813), .ZN(n815) );
  XNOR2_X1 U899 ( .A(G305), .B(n815), .ZN(n818) );
  XNOR2_X1 U900 ( .A(G166), .B(n816), .ZN(n817) );
  XNOR2_X1 U901 ( .A(n818), .B(n817), .ZN(n819) );
  XNOR2_X1 U902 ( .A(n819), .B(G290), .ZN(n915) );
  XNOR2_X1 U903 ( .A(n847), .B(n915), .ZN(n820) );
  NAND2_X1 U904 ( .A1(n820), .A2(G868), .ZN(n823) );
  NAND2_X1 U905 ( .A1(n821), .A2(n845), .ZN(n822) );
  NAND2_X1 U906 ( .A1(n823), .A2(n822), .ZN(G295) );
  NAND2_X1 U907 ( .A1(G2078), .A2(G2084), .ZN(n825) );
  XOR2_X1 U908 ( .A(KEYINPUT86), .B(KEYINPUT20), .Z(n824) );
  XNOR2_X1 U909 ( .A(n825), .B(n824), .ZN(n826) );
  NAND2_X1 U910 ( .A1(G2090), .A2(n826), .ZN(n827) );
  XNOR2_X1 U911 ( .A(KEYINPUT21), .B(n827), .ZN(n828) );
  NAND2_X1 U912 ( .A1(n828), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U913 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U914 ( .A1(G120), .A2(G69), .ZN(n829) );
  NOR2_X1 U915 ( .A1(G237), .A2(n829), .ZN(n830) );
  XNOR2_X1 U916 ( .A(KEYINPUT88), .B(n830), .ZN(n831) );
  NAND2_X1 U917 ( .A1(n831), .A2(G108), .ZN(n850) );
  NAND2_X1 U918 ( .A1(n850), .A2(G567), .ZN(n837) );
  XOR2_X1 U919 ( .A(KEYINPUT87), .B(KEYINPUT22), .Z(n833) );
  NAND2_X1 U920 ( .A1(G132), .A2(G82), .ZN(n832) );
  XNOR2_X1 U921 ( .A(n833), .B(n832), .ZN(n834) );
  NOR2_X1 U922 ( .A1(n834), .A2(G218), .ZN(n835) );
  NAND2_X1 U923 ( .A1(G96), .A2(n835), .ZN(n851) );
  NAND2_X1 U924 ( .A1(n851), .A2(G2106), .ZN(n836) );
  NAND2_X1 U925 ( .A1(n837), .A2(n836), .ZN(n852) );
  NAND2_X1 U926 ( .A1(G483), .A2(G661), .ZN(n838) );
  NOR2_X1 U927 ( .A1(n852), .A2(n838), .ZN(n844) );
  NAND2_X1 U928 ( .A1(n844), .A2(G36), .ZN(G176) );
  NAND2_X1 U929 ( .A1(G2106), .A2(n839), .ZN(G217) );
  NAND2_X1 U930 ( .A1(G15), .A2(G2), .ZN(n840) );
  XNOR2_X1 U931 ( .A(KEYINPUT111), .B(n840), .ZN(n841) );
  NAND2_X1 U932 ( .A1(n841), .A2(G661), .ZN(n842) );
  XNOR2_X1 U933 ( .A(KEYINPUT112), .B(n842), .ZN(G259) );
  NAND2_X1 U934 ( .A1(G3), .A2(G1), .ZN(n843) );
  NAND2_X1 U935 ( .A1(n844), .A2(n843), .ZN(G188) );
  XNOR2_X1 U937 ( .A(n845), .B(KEYINPUT82), .ZN(n849) );
  NAND2_X1 U938 ( .A1(n847), .A2(n846), .ZN(n848) );
  XNOR2_X1 U939 ( .A(n849), .B(n848), .ZN(G145) );
  INV_X1 U940 ( .A(G132), .ZN(G219) );
  INV_X1 U941 ( .A(G120), .ZN(G236) );
  INV_X1 U942 ( .A(G108), .ZN(G238) );
  INV_X1 U943 ( .A(G96), .ZN(G221) );
  INV_X1 U944 ( .A(G82), .ZN(G220) );
  INV_X1 U945 ( .A(G69), .ZN(G235) );
  NOR2_X1 U946 ( .A1(n851), .A2(n850), .ZN(G325) );
  INV_X1 U947 ( .A(G325), .ZN(G261) );
  INV_X1 U948 ( .A(n852), .ZN(G319) );
  XOR2_X1 U949 ( .A(G1961), .B(G1986), .Z(n854) );
  XNOR2_X1 U950 ( .A(G1996), .B(G1991), .ZN(n853) );
  XNOR2_X1 U951 ( .A(n854), .B(n853), .ZN(n864) );
  XOR2_X1 U952 ( .A(G2474), .B(KEYINPUT115), .Z(n856) );
  XNOR2_X1 U953 ( .A(G1956), .B(KEYINPUT114), .ZN(n855) );
  XNOR2_X1 U954 ( .A(n856), .B(n855), .ZN(n860) );
  XOR2_X1 U955 ( .A(G1976), .B(G1981), .Z(n858) );
  XNOR2_X1 U956 ( .A(G1971), .B(G1966), .ZN(n857) );
  XNOR2_X1 U957 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U958 ( .A(n860), .B(n859), .Z(n862) );
  XNOR2_X1 U959 ( .A(KEYINPUT41), .B(KEYINPUT113), .ZN(n861) );
  XNOR2_X1 U960 ( .A(n862), .B(n861), .ZN(n863) );
  XOR2_X1 U961 ( .A(n864), .B(n863), .Z(G229) );
  XOR2_X1 U962 ( .A(G2100), .B(G2096), .Z(n866) );
  XNOR2_X1 U963 ( .A(KEYINPUT42), .B(G2678), .ZN(n865) );
  XNOR2_X1 U964 ( .A(n866), .B(n865), .ZN(n870) );
  XOR2_X1 U965 ( .A(KEYINPUT43), .B(G2072), .Z(n868) );
  XNOR2_X1 U966 ( .A(G2067), .B(G2090), .ZN(n867) );
  XNOR2_X1 U967 ( .A(n868), .B(n867), .ZN(n869) );
  XOR2_X1 U968 ( .A(n870), .B(n869), .Z(n872) );
  XNOR2_X1 U969 ( .A(G2078), .B(G2084), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n872), .B(n871), .ZN(G227) );
  NAND2_X1 U971 ( .A1(G124), .A2(n899), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT44), .ZN(n875) );
  NAND2_X1 U973 ( .A1(n903), .A2(G100), .ZN(n874) );
  NAND2_X1 U974 ( .A1(n875), .A2(n874), .ZN(n879) );
  NAND2_X1 U975 ( .A1(G112), .A2(n898), .ZN(n877) );
  NAND2_X1 U976 ( .A1(G136), .A2(n906), .ZN(n876) );
  NAND2_X1 U977 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U978 ( .A1(n879), .A2(n878), .ZN(G162) );
  XOR2_X1 U979 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n881) );
  XNOR2_X1 U980 ( .A(G162), .B(KEYINPUT118), .ZN(n880) );
  XNOR2_X1 U981 ( .A(n881), .B(n880), .ZN(n893) );
  NAND2_X1 U982 ( .A1(G106), .A2(n903), .ZN(n883) );
  NAND2_X1 U983 ( .A1(G142), .A2(n906), .ZN(n882) );
  NAND2_X1 U984 ( .A1(n883), .A2(n882), .ZN(n884) );
  XNOR2_X1 U985 ( .A(n884), .B(KEYINPUT45), .ZN(n889) );
  NAND2_X1 U986 ( .A1(G118), .A2(n898), .ZN(n886) );
  NAND2_X1 U987 ( .A1(G130), .A2(n899), .ZN(n885) );
  NAND2_X1 U988 ( .A1(n886), .A2(n885), .ZN(n887) );
  XOR2_X1 U989 ( .A(KEYINPUT116), .B(n887), .Z(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n891), .B(n890), .ZN(n892) );
  XOR2_X1 U992 ( .A(n893), .B(n892), .Z(n897) );
  XOR2_X1 U993 ( .A(n895), .B(n894), .Z(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n913) );
  NAND2_X1 U995 ( .A1(G115), .A2(n898), .ZN(n901) );
  NAND2_X1 U996 ( .A1(G127), .A2(n899), .ZN(n900) );
  NAND2_X1 U997 ( .A1(n901), .A2(n900), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n902), .B(KEYINPUT47), .ZN(n905) );
  NAND2_X1 U999 ( .A1(G103), .A2(n903), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(n909) );
  NAND2_X1 U1001 ( .A1(G139), .A2(n906), .ZN(n907) );
  XNOR2_X1 U1002 ( .A(KEYINPUT117), .B(n907), .ZN(n908) );
  NOR2_X1 U1003 ( .A1(n909), .A2(n908), .ZN(n960) );
  XOR2_X1 U1004 ( .A(G160), .B(n960), .Z(n910) );
  XNOR2_X1 U1005 ( .A(n958), .B(n910), .ZN(n911) );
  XOR2_X1 U1006 ( .A(G164), .B(n911), .Z(n912) );
  XNOR2_X1 U1007 ( .A(n913), .B(n912), .ZN(n914) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n914), .ZN(G395) );
  XNOR2_X1 U1009 ( .A(n997), .B(n915), .ZN(n917) );
  XNOR2_X1 U1010 ( .A(G301), .B(n988), .ZN(n916) );
  XNOR2_X1 U1011 ( .A(n917), .B(n916), .ZN(n918) );
  XOR2_X1 U1012 ( .A(G286), .B(n918), .Z(n919) );
  NOR2_X1 U1013 ( .A1(G37), .A2(n919), .ZN(G397) );
  XOR2_X1 U1014 ( .A(G2443), .B(G2427), .Z(n921) );
  XNOR2_X1 U1015 ( .A(G2438), .B(G2454), .ZN(n920) );
  XNOR2_X1 U1016 ( .A(n921), .B(n920), .ZN(n922) );
  XOR2_X1 U1017 ( .A(n922), .B(G2435), .Z(n924) );
  XNOR2_X1 U1018 ( .A(G1348), .B(G1341), .ZN(n923) );
  XNOR2_X1 U1019 ( .A(n924), .B(n923), .ZN(n928) );
  XOR2_X1 U1020 ( .A(G2430), .B(G2446), .Z(n926) );
  XNOR2_X1 U1021 ( .A(KEYINPUT110), .B(G2451), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(n926), .B(n925), .ZN(n927) );
  XOR2_X1 U1023 ( .A(n928), .B(n927), .Z(n929) );
  NAND2_X1 U1024 ( .A1(G14), .A2(n929), .ZN(n935) );
  NAND2_X1 U1025 ( .A1(G319), .A2(n935), .ZN(n932) );
  NOR2_X1 U1026 ( .A1(G229), .A2(G227), .ZN(n930) );
  XNOR2_X1 U1027 ( .A(KEYINPUT49), .B(n930), .ZN(n931) );
  NOR2_X1 U1028 ( .A1(n932), .A2(n931), .ZN(n934) );
  NOR2_X1 U1029 ( .A1(G395), .A2(G397), .ZN(n933) );
  NAND2_X1 U1030 ( .A1(n934), .A2(n933), .ZN(G225) );
  INV_X1 U1031 ( .A(G225), .ZN(G308) );
  INV_X1 U1032 ( .A(n935), .ZN(G401) );
  XNOR2_X1 U1033 ( .A(KEYINPUT55), .B(KEYINPUT121), .ZN(n957) );
  XOR2_X1 U1034 ( .A(KEYINPUT54), .B(G34), .Z(n936) );
  XNOR2_X1 U1035 ( .A(n936), .B(G2084), .ZN(n953) );
  XNOR2_X1 U1036 ( .A(G2090), .B(G35), .ZN(n951) );
  XNOR2_X1 U1037 ( .A(G1996), .B(G32), .ZN(n938) );
  XNOR2_X1 U1038 ( .A(G33), .B(G2072), .ZN(n937) );
  NOR2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n945) );
  XOR2_X1 U1040 ( .A(G2067), .B(G26), .Z(n939) );
  NAND2_X1 U1041 ( .A1(n939), .A2(G28), .ZN(n943) );
  XOR2_X1 U1042 ( .A(G25), .B(n940), .Z(n941) );
  XNOR2_X1 U1043 ( .A(KEYINPUT122), .B(n941), .ZN(n942) );
  NOR2_X1 U1044 ( .A1(n943), .A2(n942), .ZN(n944) );
  NAND2_X1 U1045 ( .A1(n945), .A2(n944), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G27), .B(n946), .ZN(n947) );
  NOR2_X1 U1047 ( .A1(n948), .A2(n947), .ZN(n949) );
  XNOR2_X1 U1048 ( .A(KEYINPUT53), .B(n949), .ZN(n950) );
  NOR2_X1 U1049 ( .A1(n951), .A2(n950), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n953), .A2(n952), .ZN(n955) );
  INV_X1 U1051 ( .A(G29), .ZN(n954) );
  NAND2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1053 ( .A(n957), .B(n956), .ZN(n983) );
  XNOR2_X1 U1054 ( .A(G160), .B(G2084), .ZN(n959) );
  NAND2_X1 U1055 ( .A1(n959), .A2(n958), .ZN(n966) );
  XOR2_X1 U1056 ( .A(G2072), .B(n960), .Z(n962) );
  XOR2_X1 U1057 ( .A(G164), .B(G2078), .Z(n961) );
  NOR2_X1 U1058 ( .A1(n962), .A2(n961), .ZN(n963) );
  XOR2_X1 U1059 ( .A(KEYINPUT50), .B(n963), .Z(n964) );
  XNOR2_X1 U1060 ( .A(KEYINPUT120), .B(n964), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NOR2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n976) );
  XNOR2_X1 U1064 ( .A(G2090), .B(G162), .ZN(n971) );
  XNOR2_X1 U1065 ( .A(n971), .B(KEYINPUT119), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n974) );
  XOR2_X1 U1067 ( .A(KEYINPUT51), .B(n974), .Z(n975) );
  NAND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NOR2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n980) );
  NAND2_X1 U1070 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1071 ( .A(KEYINPUT52), .B(n981), .ZN(n982) );
  NAND2_X1 U1072 ( .A1(n983), .A2(n522), .ZN(n1036) );
  XNOR2_X1 U1073 ( .A(G16), .B(KEYINPUT56), .ZN(n1006) );
  XNOR2_X1 U1074 ( .A(G301), .B(G1961), .ZN(n984) );
  NOR2_X1 U1075 ( .A1(n985), .A2(n984), .ZN(n996) );
  NAND2_X1 U1076 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n987), .A2(n986), .ZN(n994) );
  XOR2_X1 U1078 ( .A(G1348), .B(n988), .Z(n990) );
  XNOR2_X1 U1079 ( .A(G299), .B(G1956), .ZN(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NOR2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n995) );
  NAND2_X1 U1083 ( .A1(n996), .A2(n995), .ZN(n999) );
  XNOR2_X1 U1084 ( .A(G1341), .B(n997), .ZN(n998) );
  NOR2_X1 U1085 ( .A1(n999), .A2(n998), .ZN(n1004) );
  XNOR2_X1 U1086 ( .A(G168), .B(G1966), .ZN(n1001) );
  NAND2_X1 U1087 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  XNOR2_X1 U1088 ( .A(n1002), .B(KEYINPUT57), .ZN(n1003) );
  NAND2_X1 U1089 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NAND2_X1 U1090 ( .A1(n1006), .A2(n1005), .ZN(n1033) );
  XNOR2_X1 U1091 ( .A(KEYINPUT123), .B(G16), .ZN(n1031) );
  XNOR2_X1 U1092 ( .A(G1961), .B(G5), .ZN(n1008) );
  XNOR2_X1 U1093 ( .A(G21), .B(G1966), .ZN(n1007) );
  NOR2_X1 U1094 ( .A1(n1008), .A2(n1007), .ZN(n1020) );
  XOR2_X1 U1095 ( .A(G4), .B(KEYINPUT124), .Z(n1010) );
  XNOR2_X1 U1096 ( .A(G1348), .B(KEYINPUT59), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1010), .B(n1009), .ZN(n1017) );
  XNOR2_X1 U1098 ( .A(G20), .B(n1011), .ZN(n1015) );
  XNOR2_X1 U1099 ( .A(G1341), .B(G19), .ZN(n1013) );
  XNOR2_X1 U1100 ( .A(G1981), .B(G6), .ZN(n1012) );
  NOR2_X1 U1101 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(n1018), .B(KEYINPUT60), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1027) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1022) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1024) );
  XOR2_X1 U1109 ( .A(G1986), .B(G24), .Z(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XNOR2_X1 U1111 ( .A(KEYINPUT58), .B(n1025), .ZN(n1026) );
  NOR2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  XOR2_X1 U1113 ( .A(n1028), .B(KEYINPUT125), .Z(n1029) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1029), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  NAND2_X1 U1116 ( .A1(n1033), .A2(n1032), .ZN(n1034) );
  XNOR2_X1 U1117 ( .A(KEYINPUT126), .B(n1034), .ZN(n1035) );
  NOR2_X1 U1118 ( .A1(n1036), .A2(n1035), .ZN(n1037) );
  NAND2_X1 U1119 ( .A1(n1037), .A2(G11), .ZN(n1038) );
  XNOR2_X1 U1120 ( .A(n1038), .B(KEYINPUT127), .ZN(n1039) );
  XNOR2_X1 U1121 ( .A(KEYINPUT62), .B(n1039), .ZN(G311) );
  INV_X1 U1122 ( .A(G311), .ZN(G150) );
endmodule

