//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:11 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1270, new_n1271, new_n1272,
    new_n1273, new_n1274, new_n1275, new_n1276, new_n1277, new_n1279,
    new_n1280, new_n1281, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1341,
    new_n1342, new_n1343, new_n1344, new_n1345, new_n1346, new_n1347;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G77), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT66), .ZN(G353));
  OAI21_X1  g0011(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0012(.A(G1), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n216), .A2(G13), .ZN(new_n217));
  OAI211_X1 g0017(.A(new_n217), .B(G250), .C1(G257), .C2(G264), .ZN(new_n218));
  XNOR2_X1  g0018(.A(new_n218), .B(KEYINPUT0), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT70), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n216), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n226), .A2(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g0028(.A1(new_n219), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n206), .A2(new_n207), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT68), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT69), .Z(new_n232));
  AND2_X1   g0032(.A1(KEYINPUT67), .A2(G20), .ZN(new_n233));
  NOR2_X1   g0033(.A1(KEYINPUT67), .A2(G20), .ZN(new_n234));
  NOR2_X1   g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND2_X1  g0035(.A1(G1), .A2(G13), .ZN(new_n236));
  NOR2_X1   g0036(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AOI21_X1  g0037(.A(new_n229), .B1(new_n232), .B2(new_n237), .ZN(G361));
  XNOR2_X1  g0038(.A(G238), .B(G244), .ZN(new_n239));
  INV_X1    g0039(.A(G232), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(KEYINPUT2), .B(G226), .Z(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XNOR2_X1  g0047(.A(G50), .B(G68), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT71), .ZN(new_n249));
  XOR2_X1   g0049(.A(G58), .B(G77), .Z(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n252), .B(KEYINPUT72), .ZN(new_n253));
  XNOR2_X1  g0053(.A(G107), .B(G116), .ZN(new_n254));
  XNOR2_X1  g0054(.A(new_n253), .B(new_n254), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n251), .B(new_n255), .ZN(G351));
  AOI21_X1  g0056(.A(new_n236), .B1(G33), .B2(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G274), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n213), .B1(G41), .B2(G45), .ZN(new_n259));
  OR3_X1    g0059(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT73), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g0062(.A(G33), .ZN(new_n263));
  INV_X1    g0063(.A(G41), .ZN(new_n264));
  OAI211_X1 g0064(.A(G1), .B(G13), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  OAI211_X1 g0065(.A(new_n213), .B(KEYINPUT73), .C1(G41), .C2(G45), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G238), .ZN(new_n268));
  OAI21_X1  g0068(.A(new_n260), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(G33), .A2(G97), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n240), .A2(G1698), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n271), .B1(G226), .B2(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT3), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n270), .B1(new_n272), .B2(new_n276), .ZN(new_n277));
  OR2_X1    g0077(.A1(new_n277), .A2(KEYINPUT76), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n265), .B1(new_n277), .B2(KEYINPUT76), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n269), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g0080(.A(new_n280), .B(KEYINPUT13), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT14), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n282), .A2(new_n283), .A3(G169), .ZN(new_n284));
  INV_X1    g0084(.A(G169), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT14), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n281), .A2(G179), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n284), .A2(new_n286), .A3(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(G20), .A2(G33), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n289), .A2(G50), .B1(G20), .B2(new_n202), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n235), .A2(G33), .ZN(new_n291));
  INV_X1    g0091(.A(G77), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n290), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n294), .A2(new_n236), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OR2_X1    g0096(.A1(new_n296), .A2(KEYINPUT11), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(KEYINPUT11), .ZN(new_n298));
  INV_X1    g0098(.A(G13), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G20), .ZN(new_n301));
  OR3_X1    g0101(.A1(new_n301), .A2(KEYINPUT12), .A3(G68), .ZN(new_n302));
  OAI21_X1  g0102(.A(KEYINPUT12), .B1(new_n301), .B2(G68), .ZN(new_n303));
  NOR3_X1   g0103(.A1(new_n299), .A2(new_n214), .A3(G1), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n304), .A2(new_n295), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n202), .B1(new_n213), .B2(G20), .ZN(new_n306));
  AOI22_X1  g0106(.A1(new_n302), .A2(new_n303), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n297), .A2(new_n298), .A3(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n288), .A2(new_n309), .ZN(new_n310));
  AND3_X1   g0110(.A1(new_n273), .A2(new_n275), .A3(G1698), .ZN(new_n311));
  AOI22_X1  g0111(.A1(new_n311), .A2(G223), .B1(G77), .B2(new_n276), .ZN(new_n312));
  XNOR2_X1  g0112(.A(KEYINPUT3), .B(G33), .ZN(new_n313));
  INV_X1    g0113(.A(G1698), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n313), .A2(G222), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n312), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n316), .A2(new_n257), .ZN(new_n317));
  NOR3_X1   g0117(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n262), .A2(new_n265), .A3(new_n266), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n318), .B1(new_n319), .B2(G226), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G200), .ZN(new_n322));
  INV_X1    g0122(.A(G190), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n321), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n295), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n209), .A2(G20), .ZN(new_n327));
  XNOR2_X1  g0127(.A(KEYINPUT8), .B(G58), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n291), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g0129(.A(new_n329), .B1(G150), .B2(new_n289), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n326), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n213), .A2(G20), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n305), .A2(G50), .A3(new_n332), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n333), .B1(G50), .B2(new_n301), .ZN(new_n334));
  OAI21_X1  g0134(.A(KEYINPUT9), .B1(new_n331), .B2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  NOR3_X1   g0136(.A1(new_n331), .A2(KEYINPUT9), .A3(new_n334), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n325), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n338), .A2(KEYINPUT10), .ZN(new_n339));
  INV_X1    g0139(.A(new_n337), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(new_n335), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT10), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n341), .A2(new_n342), .A3(new_n325), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n282), .A2(G200), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n281), .A2(G190), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n345), .A2(new_n308), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n326), .A2(new_n301), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n332), .A2(G77), .ZN(new_n349));
  OAI22_X1  g0149(.A1(new_n348), .A2(new_n349), .B1(G77), .B2(new_n301), .ZN(new_n350));
  OR2_X1    g0150(.A1(KEYINPUT67), .A2(G20), .ZN(new_n351));
  NAND2_X1  g0151(.A1(KEYINPUT67), .A2(G20), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n214), .A2(new_n263), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI221_X1 g0156(.A(new_n354), .B1(new_n355), .B2(new_n328), .C1(new_n291), .C2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n350), .B1(new_n357), .B2(new_n295), .ZN(new_n358));
  AOI21_X1  g0158(.A(new_n318), .B1(new_n319), .B2(G244), .ZN(new_n359));
  NAND4_X1  g0159(.A1(new_n273), .A2(new_n275), .A3(G238), .A4(G1698), .ZN(new_n360));
  INV_X1    g0160(.A(G107), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n360), .B1(new_n361), .B2(new_n313), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n273), .A2(new_n275), .A3(G232), .A4(new_n314), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT74), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n313), .A2(KEYINPUT74), .A3(G232), .A4(new_n314), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n362), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n359), .B1(new_n367), .B2(new_n265), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n358), .B1(new_n368), .B2(new_n285), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT75), .ZN(new_n370));
  OAI22_X1  g0170(.A1(new_n369), .A2(new_n370), .B1(G179), .B2(new_n368), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n365), .A2(new_n366), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n311), .A2(G238), .B1(G107), .B2(new_n276), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n265), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g0174(.A(G244), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n260), .B1(new_n267), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n285), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n358), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g0179(.A1(new_n379), .A2(KEYINPUT75), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n371), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n321), .A2(new_n285), .ZN(new_n382));
  OAI21_X1  g0182(.A(new_n382), .B1(G179), .B2(new_n321), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n331), .A2(new_n334), .ZN(new_n384));
  NOR2_X1   g0184(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(G190), .B(new_n359), .C1(new_n367), .C2(new_n265), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n386), .A2(new_n358), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n387), .B1(G200), .B2(new_n368), .ZN(new_n388));
  NOR3_X1   g0188(.A1(new_n381), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  AND4_X1   g0189(.A1(new_n310), .A2(new_n344), .A3(new_n347), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT80), .ZN(new_n391));
  INV_X1    g0191(.A(new_n328), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n332), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n393), .A2(new_n348), .B1(new_n301), .B2(new_n392), .ZN(new_n394));
  NOR2_X1   g0194(.A1(new_n274), .A2(G33), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n263), .A2(KEYINPUT3), .ZN(new_n396));
  OAI21_X1  g0196(.A(KEYINPUT77), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT77), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n273), .A2(new_n275), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(new_n235), .A3(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT7), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n400), .A2(KEYINPUT78), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n276), .A2(KEYINPUT7), .A3(new_n214), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(KEYINPUT78), .B1(new_n400), .B2(new_n401), .ZN(new_n405));
  OAI21_X1  g0205(.A(G68), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(G58), .A2(G68), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n203), .A2(new_n205), .A3(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(G20), .ZN(new_n409));
  INV_X1    g0209(.A(G159), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT79), .B1(new_n355), .B2(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT79), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n289), .A2(new_n412), .A3(G159), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n409), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n406), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n401), .B1(new_n276), .B2(new_n235), .ZN(new_n419));
  AOI211_X1 g0219(.A(KEYINPUT7), .B(G20), .C1(new_n273), .C2(new_n275), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n415), .B1(new_n421), .B2(G68), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n295), .B1(new_n422), .B2(KEYINPUT16), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n394), .B1(new_n418), .B2(new_n424), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n318), .B1(new_n319), .B2(G232), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n313), .A2(G226), .A3(G1698), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n273), .A2(new_n275), .A3(G223), .A4(new_n314), .ZN(new_n428));
  NAND2_X1  g0228(.A1(G33), .A2(G87), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n430), .A2(new_n257), .ZN(new_n431));
  AOI21_X1  g0231(.A(G200), .B1(new_n426), .B2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n426), .A2(new_n431), .A3(new_n323), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT17), .B1(new_n425), .B2(new_n435), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n423), .B1(new_n406), .B2(new_n417), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  AND3_X1   g0238(.A1(new_n426), .A2(new_n431), .A3(new_n323), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(new_n432), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n437), .A2(new_n438), .A3(new_n394), .A4(new_n440), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n391), .B1(new_n436), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n426), .A2(new_n431), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(G169), .ZN(new_n444));
  INV_X1    g0244(.A(G179), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n445), .B2(new_n443), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  NOR3_X1   g0247(.A1(new_n425), .A2(KEYINPUT18), .A3(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT18), .ZN(new_n449));
  INV_X1    g0249(.A(new_n394), .ZN(new_n450));
  INV_X1    g0250(.A(new_n417), .ZN(new_n451));
  INV_X1    g0251(.A(KEYINPUT78), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n273), .A2(new_n275), .A3(new_n398), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n398), .B1(new_n273), .B2(new_n275), .ZN(new_n454));
  NOR3_X1   g0254(.A1(new_n453), .A2(new_n454), .A3(new_n353), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n452), .B1(new_n455), .B2(KEYINPUT7), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n456), .A2(new_n403), .A3(new_n402), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n451), .B1(new_n457), .B2(G68), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n450), .B1(new_n458), .B2(new_n423), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n449), .B1(new_n459), .B2(new_n446), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n448), .A2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n450), .B(new_n435), .C1(new_n458), .C2(new_n423), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n462), .A2(new_n438), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n418), .A2(new_n424), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n464), .A2(KEYINPUT17), .A3(new_n450), .A4(new_n435), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT80), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n442), .A2(new_n461), .A3(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n390), .A2(new_n468), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  AND4_X1   g0270(.A1(new_n351), .A2(new_n273), .A3(new_n275), .A4(new_n352), .ZN(new_n471));
  XNOR2_X1  g0271(.A(KEYINPUT84), .B(KEYINPUT19), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n351), .A2(G33), .A3(G97), .A4(new_n352), .ZN(new_n473));
  AOI22_X1  g0273(.A1(new_n471), .A2(G68), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n235), .B(KEYINPUT85), .C1(new_n472), .C2(new_n270), .ZN(new_n475));
  INV_X1    g0275(.A(G87), .ZN(new_n476));
  INV_X1    g0276(.A(G97), .ZN(new_n477));
  NAND3_X1  g0277(.A1(new_n476), .A2(new_n477), .A3(new_n361), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(new_n270), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT19), .ZN(new_n481));
  AND2_X1   g0281(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n481), .A2(KEYINPUT84), .ZN(new_n483));
  OAI21_X1  g0283(.A(new_n480), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(KEYINPUT85), .B1(new_n484), .B2(new_n235), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n474), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(KEYINPUT86), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT86), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n474), .B(new_n488), .C1(new_n479), .C2(new_n485), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n487), .A2(new_n295), .A3(new_n489), .ZN(new_n490));
  INV_X1    g0290(.A(new_n356), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n301), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n305), .B1(G1), .B2(new_n263), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(new_n476), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n375), .A2(G1698), .ZN(new_n497));
  OAI211_X1 g0297(.A(new_n313), .B(new_n497), .C1(G238), .C2(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G116), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n265), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(G45), .ZN(new_n501));
  NOR2_X1   g0301(.A1(new_n501), .A2(G1), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n265), .A2(G274), .A3(new_n502), .ZN(new_n503));
  OAI21_X1  g0303(.A(G250), .B1(new_n501), .B2(G1), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n503), .B1(new_n257), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n500), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n506), .A2(G190), .ZN(new_n507));
  INV_X1    g0307(.A(G200), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n506), .ZN(new_n509));
  NOR3_X1   g0309(.A1(new_n494), .A2(new_n496), .A3(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(new_n495), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n491), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n490), .A2(new_n512), .A3(new_n493), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT87), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n506), .A2(new_n445), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n285), .B1(new_n500), .B2(new_n505), .ZN(new_n516));
  AND2_X1   g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n510), .B1(new_n514), .B2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(G116), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n304), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n520), .B1(new_n495), .B2(new_n519), .ZN(new_n521));
  NAND2_X1  g0321(.A1(G33), .A2(G283), .ZN(new_n522));
  OAI211_X1 g0322(.A(new_n235), .B(new_n522), .C1(G33), .C2(new_n477), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n519), .A2(G20), .ZN(new_n524));
  AND3_X1   g0324(.A1(new_n295), .A2(KEYINPUT88), .A3(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(KEYINPUT88), .B1(new_n295), .B2(new_n524), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n523), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT20), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n523), .B(KEYINPUT20), .C1(new_n525), .C2(new_n526), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n313), .A2(G264), .A3(G1698), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n276), .A2(G303), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n273), .A2(new_n275), .A3(G257), .A4(new_n314), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n532), .A2(new_n533), .A3(new_n534), .ZN(new_n535));
  AND2_X1   g0335(.A1(new_n535), .A2(new_n257), .ZN(new_n536));
  XNOR2_X1  g0336(.A(KEYINPUT5), .B(G41), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n257), .B1(new_n502), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(G270), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n537), .A2(new_n265), .A3(G274), .A4(new_n502), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g0341(.A(G169), .B1(new_n536), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n531), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(new_n531), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n535), .A2(new_n257), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n545), .A2(new_n540), .A3(new_n539), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n546), .A2(new_n445), .ZN(new_n547));
  AOI22_X1  g0347(.A1(new_n543), .A2(KEYINPUT21), .B1(new_n544), .B2(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n549), .B1(new_n531), .B2(new_n542), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n546), .A2(G200), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n531), .B(new_n551), .C1(new_n323), .C2(new_n546), .ZN(new_n552));
  AND3_X1   g0352(.A1(new_n548), .A2(new_n550), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n235), .A2(new_n313), .A3(G87), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n554), .A2(KEYINPUT22), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT22), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n235), .A2(new_n313), .A3(new_n556), .A4(G87), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(KEYINPUT23), .A2(G107), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n353), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(KEYINPUT23), .A2(G107), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n263), .A2(new_n519), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n214), .B1(new_n562), .B2(KEYINPUT23), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n560), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n558), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT90), .ZN(new_n567));
  XOR2_X1   g0367(.A(KEYINPUT89), .B(KEYINPUT24), .Z(new_n568));
  NAND3_X1  g0368(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n568), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n564), .B1(new_n555), .B2(new_n557), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n570), .B1(new_n571), .B2(KEYINPUT90), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n558), .A2(KEYINPUT90), .A3(new_n565), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n295), .B(new_n569), .C1(new_n572), .C2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n313), .A2(G257), .A3(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n313), .A2(G250), .A3(new_n314), .ZN(new_n576));
  NAND2_X1  g0376(.A1(G33), .A2(G294), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(new_n257), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n538), .A2(G264), .ZN(new_n580));
  AND4_X1   g0380(.A1(G190), .A2(new_n579), .A3(new_n540), .A4(new_n580), .ZN(new_n581));
  AOI22_X1  g0381(.A1(new_n578), .A2(new_n257), .B1(G264), .B2(new_n538), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n508), .B1(new_n582), .B2(new_n540), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(KEYINPUT25), .B1(new_n304), .B2(new_n361), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n304), .A2(KEYINPUT25), .A3(new_n361), .ZN(new_n586));
  INV_X1    g0386(.A(new_n586), .ZN(new_n587));
  OAI22_X1  g0387(.A1(new_n495), .A2(new_n361), .B1(new_n585), .B2(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n574), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n289), .A2(G77), .ZN(new_n591));
  XNOR2_X1  g0391(.A(new_n591), .B(KEYINPUT81), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n361), .A2(KEYINPUT6), .A3(G97), .ZN(new_n593));
  XOR2_X1   g0393(.A(G97), .B(G107), .Z(new_n594));
  OAI21_X1  g0394(.A(new_n593), .B1(new_n594), .B2(KEYINPUT6), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n592), .B1(new_n353), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n421), .A2(G107), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n598), .A2(new_n295), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n301), .A2(G97), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n495), .B2(new_n477), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n538), .A2(G257), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(new_n540), .ZN(new_n606));
  INV_X1    g0406(.A(new_n606), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n273), .A2(new_n275), .A3(G244), .A4(new_n314), .ZN(new_n608));
  INV_X1    g0408(.A(KEYINPUT82), .ZN(new_n609));
  OR2_X1    g0409(.A1(new_n609), .A2(KEYINPUT4), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n313), .A2(G244), .A3(new_n610), .A4(new_n314), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n313), .A2(G250), .A3(G1698), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n612), .A2(new_n613), .A3(new_n522), .A4(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT83), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n616), .A3(new_n257), .ZN(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n615), .B2(new_n257), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n445), .B(new_n607), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n615), .A2(new_n257), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n607), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(new_n285), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n604), .A2(new_n620), .A3(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n602), .B1(new_n598), .B2(new_n295), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n606), .B1(new_n257), .B2(new_n615), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G190), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n621), .A2(KEYINPUT83), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n606), .B1(new_n628), .B2(new_n617), .ZN(new_n629));
  OAI211_X1 g0429(.A(new_n625), .B(new_n627), .C1(new_n629), .C2(new_n508), .ZN(new_n630));
  AND3_X1   g0430(.A1(new_n590), .A2(new_n624), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n574), .A2(new_n589), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n582), .A2(new_n540), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G169), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n634), .B1(new_n445), .B2(new_n633), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  AND3_X1   g0436(.A1(new_n553), .A2(new_n631), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n470), .A2(new_n518), .A3(new_n637), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n638), .B(KEYINPUT91), .ZN(G372));
  INV_X1    g0439(.A(new_n385), .ZN(new_n640));
  INV_X1    g0440(.A(new_n461), .ZN(new_n641));
  INV_X1    g0441(.A(new_n347), .ZN(new_n642));
  INV_X1    g0442(.A(new_n381), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n642), .B1(new_n310), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g0444(.A1(new_n463), .A2(KEYINPUT80), .A3(new_n465), .ZN(new_n645));
  AOI21_X1  g0445(.A(KEYINPUT80), .B1(new_n463), .B2(new_n465), .ZN(new_n646));
  NOR2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n641), .B1(new_n644), .B2(new_n647), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n342), .B1(new_n341), .B2(new_n325), .ZN(new_n649));
  AOI211_X1 g0449(.A(KEYINPUT10), .B(new_n324), .C1(new_n340), .C2(new_n335), .ZN(new_n650));
  INV_X1    g0450(.A(KEYINPUT94), .ZN(new_n651));
  NOR3_X1   g0451(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(KEYINPUT94), .B1(new_n339), .B2(new_n343), .ZN(new_n653));
  NOR2_X1   g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n640), .B1(new_n648), .B2(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n516), .A2(KEYINPUT92), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n516), .A2(KEYINPUT92), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n657), .A2(new_n515), .A3(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n513), .A2(KEYINPUT87), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT87), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n326), .B1(new_n486), .B2(KEYINPUT86), .ZN(new_n662));
  AOI21_X1  g0462(.A(new_n492), .B1(new_n662), .B2(new_n489), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n661), .B1(new_n663), .B2(new_n512), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n659), .B1(new_n660), .B2(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(new_n635), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n571), .A2(KEYINPUT90), .ZN(new_n667));
  AOI21_X1  g0467(.A(new_n326), .B1(new_n667), .B2(new_n568), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n566), .A2(new_n567), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n571), .A2(KEYINPUT90), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n669), .A2(new_n670), .A3(new_n570), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n588), .B1(new_n668), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n548), .B(new_n550), .C1(new_n666), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n510), .ZN(new_n674));
  NAND4_X1  g0474(.A1(new_n665), .A2(new_n631), .A3(new_n673), .A4(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT26), .ZN(new_n676));
  INV_X1    g0476(.A(new_n624), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n665), .A2(new_n676), .A3(new_n677), .A4(new_n674), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n665), .A2(KEYINPUT93), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT93), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n514), .A2(new_n680), .A3(new_n659), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n675), .A2(new_n678), .A3(new_n679), .A4(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n676), .B1(new_n518), .B2(new_n677), .ZN(new_n683));
  OR2_X1    g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n470), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n656), .A2(new_n685), .ZN(G369));
  NAND2_X1  g0486(.A1(new_n548), .A2(new_n550), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n235), .A2(new_n300), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(KEYINPUT27), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(G213), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(G343), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n544), .A2(new_n693), .ZN(new_n694));
  MUX2_X1   g0494(.A(new_n687), .B(new_n553), .S(new_n694), .Z(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n632), .A2(new_n693), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n636), .A2(new_n697), .A3(new_n590), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT95), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n636), .A2(new_n697), .A3(KEYINPUT95), .A4(new_n590), .ZN(new_n701));
  INV_X1    g0501(.A(new_n693), .ZN(new_n702));
  OR3_X1    g0502(.A1(new_n636), .A2(KEYINPUT96), .A3(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT96), .B1(new_n636), .B2(new_n702), .ZN(new_n704));
  AOI22_X1  g0504(.A1(new_n700), .A2(new_n701), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n696), .A2(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n636), .A2(new_n693), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n700), .A2(new_n701), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n703), .A2(new_n704), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n687), .A2(new_n702), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n708), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n707), .A2(new_n714), .ZN(G399));
  INV_X1    g0515(.A(new_n217), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G41), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n478), .A2(G116), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n718), .A2(G1), .A3(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n231), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n718), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT28), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n665), .A2(new_n674), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n676), .B1(new_n725), .B2(new_n677), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n517), .B1(new_n660), .B2(new_n664), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n727), .A2(new_n676), .A3(new_n674), .A4(new_n677), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n675), .A2(new_n728), .A3(new_n679), .A4(new_n681), .ZN(new_n729));
  OAI21_X1  g0529(.A(new_n702), .B1(new_n726), .B2(new_n729), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n684), .A2(new_n702), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n732), .B2(KEYINPUT29), .ZN(new_n733));
  INV_X1    g0533(.A(G330), .ZN(new_n734));
  NAND3_X1  g0534(.A1(new_n637), .A2(new_n518), .A3(new_n702), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n547), .A2(new_n626), .A3(new_n506), .A4(new_n582), .ZN(new_n736));
  INV_X1    g0536(.A(KEYINPUT30), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n629), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n506), .A2(G179), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n739), .A2(new_n546), .A3(new_n633), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n736), .A2(new_n737), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n738), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AND3_X1   g0543(.A1(new_n743), .A2(KEYINPUT31), .A3(new_n693), .ZN(new_n744));
  AOI21_X1  g0544(.A(KEYINPUT31), .B1(new_n743), .B2(new_n693), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n734), .B1(new_n735), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n733), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n723), .B1(new_n748), .B2(G1), .ZN(G364));
  NOR2_X1   g0549(.A1(new_n353), .A2(new_n299), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n213), .B1(new_n750), .B2(G45), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n717), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n217), .A2(new_n313), .ZN(new_n754));
  INV_X1    g0554(.A(G355), .ZN(new_n755));
  OAI22_X1  g0555(.A1(new_n754), .A2(new_n755), .B1(G116), .B2(new_n217), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n232), .A2(new_n501), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n453), .A2(new_n454), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(new_n716), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n761), .B1(new_n251), .B2(G45), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n756), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n236), .B1(G20), .B2(new_n285), .ZN(new_n764));
  OR2_X1    g0564(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(KEYINPUT97), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G13), .A2(G33), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n770), .A2(G20), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n753), .B1(new_n763), .B2(new_n773), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n445), .A2(G200), .ZN(new_n775));
  XNOR2_X1  g0575(.A(new_n775), .B(KEYINPUT98), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n214), .A2(new_n323), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(new_n476), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n235), .A2(G190), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n776), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G107), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n313), .ZN(new_n784));
  NOR3_X1   g0584(.A1(G179), .A2(G190), .A3(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n353), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G159), .ZN(new_n788));
  AOI211_X1 g0588(.A(new_n779), .B(new_n784), .C1(KEYINPUT32), .C2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n235), .A2(new_n445), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n323), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n791), .A2(G190), .ZN(new_n793));
  AOI22_X1  g0593(.A1(G50), .A2(new_n792), .B1(new_n793), .B2(G68), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n323), .A2(G200), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n235), .B1(new_n445), .B2(new_n795), .ZN(new_n796));
  XOR2_X1   g0596(.A(new_n796), .B(KEYINPUT99), .Z(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n798), .A2(G97), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n790), .A2(new_n795), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n788), .A2(KEYINPUT32), .B1(new_n800), .B2(new_n201), .ZN(new_n801));
  NOR2_X1   g0601(.A1(G190), .A2(G200), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n790), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n801), .B1(G77), .B2(new_n804), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n789), .A2(new_n794), .A3(new_n799), .A4(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT33), .B(G317), .ZN(new_n807));
  INV_X1    g0607(.A(new_n800), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n793), .A2(new_n807), .B1(new_n808), .B2(G322), .ZN(new_n809));
  XNOR2_X1  g0609(.A(new_n809), .B(KEYINPUT100), .ZN(new_n810));
  INV_X1    g0610(.A(G283), .ZN(new_n811));
  INV_X1    g0611(.A(G303), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n811), .A2(new_n781), .B1(new_n778), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n796), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n813), .B1(G294), .B2(new_n814), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n313), .B1(new_n787), .B2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(G311), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n803), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(G326), .B2(new_n792), .ZN(new_n819));
  NAND3_X1  g0619(.A1(new_n810), .A2(new_n815), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n768), .B1(new_n806), .B2(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n774), .A2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n695), .B2(new_n772), .ZN(new_n823));
  INV_X1    g0623(.A(new_n753), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n696), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n695), .A2(G330), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n823), .B1(new_n825), .B2(new_n826), .ZN(G396));
  OAI21_X1  g0627(.A(new_n388), .B1(new_n371), .B2(new_n380), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n368), .A2(G179), .ZN(new_n829));
  AOI21_X1  g0629(.A(new_n829), .B1(new_n379), .B2(KEYINPUT75), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n369), .A2(new_n370), .ZN(new_n831));
  AOI21_X1  g0631(.A(KEYINPUT104), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n702), .A2(new_n358), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n828), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n833), .ZN(new_n835));
  AOI211_X1 g0635(.A(KEYINPUT104), .B(new_n835), .C1(new_n830), .C2(new_n831), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT105), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n381), .B2(KEYINPUT104), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n832), .A2(new_n833), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT105), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n838), .A2(new_n839), .A3(new_n840), .A4(new_n828), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n769), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n768), .A2(new_n770), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n753), .B1(new_n845), .B2(G77), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n276), .B1(new_n786), .B2(new_n817), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n781), .A2(new_n476), .ZN(new_n848));
  AOI211_X1 g0648(.A(new_n847), .B(new_n848), .C1(G303), .C2(new_n792), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT101), .B(G283), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n793), .A2(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n778), .A2(new_n361), .B1(new_n803), .B2(new_n519), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(G294), .B2(new_n808), .ZN(new_n854));
  NAND4_X1  g0654(.A1(new_n799), .A2(new_n849), .A3(new_n852), .A4(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G137), .A2(new_n792), .B1(new_n793), .B2(G150), .ZN(new_n856));
  XOR2_X1   g0656(.A(new_n856), .B(KEYINPUT102), .Z(new_n857));
  AOI22_X1  g0657(.A1(new_n804), .A2(G159), .B1(new_n808), .B2(G143), .ZN(new_n858));
  XOR2_X1   g0658(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n859));
  NAND3_X1  g0659(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n781), .A2(new_n202), .ZN(new_n861));
  INV_X1    g0661(.A(G132), .ZN(new_n862));
  OAI221_X1 g0662(.A(new_n759), .B1(new_n862), .B2(new_n786), .C1(new_n778), .C2(new_n207), .ZN(new_n863));
  AOI211_X1 g0663(.A(new_n861), .B(new_n863), .C1(G58), .C2(new_n814), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n860), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n859), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n855), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n846), .B1(new_n867), .B2(new_n767), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n844), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n732), .A2(new_n843), .ZN(new_n870));
  OAI211_X1 g0670(.A(new_n842), .B(new_n702), .C1(new_n682), .C2(new_n683), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n870), .A2(new_n747), .A3(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT106), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT106), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  NAND4_X1  g0676(.A1(new_n874), .A2(KEYINPUT107), .A3(new_n824), .A4(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n870), .A2(new_n871), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n735), .A2(new_n746), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(G330), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n877), .A2(new_n881), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n753), .B1(new_n873), .B2(KEYINPUT106), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT107), .B1(new_n883), .B2(new_n876), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n869), .B1(new_n882), .B2(new_n884), .ZN(G384));
  OR2_X1    g0685(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n595), .A2(KEYINPUT35), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n886), .A2(G116), .A3(new_n237), .A4(new_n887), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n888), .B(KEYINPUT36), .Z(new_n889));
  NAND3_X1  g0689(.A1(new_n231), .A2(G77), .A3(new_n407), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n890), .B1(G50), .B2(new_n202), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n213), .A2(G13), .ZN(new_n892));
  AOI21_X1  g0692(.A(new_n889), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n418), .A2(new_n295), .ZN(new_n894));
  INV_X1    g0694(.A(new_n415), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT16), .B1(new_n406), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n450), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(new_n691), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n406), .A2(new_n895), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n416), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n326), .B1(new_n406), .B2(new_n417), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n394), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n462), .B1(new_n904), .B2(new_n691), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n904), .A2(new_n447), .ZN(new_n906));
  OAI21_X1  g0706(.A(KEYINPUT37), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n425), .A2(new_n691), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT37), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n459), .A2(new_n446), .ZN(new_n911));
  NAND4_X1  g0711(.A1(new_n909), .A2(new_n910), .A3(new_n911), .A4(new_n462), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n467), .A2(new_n900), .B1(new_n907), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(KEYINPUT109), .B1(new_n913), .B2(KEYINPUT38), .ZN(new_n914));
  INV_X1    g0714(.A(KEYINPUT109), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT38), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n899), .B1(new_n647), .B2(new_n461), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n911), .A2(new_n462), .ZN(new_n918));
  NOR3_X1   g0718(.A1(new_n918), .A2(KEYINPUT37), .A3(new_n908), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n899), .B(new_n462), .C1(new_n447), .C2(new_n904), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n919), .B1(KEYINPUT37), .B2(new_n920), .ZN(new_n921));
  OAI211_X1 g0721(.A(new_n915), .B(new_n916), .C1(new_n917), .C2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n916), .B1(new_n907), .B2(new_n912), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n467), .A2(new_n900), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n923), .A2(new_n924), .A3(KEYINPUT108), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT108), .B1(new_n923), .B2(new_n924), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n914), .B(new_n922), .C1(new_n925), .C2(new_n926), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n310), .B(new_n347), .C1(new_n308), .C2(new_n702), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n309), .B(new_n693), .C1(new_n642), .C2(new_n288), .ZN(new_n929));
  AND2_X1   g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n879), .ZN(new_n931));
  NOR3_X1   g0731(.A1(new_n930), .A2(new_n931), .A3(new_n843), .ZN(new_n932));
  AOI21_X1  g0732(.A(KEYINPUT40), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n923), .A2(new_n924), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n463), .A2(new_n465), .A3(KEYINPUT110), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n461), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g0736(.A(KEYINPUT110), .B1(new_n463), .B2(new_n465), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n908), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(KEYINPUT37), .B1(new_n918), .B2(new_n908), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n912), .A2(new_n939), .ZN(new_n940));
  AOI21_X1  g0740(.A(KEYINPUT38), .B1(new_n938), .B2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n934), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n928), .A2(new_n929), .ZN(new_n944));
  NAND4_X1  g0744(.A1(new_n944), .A2(new_n879), .A3(KEYINPUT40), .A4(new_n842), .ZN(new_n945));
  INV_X1    g0745(.A(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n933), .B1(new_n943), .B2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n469), .A2(new_n931), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n734), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n949), .B1(new_n947), .B2(new_n948), .ZN(new_n950));
  XOR2_X1   g0750(.A(new_n950), .B(KEYINPUT111), .Z(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n643), .A2(new_n693), .ZN(new_n953));
  INV_X1    g0753(.A(new_n953), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n930), .B1(new_n871), .B2(new_n954), .ZN(new_n955));
  AOI22_X1  g0755(.A1(new_n927), .A2(new_n955), .B1(new_n641), .B2(new_n691), .ZN(new_n956));
  NOR3_X1   g0756(.A1(new_n934), .A2(new_n941), .A3(KEYINPUT39), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n957), .B1(new_n927), .B2(KEYINPUT39), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n288), .A2(new_n309), .A3(new_n702), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n655), .B1(new_n733), .B2(new_n470), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n960), .B(new_n961), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(new_n962), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n951), .A2(new_n964), .B1(new_n213), .B2(new_n750), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n893), .B1(new_n963), .B2(new_n965), .ZN(G367));
  AND2_X1   g0766(.A1(new_n681), .A2(new_n679), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n693), .B1(new_n494), .B2(new_n496), .ZN(new_n968));
  MUX2_X1   g0768(.A(new_n967), .B(new_n724), .S(new_n968), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(new_n771), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n761), .A2(new_n246), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n773), .B1(new_n716), .B2(new_n491), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n824), .B1(new_n971), .B2(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n782), .A2(G97), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n974), .B1(new_n812), .B2(new_n800), .C1(new_n803), .C2(new_n850), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n759), .B1(G317), .B2(new_n787), .ZN(new_n976));
  INV_X1    g0776(.A(new_n793), .ZN(new_n977));
  INV_X1    g0777(.A(G294), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n976), .B1(new_n361), .B2(new_n796), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n975), .B(new_n979), .C1(G311), .C2(new_n792), .ZN(new_n980));
  INV_X1    g0780(.A(new_n778), .ZN(new_n981));
  AOI21_X1  g0781(.A(KEYINPUT113), .B1(new_n981), .B2(G116), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n982), .B(KEYINPUT46), .ZN(new_n983));
  INV_X1    g0783(.A(G137), .ZN(new_n984));
  INV_X1    g0784(.A(G150), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n313), .B1(new_n984), .B2(new_n786), .C1(new_n800), .C2(new_n985), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n977), .A2(new_n410), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n986), .B(new_n987), .C1(G143), .C2(new_n792), .ZN(new_n988));
  NOR2_X1   g0788(.A1(new_n781), .A2(new_n292), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G58), .B2(new_n981), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(new_n207), .B2(new_n803), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(G68), .B2(new_n798), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n980), .A2(new_n983), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n993), .A2(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n767), .ZN(new_n996));
  OAI211_X1 g0796(.A(new_n970), .B(new_n973), .C1(new_n994), .C2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT44), .ZN(new_n998));
  INV_X1    g0798(.A(new_n630), .ZN(new_n999));
  NOR2_X1   g0799(.A1(new_n999), .A2(new_n677), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n604), .A2(new_n693), .ZN(new_n1001));
  AOI22_X1  g0801(.A1(new_n1000), .A2(new_n1001), .B1(new_n677), .B2(new_n693), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n998), .B1(new_n714), .B2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n705), .A2(new_n712), .ZN(new_n1005));
  OAI211_X1 g0805(.A(KEYINPUT44), .B(new_n1002), .C1(new_n1005), .C2(new_n708), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n714), .A2(KEYINPUT45), .A3(new_n1003), .ZN(new_n1007));
  INV_X1    g0807(.A(new_n708), .ZN(new_n1008));
  OAI211_X1 g0808(.A(new_n1008), .B(new_n1003), .C1(new_n705), .C2(new_n712), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1004), .A2(new_n1006), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT112), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n707), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1007), .A2(new_n1011), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1017), .A2(KEYINPUT112), .A3(new_n706), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n711), .A2(new_n713), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n1019), .A2(new_n1005), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(new_n696), .ZN(new_n1021));
  NAND4_X1  g0821(.A1(new_n1014), .A2(new_n1018), .A3(new_n748), .A4(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n748), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n717), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n752), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(KEYINPUT43), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n969), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g0828(.A(new_n624), .B1(new_n636), .B2(new_n999), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1029), .A2(new_n702), .ZN(new_n1030));
  INV_X1    g0830(.A(new_n1030), .ZN(new_n1031));
  NOR3_X1   g0831(.A1(new_n705), .A2(new_n712), .A3(new_n1002), .ZN(new_n1032));
  INV_X1    g0832(.A(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1031), .B1(new_n1033), .B2(KEYINPUT42), .ZN(new_n1034));
  INV_X1    g0834(.A(KEYINPUT42), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1032), .A2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1028), .B1(new_n1034), .B2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n969), .A2(new_n1027), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1034), .A2(new_n1027), .A3(new_n969), .A4(new_n1036), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g0841(.A1(new_n707), .A2(new_n1002), .ZN(new_n1042));
  INV_X1    g0842(.A(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g0843(.A(new_n1041), .B(new_n1043), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n997), .B1(new_n1026), .B2(new_n1044), .ZN(G387));
  NAND2_X1  g0845(.A1(new_n705), .A2(new_n771), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n754), .A2(new_n719), .B1(G107), .B2(new_n217), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n243), .A2(new_n501), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT114), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n328), .A2(G50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT50), .ZN(new_n1051));
  INV_X1    g0851(.A(new_n719), .ZN(new_n1052));
  AOI211_X1 g0852(.A(G45), .B(new_n1052), .C1(G68), .C2(G77), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n761), .B1(new_n1051), .B2(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1047), .B1(new_n1049), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n753), .B1(new_n1055), .B2(new_n773), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n981), .A2(G77), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n758), .B1(G150), .B2(new_n787), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n974), .A2(new_n1057), .A3(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(new_n1059), .B(KEYINPUT115), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n804), .A2(G68), .B1(new_n808), .B2(G50), .ZN(new_n1061));
  OAI21_X1  g0861(.A(new_n1061), .B1(new_n328), .B2(new_n977), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n1062), .B1(G159), .B2(new_n792), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n798), .A2(new_n491), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n759), .B1(G326), .B2(new_n787), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n804), .A2(G303), .B1(new_n808), .B2(G317), .ZN(new_n1067));
  INV_X1    g0867(.A(G322), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n792), .ZN(new_n1069));
  OAI221_X1 g0869(.A(new_n1067), .B1(new_n977), .B2(new_n817), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT48), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(new_n981), .A2(G294), .B1(new_n814), .B2(new_n851), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n1072), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(KEYINPUT49), .ZN(new_n1076));
  OAI221_X1 g0876(.A(new_n1066), .B1(new_n519), .B2(new_n781), .C1(new_n1075), .C2(new_n1076), .ZN(new_n1077));
  AND2_X1   g0877(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1065), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n1056), .B1(new_n1079), .B2(new_n767), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n1021), .A2(new_n752), .B1(new_n1046), .B2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n748), .A2(new_n1021), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n717), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n748), .A2(new_n1021), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1081), .B1(new_n1083), .B2(new_n1084), .ZN(G393));
  INV_X1    g0885(.A(KEYINPUT116), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n706), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n707), .A2(KEYINPUT116), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n1017), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1012), .A2(new_n1086), .A3(new_n706), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1082), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1022), .A2(new_n717), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n773), .B1(G97), .B2(new_n716), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n255), .A2(new_n760), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n824), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n783), .B(new_n276), .C1(new_n1068), .C2(new_n786), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n981), .A2(new_n851), .B1(new_n804), .B2(G294), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n519), .B2(new_n796), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(G303), .C2(new_n793), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n792), .A2(G317), .B1(new_n808), .B2(G311), .ZN(new_n1100));
  XOR2_X1   g0900(.A(new_n1100), .B(KEYINPUT52), .Z(new_n1101));
  AOI22_X1  g0901(.A1(new_n792), .A2(G150), .B1(new_n808), .B2(G159), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT51), .Z(new_n1103));
  AOI22_X1  g0903(.A1(G68), .A2(new_n981), .B1(new_n804), .B2(new_n392), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n848), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n793), .A2(G50), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n758), .B1(G143), .B2(new_n787), .ZN(new_n1107));
  NAND4_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1108), .B1(G77), .B2(new_n798), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n1099), .A2(new_n1101), .B1(new_n1103), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1095), .B1(new_n1110), .B2(new_n768), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1111), .B1(new_n771), .B2(new_n1002), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n752), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1092), .A2(new_n1114), .ZN(G390));
  NAND2_X1  g0915(.A1(new_n927), .A2(KEYINPUT39), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n957), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n871), .A2(new_n954), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n944), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n959), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1116), .A2(new_n1117), .A3(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n702), .B(new_n842), .C1(new_n726), .C2(new_n729), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n930), .B1(new_n1122), .B2(new_n954), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n959), .B1(new_n934), .B2(new_n941), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1121), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n747), .A2(new_n842), .A3(new_n944), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n944), .B1(new_n747), .B2(new_n842), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1118), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n930), .B1(new_n880), .B2(new_n843), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1133), .A2(new_n954), .A3(new_n1128), .A4(new_n1122), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1132), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n470), .A2(new_n747), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1135), .A2(new_n961), .A3(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1121), .A2(new_n1128), .A3(new_n1126), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1130), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI211_X1 g0940(.A(new_n1129), .B(new_n1125), .C1(new_n958), .C2(new_n1120), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1128), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1137), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n1140), .A2(new_n1143), .A3(new_n717), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n861), .B1(G116), .B2(new_n808), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1145), .B1(new_n477), .B2(new_n803), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(G77), .B2(new_n798), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n276), .B1(new_n978), .B2(new_n786), .C1(new_n778), .C2(new_n476), .ZN(new_n1148));
  NOR2_X1   g0948(.A1(new_n1069), .A2(new_n811), .ZN(new_n1149));
  AOI211_X1 g0949(.A(new_n1148), .B(new_n1149), .C1(G107), .C2(new_n793), .ZN(new_n1150));
  INV_X1    g0950(.A(G128), .ZN(new_n1151));
  OAI22_X1  g0951(.A1(new_n1151), .A2(new_n1069), .B1(new_n977), .B2(new_n984), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n276), .B1(new_n787), .B2(G125), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1153), .B1(new_n862), .B2(new_n800), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT54), .B(G143), .ZN(new_n1155));
  OAI22_X1  g0955(.A1(new_n781), .A2(new_n207), .B1(new_n803), .B2(new_n1155), .ZN(new_n1156));
  NOR3_X1   g0956(.A1(new_n1152), .A2(new_n1154), .A3(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT53), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n1158), .B1(new_n778), .B2(new_n985), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n981), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n798), .A2(G159), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1147), .A2(new_n1150), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  OAI221_X1 g0962(.A(new_n753), .B1(new_n392), .B2(new_n845), .C1(new_n1162), .C2(new_n768), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n958), .B2(new_n769), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1141), .A2(new_n1142), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1164), .B1(new_n1165), .B2(new_n752), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT117), .ZN(new_n1167));
  NAND3_X1  g0967(.A1(new_n1144), .A2(new_n1166), .A3(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1144), .B2(new_n1166), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(G378));
  INV_X1    g0971(.A(KEYINPUT57), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n733), .A2(new_n470), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1173), .A2(new_n656), .A3(new_n1136), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(new_n1165), .B2(new_n1138), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n384), .A2(new_n691), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n654), .B2(new_n385), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n651), .B1(new_n649), .B2(new_n650), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n339), .A2(new_n343), .A3(KEYINPUT94), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1176), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n640), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n1182), .A3(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1181), .B1(new_n1180), .B2(new_n640), .ZN(new_n1186));
  AOI211_X1 g0986(.A(new_n385), .B(new_n1176), .C1(new_n1178), .C2(new_n1179), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n927), .A2(new_n932), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT40), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  OAI21_X1  g0992(.A(G330), .B1(new_n942), .B2(new_n945), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1189), .B1(new_n1192), .B2(new_n1194), .ZN(new_n1195));
  AND2_X1   g0995(.A1(new_n1184), .A2(new_n1188), .ZN(new_n1196));
  NOR3_X1   g0996(.A1(new_n933), .A2(new_n1196), .A3(new_n1193), .ZN(new_n1197));
  NOR3_X1   g0997(.A1(new_n1195), .A2(new_n1197), .A3(new_n960), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1192), .A2(new_n1194), .A3(new_n1189), .ZN(new_n1199));
  OAI21_X1  g0999(.A(new_n1196), .B1(new_n933), .B2(new_n1193), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n959), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(new_n1199), .A2(new_n1200), .B1(new_n1203), .B2(new_n956), .ZN(new_n1204));
  NOR2_X1   g1004(.A1(new_n1198), .A2(new_n1204), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1172), .B1(new_n1175), .B2(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1174), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1140), .A2(new_n1207), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n960), .B1(new_n1195), .B2(new_n1197), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1199), .A2(new_n1203), .A3(new_n1200), .A4(new_n956), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n1172), .B1(new_n1209), .B2(new_n1210), .ZN(new_n1211));
  AOI21_X1  g1011(.A(new_n718), .B1(new_n1208), .B2(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1206), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1196), .A2(new_n769), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n753), .B1(new_n845), .B2(G50), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n778), .A2(new_n1155), .B1(new_n800), .B2(new_n1151), .ZN(new_n1217));
  XOR2_X1   g1017(.A(new_n1217), .B(KEYINPUT119), .Z(new_n1218));
  AOI22_X1  g1018(.A1(new_n792), .A2(G125), .B1(new_n804), .B2(G137), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1219), .B1(new_n862), .B2(new_n977), .C1(new_n797), .C2(new_n985), .ZN(new_n1220));
  NOR2_X1   g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  XNOR2_X1  g1021(.A(new_n1221), .B(KEYINPUT59), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT120), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT120), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n782), .A2(G159), .ZN(new_n1226));
  AOI211_X1 g1026(.A(G33), .B(G41), .C1(new_n787), .C2(G124), .ZN(new_n1227));
  NAND4_X1  g1027(.A1(new_n1224), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1057), .B1(new_n811), .B2(new_n786), .C1(new_n977), .C2(new_n477), .ZN(new_n1229));
  NOR2_X1   g1029(.A1(new_n797), .A2(new_n202), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n758), .A2(new_n264), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(G107), .B2(new_n808), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n804), .A2(new_n491), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n782), .A2(G58), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1232), .A2(new_n1233), .A3(new_n1234), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1069), .A2(new_n519), .ZN(new_n1236));
  NOR4_X1   g1036(.A1(new_n1229), .A2(new_n1230), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1238));
  OR2_X1    g1038(.A1(new_n1237), .A2(KEYINPUT58), .ZN(new_n1239));
  OAI211_X1 g1039(.A(new_n1231), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1240));
  XOR2_X1   g1040(.A(new_n1240), .B(KEYINPUT118), .Z(new_n1241));
  NAND4_X1  g1041(.A1(new_n1228), .A2(new_n1238), .A3(new_n1239), .A4(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1216), .B1(new_n1242), .B2(new_n767), .ZN(new_n1243));
  AOI22_X1  g1043(.A1(new_n1214), .A2(new_n752), .B1(new_n1215), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1213), .A2(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(KEYINPUT121), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1244), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1248), .B1(new_n1206), .B2(new_n1212), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(KEYINPUT121), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1247), .A2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(G375));
  NAND2_X1  g1052(.A1(new_n930), .A2(new_n769), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n753), .B1(new_n845), .B2(G68), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n313), .B(new_n989), .C1(G303), .C2(new_n787), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n519), .B2(new_n977), .C1(new_n978), .C2(new_n1069), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G97), .A2(new_n981), .B1(new_n804), .B2(G107), .ZN(new_n1257));
  OAI211_X1 g1057(.A(new_n1064), .B(new_n1257), .C1(new_n811), .C2(new_n800), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n758), .B1(G128), .B2(new_n787), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1234), .A2(new_n1259), .ZN(new_n1260));
  OAI221_X1 g1060(.A(new_n1260), .B1(new_n862), .B2(new_n1069), .C1(new_n977), .C2(new_n1155), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(G159), .A2(new_n981), .B1(new_n804), .B2(G150), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n984), .B2(new_n800), .C1(new_n797), .C2(new_n207), .ZN(new_n1263));
  OAI22_X1  g1063(.A1(new_n1256), .A2(new_n1258), .B1(new_n1261), .B2(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1254), .B1(new_n1264), .B2(new_n767), .ZN(new_n1265));
  AOI22_X1  g1065(.A1(new_n1135), .A2(new_n752), .B1(new_n1253), .B2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1207), .A2(new_n1135), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1137), .A2(new_n1025), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1267), .B2(new_n1268), .ZN(G381));
  NOR3_X1   g1069(.A1(G387), .A2(G390), .A3(G381), .ZN(new_n1270));
  OR3_X1    g1070(.A1(G384), .A2(G396), .A3(G393), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1270), .B1(KEYINPUT122), .B2(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(KEYINPUT122), .B2(new_n1271), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT123), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1144), .A2(new_n1274), .A3(new_n1166), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1144), .B2(new_n1166), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  NAND3_X1  g1077(.A1(new_n1273), .A2(new_n1251), .A3(new_n1277), .ZN(G407));
  INV_X1    g1078(.A(G213), .ZN(new_n1279));
  NOR2_X1   g1079(.A1(new_n1279), .A2(G343), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1251), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(G407), .A2(G213), .A3(new_n1281), .ZN(G409));
  INV_X1    g1082(.A(G390), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(G387), .A2(new_n1283), .ZN(new_n1284));
  OAI211_X1 g1084(.A(G390), .B(new_n997), .C1(new_n1026), .C2(new_n1044), .ZN(new_n1285));
  XOR2_X1   g1085(.A(G393), .B(G396), .Z(new_n1286));
  AND4_X1   g1086(.A1(KEYINPUT126), .A2(new_n1284), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT126), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1285), .A2(new_n1288), .ZN(new_n1289));
  AOI22_X1  g1089(.A1(new_n1289), .A2(new_n1286), .B1(new_n1284), .B2(new_n1285), .ZN(new_n1290));
  NOR2_X1   g1090(.A1(new_n1287), .A2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1291), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1174), .A2(KEYINPUT60), .A3(new_n1132), .A4(new_n1134), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1293), .A2(new_n717), .ZN(new_n1294));
  AND2_X1   g1094(.A1(new_n1137), .A2(KEYINPUT60), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1294), .B1(new_n1267), .B2(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n1266), .ZN(new_n1297));
  INV_X1    g1097(.A(G384), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1296), .A2(G384), .A3(new_n1266), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1280), .A2(G2897), .ZN(new_n1301));
  AND3_X1   g1101(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1302));
  AOI21_X1  g1102(.A(new_n1301), .B1(new_n1299), .B2(new_n1300), .ZN(new_n1303));
  NOR2_X1   g1103(.A1(new_n1302), .A2(new_n1303), .ZN(new_n1304));
  INV_X1    g1104(.A(KEYINPUT124), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1214), .A2(new_n1025), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1175), .ZN(new_n1307));
  NAND4_X1  g1107(.A1(new_n1208), .A2(KEYINPUT124), .A3(new_n1025), .A4(new_n1214), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1307), .A2(new_n1244), .A3(new_n1308), .ZN(new_n1309));
  AOI22_X1  g1109(.A1(G378), .A2(new_n1249), .B1(new_n1277), .B2(new_n1309), .ZN(new_n1310));
  OAI21_X1  g1110(.A(new_n1304), .B1(new_n1310), .B2(new_n1280), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT61), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1277), .A2(new_n1309), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1144), .A2(new_n1166), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1315), .A2(KEYINPUT117), .ZN(new_n1316));
  NAND4_X1  g1116(.A1(new_n1213), .A2(new_n1316), .A3(new_n1168), .A4(new_n1244), .ZN(new_n1317));
  AOI211_X1 g1117(.A(new_n1280), .B(new_n1313), .C1(new_n1314), .C2(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1311), .B(new_n1312), .C1(new_n1318), .C2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1314), .A2(new_n1317), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1280), .ZN(new_n1322));
  INV_X1    g1122(.A(new_n1313), .ZN(new_n1323));
  NAND3_X1  g1123(.A1(new_n1321), .A2(new_n1322), .A3(new_n1323), .ZN(new_n1324));
  XNOR2_X1  g1124(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n1325));
  NOR2_X1   g1125(.A1(new_n1324), .A2(new_n1325), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1292), .B1(new_n1320), .B2(new_n1326), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1280), .B1(new_n1314), .B2(new_n1317), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1303), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1299), .A2(new_n1300), .A3(new_n1301), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1331));
  OAI211_X1 g1131(.A(new_n1291), .B(new_n1312), .C1(new_n1328), .C2(new_n1331), .ZN(new_n1332));
  INV_X1    g1132(.A(new_n1332), .ZN(new_n1333));
  OAI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1318), .B2(KEYINPUT63), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1318), .A2(KEYINPUT63), .ZN(new_n1335));
  INV_X1    g1135(.A(KEYINPUT125), .ZN(new_n1336));
  INV_X1    g1136(.A(KEYINPUT63), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1324), .A2(new_n1336), .A3(new_n1337), .ZN(new_n1338));
  NAND4_X1  g1138(.A1(new_n1333), .A2(new_n1334), .A3(new_n1335), .A4(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1327), .A2(new_n1339), .ZN(G405));
  NAND3_X1  g1140(.A1(new_n1247), .A2(new_n1250), .A3(new_n1277), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1341), .A2(new_n1317), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(new_n1323), .ZN(new_n1343));
  NAND3_X1  g1143(.A1(new_n1341), .A2(new_n1317), .A3(new_n1313), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1345), .A2(new_n1292), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1343), .A2(new_n1291), .A3(new_n1344), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(G402));
endmodule


