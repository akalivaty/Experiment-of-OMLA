

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  AND2_X1 U552 ( .A1(n545), .A2(G2104), .ZN(n867) );
  NOR2_X1 U553 ( .A1(G651), .A2(n632), .ZN(n650) );
  NOR2_X2 U554 ( .A1(G1966), .A2(n775), .ZN(n687) );
  AND2_X2 U555 ( .A1(n705), .A2(G8), .ZN(n683) );
  NOR2_X1 U556 ( .A1(n744), .A2(n688), .ZN(n690) );
  NOR2_X1 U557 ( .A1(n953), .A2(n704), .ZN(n703) );
  INV_X1 U558 ( .A(KEYINPUT28), .ZN(n702) );
  INV_X1 U559 ( .A(KEYINPUT29), .ZN(n725) );
  XNOR2_X1 U560 ( .A(n726), .B(n725), .ZN(n729) );
  NAND2_X1 U561 ( .A1(n729), .A2(n728), .ZN(n746) );
  INV_X1 U562 ( .A(n960), .ZN(n753) );
  AND2_X1 U563 ( .A1(n774), .A2(n753), .ZN(n758) );
  AND2_X1 U564 ( .A1(n766), .A2(n765), .ZN(n767) );
  NAND2_X1 U565 ( .A1(n680), .A2(G40), .ZN(n793) );
  NOR2_X1 U566 ( .A1(G2105), .A2(G2104), .ZN(n549) );
  NOR2_X2 U567 ( .A1(G2104), .A2(n545), .ZN(n870) );
  AND2_X1 U568 ( .A1(n828), .A2(n827), .ZN(n829) );
  XOR2_X1 U569 ( .A(G2443), .B(G2446), .Z(n520) );
  XNOR2_X1 U570 ( .A(G2427), .B(G2451), .ZN(n519) );
  XNOR2_X1 U571 ( .A(n520), .B(n519), .ZN(n526) );
  XOR2_X1 U572 ( .A(G2430), .B(G2454), .Z(n522) );
  XNOR2_X1 U573 ( .A(G1348), .B(G1341), .ZN(n521) );
  XNOR2_X1 U574 ( .A(n522), .B(n521), .ZN(n524) );
  XOR2_X1 U575 ( .A(G2435), .B(G2438), .Z(n523) );
  XNOR2_X1 U576 ( .A(n524), .B(n523), .ZN(n525) );
  XOR2_X1 U577 ( .A(n526), .B(n525), .Z(n527) );
  AND2_X1 U578 ( .A1(G14), .A2(n527), .ZN(G401) );
  NOR2_X1 U579 ( .A1(G651), .A2(G543), .ZN(n643) );
  NAND2_X1 U580 ( .A1(G85), .A2(n643), .ZN(n529) );
  XOR2_X1 U581 ( .A(KEYINPUT0), .B(G543), .Z(n632) );
  INV_X1 U582 ( .A(G651), .ZN(n530) );
  NOR2_X1 U583 ( .A1(n632), .A2(n530), .ZN(n646) );
  NAND2_X1 U584 ( .A1(G72), .A2(n646), .ZN(n528) );
  NAND2_X1 U585 ( .A1(n529), .A2(n528), .ZN(n535) );
  NOR2_X1 U586 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n531), .Z(n642) );
  NAND2_X1 U588 ( .A1(G60), .A2(n642), .ZN(n533) );
  NAND2_X1 U589 ( .A1(G47), .A2(n650), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  OR2_X1 U591 ( .A1(n535), .A2(n534), .ZN(G290) );
  NAND2_X1 U592 ( .A1(G64), .A2(n642), .ZN(n537) );
  NAND2_X1 U593 ( .A1(G52), .A2(n650), .ZN(n536) );
  NAND2_X1 U594 ( .A1(n537), .A2(n536), .ZN(n543) );
  NAND2_X1 U595 ( .A1(G90), .A2(n643), .ZN(n539) );
  NAND2_X1 U596 ( .A1(G77), .A2(n646), .ZN(n538) );
  NAND2_X1 U597 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X1 U598 ( .A(KEYINPUT9), .B(n540), .ZN(n541) );
  XNOR2_X1 U599 ( .A(KEYINPUT65), .B(n541), .ZN(n542) );
  NOR2_X1 U600 ( .A1(n543), .A2(n542), .ZN(G171) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G57), .ZN(G237) );
  INV_X1 U603 ( .A(G132), .ZN(G219) );
  INV_X1 U604 ( .A(G82), .ZN(G220) );
  INV_X1 U605 ( .A(G2105), .ZN(n545) );
  NAND2_X1 U606 ( .A1(G125), .A2(n870), .ZN(n544) );
  XNOR2_X1 U607 ( .A(n544), .B(KEYINPUT64), .ZN(n548) );
  NAND2_X1 U608 ( .A1(G101), .A2(n867), .ZN(n546) );
  XOR2_X1 U609 ( .A(KEYINPUT23), .B(n546), .Z(n547) );
  NAND2_X1 U610 ( .A1(n548), .A2(n547), .ZN(n553) );
  AND2_X1 U611 ( .A1(G2105), .A2(G2104), .ZN(n869) );
  NAND2_X1 U612 ( .A1(G113), .A2(n869), .ZN(n551) );
  XOR2_X2 U613 ( .A(KEYINPUT17), .B(n549), .Z(n875) );
  NAND2_X1 U614 ( .A1(G137), .A2(n875), .ZN(n550) );
  NAND2_X1 U615 ( .A1(n551), .A2(n550), .ZN(n552) );
  NOR2_X1 U616 ( .A1(n553), .A2(n552), .ZN(n680) );
  BUF_X1 U617 ( .A(n680), .Z(G160) );
  NAND2_X1 U618 ( .A1(n867), .A2(G102), .ZN(n556) );
  NAND2_X1 U619 ( .A1(G114), .A2(n869), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT77), .B(n554), .Z(n555) );
  NAND2_X1 U621 ( .A1(n556), .A2(n555), .ZN(n560) );
  NAND2_X1 U622 ( .A1(G138), .A2(n875), .ZN(n558) );
  NAND2_X1 U623 ( .A1(G126), .A2(n870), .ZN(n557) );
  NAND2_X1 U624 ( .A1(n558), .A2(n557), .ZN(n559) );
  NOR2_X1 U625 ( .A1(n560), .A2(n559), .ZN(G164) );
  NAND2_X1 U626 ( .A1(G63), .A2(n642), .ZN(n562) );
  NAND2_X1 U627 ( .A1(G51), .A2(n650), .ZN(n561) );
  NAND2_X1 U628 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(KEYINPUT6), .B(n563), .ZN(n570) );
  NAND2_X1 U630 ( .A1(n643), .A2(G89), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n564), .B(KEYINPUT4), .ZN(n566) );
  NAND2_X1 U632 ( .A1(G76), .A2(n646), .ZN(n565) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n567) );
  XNOR2_X1 U634 ( .A(KEYINPUT5), .B(n567), .ZN(n568) );
  XNOR2_X1 U635 ( .A(KEYINPUT69), .B(n568), .ZN(n569) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT7), .B(n571), .Z(G168) );
  XOR2_X1 U638 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U639 ( .A1(G7), .A2(G661), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U641 ( .A(G223), .ZN(n830) );
  NAND2_X1 U642 ( .A1(n830), .A2(G567), .ZN(n573) );
  XOR2_X1 U643 ( .A(KEYINPUT11), .B(n573), .Z(G234) );
  XOR2_X1 U644 ( .A(KEYINPUT66), .B(KEYINPUT14), .Z(n575) );
  NAND2_X1 U645 ( .A1(G56), .A2(n642), .ZN(n574) );
  XNOR2_X1 U646 ( .A(n575), .B(n574), .ZN(n583) );
  NAND2_X1 U647 ( .A1(n643), .A2(G81), .ZN(n576) );
  XNOR2_X1 U648 ( .A(n576), .B(KEYINPUT12), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G68), .A2(n646), .ZN(n577) );
  NAND2_X1 U650 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U651 ( .A(n579), .B(KEYINPUT13), .ZN(n581) );
  NAND2_X1 U652 ( .A1(G43), .A2(n650), .ZN(n580) );
  NAND2_X1 U653 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U654 ( .A1(n583), .A2(n582), .ZN(n950) );
  NAND2_X1 U655 ( .A1(n950), .A2(G860), .ZN(G153) );
  INV_X1 U656 ( .A(G171), .ZN(G301) );
  NAND2_X1 U657 ( .A1(G868), .A2(G301), .ZN(n594) );
  NAND2_X1 U658 ( .A1(G66), .A2(n642), .ZN(n585) );
  NAND2_X1 U659 ( .A1(G92), .A2(n643), .ZN(n584) );
  NAND2_X1 U660 ( .A1(n585), .A2(n584), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n650), .A2(G54), .ZN(n586) );
  XOR2_X1 U662 ( .A(KEYINPUT67), .B(n586), .Z(n588) );
  NAND2_X1 U663 ( .A1(n646), .A2(G79), .ZN(n587) );
  NAND2_X1 U664 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U665 ( .A(KEYINPUT68), .B(n589), .ZN(n590) );
  NOR2_X1 U666 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U667 ( .A(n592), .B(KEYINPUT15), .ZN(n949) );
  INV_X1 U668 ( .A(G868), .ZN(n663) );
  NAND2_X1 U669 ( .A1(n949), .A2(n663), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(G284) );
  NAND2_X1 U671 ( .A1(G65), .A2(n642), .ZN(n596) );
  NAND2_X1 U672 ( .A1(G53), .A2(n650), .ZN(n595) );
  NAND2_X1 U673 ( .A1(n596), .A2(n595), .ZN(n600) );
  NAND2_X1 U674 ( .A1(G91), .A2(n643), .ZN(n598) );
  NAND2_X1 U675 ( .A1(G78), .A2(n646), .ZN(n597) );
  NAND2_X1 U676 ( .A1(n598), .A2(n597), .ZN(n599) );
  NOR2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n953) );
  INV_X1 U678 ( .A(n953), .ZN(G299) );
  NOR2_X1 U679 ( .A1(G286), .A2(n663), .ZN(n602) );
  NOR2_X1 U680 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U681 ( .A1(n602), .A2(n601), .ZN(G297) );
  INV_X1 U682 ( .A(G860), .ZN(n603) );
  NAND2_X1 U683 ( .A1(n603), .A2(G559), .ZN(n604) );
  INV_X1 U684 ( .A(n949), .ZN(n619) );
  NAND2_X1 U685 ( .A1(n604), .A2(n619), .ZN(n605) );
  XNOR2_X1 U686 ( .A(n605), .B(KEYINPUT16), .ZN(G148) );
  INV_X1 U687 ( .A(n950), .ZN(n887) );
  NOR2_X1 U688 ( .A1(G868), .A2(n887), .ZN(n608) );
  NAND2_X1 U689 ( .A1(G868), .A2(n619), .ZN(n606) );
  NOR2_X1 U690 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U691 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U692 ( .A1(G111), .A2(n869), .ZN(n610) );
  NAND2_X1 U693 ( .A1(G99), .A2(n867), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n610), .A2(n609), .ZN(n611) );
  XNOR2_X1 U695 ( .A(KEYINPUT70), .B(n611), .ZN(n616) );
  NAND2_X1 U696 ( .A1(G123), .A2(n870), .ZN(n612) );
  XNOR2_X1 U697 ( .A(n612), .B(KEYINPUT18), .ZN(n614) );
  NAND2_X1 U698 ( .A1(n875), .A2(G135), .ZN(n613) );
  NAND2_X1 U699 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U700 ( .A1(n616), .A2(n615), .ZN(n1008) );
  XOR2_X1 U701 ( .A(G2096), .B(n1008), .Z(n617) );
  NOR2_X1 U702 ( .A1(G2100), .A2(n617), .ZN(n618) );
  XNOR2_X1 U703 ( .A(KEYINPUT71), .B(n618), .ZN(G156) );
  XOR2_X1 U704 ( .A(n950), .B(KEYINPUT72), .Z(n621) );
  NAND2_X1 U705 ( .A1(G559), .A2(n619), .ZN(n620) );
  XNOR2_X1 U706 ( .A(n621), .B(n620), .ZN(n660) );
  NOR2_X1 U707 ( .A1(G860), .A2(n660), .ZN(n628) );
  NAND2_X1 U708 ( .A1(G67), .A2(n642), .ZN(n623) );
  NAND2_X1 U709 ( .A1(G93), .A2(n643), .ZN(n622) );
  NAND2_X1 U710 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U711 ( .A1(G80), .A2(n646), .ZN(n625) );
  NAND2_X1 U712 ( .A1(G55), .A2(n650), .ZN(n624) );
  NAND2_X1 U713 ( .A1(n625), .A2(n624), .ZN(n626) );
  OR2_X1 U714 ( .A1(n627), .A2(n626), .ZN(n662) );
  XOR2_X1 U715 ( .A(n628), .B(n662), .Z(G145) );
  NAND2_X1 U716 ( .A1(G49), .A2(n650), .ZN(n630) );
  NAND2_X1 U717 ( .A1(G74), .A2(G651), .ZN(n629) );
  NAND2_X1 U718 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U719 ( .A1(n642), .A2(n631), .ZN(n634) );
  NAND2_X1 U720 ( .A1(n632), .A2(G87), .ZN(n633) );
  NAND2_X1 U721 ( .A1(n634), .A2(n633), .ZN(G288) );
  NAND2_X1 U722 ( .A1(G75), .A2(n646), .ZN(n636) );
  NAND2_X1 U723 ( .A1(G50), .A2(n650), .ZN(n635) );
  NAND2_X1 U724 ( .A1(n636), .A2(n635), .ZN(n640) );
  NAND2_X1 U725 ( .A1(G62), .A2(n642), .ZN(n638) );
  NAND2_X1 U726 ( .A1(G88), .A2(n643), .ZN(n637) );
  NAND2_X1 U727 ( .A1(n638), .A2(n637), .ZN(n639) );
  NOR2_X1 U728 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U729 ( .A(n641), .B(KEYINPUT73), .ZN(G303) );
  NAND2_X1 U730 ( .A1(G61), .A2(n642), .ZN(n645) );
  NAND2_X1 U731 ( .A1(G86), .A2(n643), .ZN(n644) );
  NAND2_X1 U732 ( .A1(n645), .A2(n644), .ZN(n649) );
  NAND2_X1 U733 ( .A1(n646), .A2(G73), .ZN(n647) );
  XOR2_X1 U734 ( .A(KEYINPUT2), .B(n647), .Z(n648) );
  NOR2_X1 U735 ( .A1(n649), .A2(n648), .ZN(n652) );
  NAND2_X1 U736 ( .A1(n650), .A2(G48), .ZN(n651) );
  NAND2_X1 U737 ( .A1(n652), .A2(n651), .ZN(G305) );
  XNOR2_X1 U738 ( .A(KEYINPUT19), .B(KEYINPUT75), .ZN(n654) );
  XNOR2_X1 U739 ( .A(G288), .B(KEYINPUT74), .ZN(n653) );
  XNOR2_X1 U740 ( .A(n654), .B(n653), .ZN(n657) );
  XNOR2_X1 U741 ( .A(n953), .B(G290), .ZN(n655) );
  XNOR2_X1 U742 ( .A(n655), .B(G303), .ZN(n656) );
  XNOR2_X1 U743 ( .A(n657), .B(n656), .ZN(n659) );
  XOR2_X1 U744 ( .A(G305), .B(n662), .Z(n658) );
  XNOR2_X1 U745 ( .A(n659), .B(n658), .ZN(n886) );
  XNOR2_X1 U746 ( .A(n660), .B(n886), .ZN(n661) );
  NAND2_X1 U747 ( .A1(n661), .A2(G868), .ZN(n665) );
  NAND2_X1 U748 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U749 ( .A1(n665), .A2(n664), .ZN(G295) );
  NAND2_X1 U750 ( .A1(G2078), .A2(G2084), .ZN(n666) );
  XOR2_X1 U751 ( .A(KEYINPUT20), .B(n666), .Z(n667) );
  NAND2_X1 U752 ( .A1(G2090), .A2(n667), .ZN(n668) );
  XNOR2_X1 U753 ( .A(KEYINPUT21), .B(n668), .ZN(n669) );
  NAND2_X1 U754 ( .A1(n669), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U755 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U756 ( .A1(G220), .A2(G219), .ZN(n670) );
  XOR2_X1 U757 ( .A(KEYINPUT22), .B(n670), .Z(n671) );
  NOR2_X1 U758 ( .A1(G218), .A2(n671), .ZN(n672) );
  NAND2_X1 U759 ( .A1(G96), .A2(n672), .ZN(n837) );
  AND2_X1 U760 ( .A1(G2106), .A2(n837), .ZN(n677) );
  NAND2_X1 U761 ( .A1(G69), .A2(G120), .ZN(n673) );
  NOR2_X1 U762 ( .A1(G237), .A2(n673), .ZN(n674) );
  NAND2_X1 U763 ( .A1(G108), .A2(n674), .ZN(n836) );
  NAND2_X1 U764 ( .A1(G567), .A2(n836), .ZN(n675) );
  XOR2_X1 U765 ( .A(KEYINPUT76), .B(n675), .Z(n676) );
  NOR2_X1 U766 ( .A1(n677), .A2(n676), .ZN(G319) );
  INV_X1 U767 ( .A(G319), .ZN(n679) );
  NAND2_X1 U768 ( .A1(G483), .A2(G661), .ZN(n678) );
  NOR2_X1 U769 ( .A1(n679), .A2(n678), .ZN(n835) );
  NAND2_X1 U770 ( .A1(n835), .A2(G36), .ZN(G176) );
  NOR2_X1 U771 ( .A1(G164), .A2(G1384), .ZN(n794) );
  INV_X1 U772 ( .A(KEYINPUT82), .ZN(n681) );
  XNOR2_X1 U773 ( .A(n793), .B(n681), .ZN(n682) );
  NAND2_X1 U774 ( .A1(n794), .A2(n682), .ZN(n705) );
  XNOR2_X2 U775 ( .A(KEYINPUT83), .B(n683), .ZN(n775) );
  NOR2_X1 U776 ( .A1(G1981), .A2(G305), .ZN(n684) );
  XOR2_X1 U777 ( .A(n684), .B(KEYINPUT24), .Z(n685) );
  NOR2_X1 U778 ( .A1(n775), .A2(n685), .ZN(n686) );
  XNOR2_X1 U779 ( .A(KEYINPUT84), .B(n686), .ZN(n771) );
  INV_X1 U780 ( .A(n705), .ZN(n712) );
  INV_X1 U781 ( .A(n712), .ZN(n730) );
  NOR2_X1 U782 ( .A1(G2084), .A2(n730), .ZN(n744) );
  XNOR2_X1 U783 ( .A(n687), .B(KEYINPUT85), .ZN(n748) );
  NAND2_X1 U784 ( .A1(G8), .A2(n748), .ZN(n688) );
  INV_X1 U785 ( .A(KEYINPUT30), .ZN(n689) );
  XNOR2_X1 U786 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U787 ( .A1(G168), .A2(n691), .ZN(n695) );
  INV_X1 U788 ( .A(G1961), .ZN(n921) );
  NAND2_X1 U789 ( .A1(n730), .A2(n921), .ZN(n693) );
  XNOR2_X1 U790 ( .A(G2078), .B(KEYINPUT25), .ZN(n977) );
  NAND2_X1 U791 ( .A1(n712), .A2(n977), .ZN(n692) );
  NAND2_X1 U792 ( .A1(n693), .A2(n692), .ZN(n727) );
  NOR2_X1 U793 ( .A1(G171), .A2(n727), .ZN(n694) );
  NOR2_X2 U794 ( .A1(n695), .A2(n694), .ZN(n696) );
  XOR2_X1 U795 ( .A(KEYINPUT31), .B(n696), .Z(n745) );
  AND2_X1 U796 ( .A1(n712), .A2(G2072), .ZN(n698) );
  XNOR2_X1 U797 ( .A(KEYINPUT27), .B(KEYINPUT86), .ZN(n697) );
  XNOR2_X1 U798 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U799 ( .A1(n705), .A2(G1956), .ZN(n699) );
  NAND2_X1 U800 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U801 ( .A(KEYINPUT87), .B(n701), .ZN(n704) );
  XNOR2_X1 U802 ( .A(n703), .B(n702), .ZN(n724) );
  NAND2_X1 U803 ( .A1(n953), .A2(n704), .ZN(n722) );
  XOR2_X1 U804 ( .A(G1996), .B(KEYINPUT88), .Z(n984) );
  NOR2_X1 U805 ( .A1(n705), .A2(n984), .ZN(n707) );
  XNOR2_X1 U806 ( .A(KEYINPUT26), .B(KEYINPUT89), .ZN(n706) );
  XNOR2_X1 U807 ( .A(n707), .B(n706), .ZN(n709) );
  NAND2_X1 U808 ( .A1(n730), .A2(G1341), .ZN(n708) );
  NAND2_X1 U809 ( .A1(n709), .A2(n708), .ZN(n710) );
  XOR2_X1 U810 ( .A(KEYINPUT90), .B(n710), .Z(n715) );
  NAND2_X1 U811 ( .A1(n715), .A2(n950), .ZN(n711) );
  NAND2_X1 U812 ( .A1(n711), .A2(n949), .ZN(n720) );
  NOR2_X1 U813 ( .A1(n712), .A2(G1348), .ZN(n714) );
  NOR2_X1 U814 ( .A1(G2067), .A2(n730), .ZN(n713) );
  NOR2_X1 U815 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U816 ( .A1(n949), .A2(n887), .ZN(n716) );
  NAND2_X1 U817 ( .A1(n716), .A2(n715), .ZN(n717) );
  NAND2_X1 U818 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U819 ( .A1(n720), .A2(n719), .ZN(n721) );
  NAND2_X1 U820 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U821 ( .A1(n724), .A2(n723), .ZN(n726) );
  NAND2_X1 U822 ( .A1(n727), .A2(G171), .ZN(n728) );
  INV_X1 U823 ( .A(G8), .ZN(n735) );
  NOR2_X1 U824 ( .A1(G1971), .A2(n775), .ZN(n732) );
  NOR2_X1 U825 ( .A1(G2090), .A2(n730), .ZN(n731) );
  NOR2_X1 U826 ( .A1(n732), .A2(n731), .ZN(n733) );
  NAND2_X1 U827 ( .A1(n733), .A2(G303), .ZN(n734) );
  OR2_X1 U828 ( .A1(n735), .A2(n734), .ZN(n737) );
  AND2_X1 U829 ( .A1(n746), .A2(n737), .ZN(n736) );
  NAND2_X1 U830 ( .A1(n745), .A2(n736), .ZN(n741) );
  INV_X1 U831 ( .A(n737), .ZN(n739) );
  AND2_X1 U832 ( .A1(G286), .A2(G8), .ZN(n738) );
  OR2_X1 U833 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U834 ( .A1(n741), .A2(n740), .ZN(n743) );
  XOR2_X1 U835 ( .A(KEYINPUT32), .B(KEYINPUT91), .Z(n742) );
  XNOR2_X1 U836 ( .A(n743), .B(n742), .ZN(n752) );
  NAND2_X1 U837 ( .A1(G8), .A2(n744), .ZN(n750) );
  NAND2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  AND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U840 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U841 ( .A1(n752), .A2(n751), .ZN(n774) );
  NOR2_X1 U842 ( .A1(G1971), .A2(G303), .ZN(n960) );
  NOR2_X1 U843 ( .A1(G288), .A2(G1976), .ZN(n754) );
  XNOR2_X1 U844 ( .A(n754), .B(KEYINPUT92), .ZN(n755) );
  INV_X1 U845 ( .A(n755), .ZN(n963) );
  INV_X1 U846 ( .A(n775), .ZN(n761) );
  NAND2_X1 U847 ( .A1(n755), .A2(n761), .ZN(n756) );
  NAND2_X1 U848 ( .A1(n756), .A2(KEYINPUT33), .ZN(n759) );
  AND2_X1 U849 ( .A1(n963), .A2(n759), .ZN(n757) );
  NAND2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n766) );
  INV_X1 U851 ( .A(n759), .ZN(n764) );
  INV_X1 U852 ( .A(KEYINPUT33), .ZN(n760) );
  NAND2_X1 U853 ( .A1(G1976), .A2(G288), .ZN(n954) );
  AND2_X1 U854 ( .A1(n760), .A2(n954), .ZN(n762) );
  AND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n763) );
  OR2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  XNOR2_X1 U857 ( .A(n767), .B(KEYINPUT93), .ZN(n768) );
  XNOR2_X1 U858 ( .A(G1981), .B(G305), .ZN(n947) );
  NOR2_X1 U859 ( .A1(n768), .A2(n947), .ZN(n769) );
  XNOR2_X1 U860 ( .A(n769), .B(KEYINPUT94), .ZN(n770) );
  NOR2_X1 U861 ( .A1(n771), .A2(n770), .ZN(n817) );
  NOR2_X1 U862 ( .A1(G2090), .A2(G303), .ZN(n772) );
  NAND2_X1 U863 ( .A1(G8), .A2(n772), .ZN(n773) );
  NAND2_X1 U864 ( .A1(n774), .A2(n773), .ZN(n776) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n815) );
  NAND2_X1 U866 ( .A1(G117), .A2(n869), .ZN(n778) );
  NAND2_X1 U867 ( .A1(G129), .A2(n870), .ZN(n777) );
  NAND2_X1 U868 ( .A1(n778), .A2(n777), .ZN(n781) );
  NAND2_X1 U869 ( .A1(n867), .A2(G105), .ZN(n779) );
  XOR2_X1 U870 ( .A(KEYINPUT38), .B(n779), .Z(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n783) );
  NAND2_X1 U872 ( .A1(n875), .A2(G141), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(n855) );
  NOR2_X1 U874 ( .A1(G1996), .A2(n855), .ZN(n1004) );
  NAND2_X1 U875 ( .A1(n855), .A2(G1996), .ZN(n792) );
  NAND2_X1 U876 ( .A1(G95), .A2(n867), .ZN(n785) );
  NAND2_X1 U877 ( .A1(G119), .A2(n870), .ZN(n784) );
  NAND2_X1 U878 ( .A1(n785), .A2(n784), .ZN(n788) );
  NAND2_X1 U879 ( .A1(n869), .A2(G107), .ZN(n786) );
  XOR2_X1 U880 ( .A(KEYINPUT80), .B(n786), .Z(n787) );
  NOR2_X1 U881 ( .A1(n788), .A2(n787), .ZN(n790) );
  NAND2_X1 U882 ( .A1(n875), .A2(G131), .ZN(n789) );
  NAND2_X1 U883 ( .A1(n790), .A2(n789), .ZN(n851) );
  NAND2_X1 U884 ( .A1(G1991), .A2(n851), .ZN(n791) );
  NAND2_X1 U885 ( .A1(n792), .A2(n791), .ZN(n1007) );
  NOR2_X1 U886 ( .A1(n794), .A2(n793), .ZN(n819) );
  AND2_X1 U887 ( .A1(n1007), .A2(n819), .ZN(n820) );
  NOR2_X1 U888 ( .A1(G1991), .A2(n851), .ZN(n1009) );
  NOR2_X1 U889 ( .A1(G1986), .A2(G290), .ZN(n795) );
  XOR2_X1 U890 ( .A(n795), .B(KEYINPUT95), .Z(n796) );
  NOR2_X1 U891 ( .A1(n1009), .A2(n796), .ZN(n797) );
  NOR2_X1 U892 ( .A1(n820), .A2(n797), .ZN(n798) );
  NOR2_X1 U893 ( .A1(n1004), .A2(n798), .ZN(n799) );
  XNOR2_X1 U894 ( .A(KEYINPUT39), .B(n799), .ZN(n811) );
  XOR2_X1 U895 ( .A(KEYINPUT37), .B(G2067), .Z(n812) );
  NAND2_X1 U896 ( .A1(G104), .A2(n867), .ZN(n801) );
  NAND2_X1 U897 ( .A1(G140), .A2(n875), .ZN(n800) );
  NAND2_X1 U898 ( .A1(n801), .A2(n800), .ZN(n802) );
  XNOR2_X1 U899 ( .A(KEYINPUT34), .B(n802), .ZN(n808) );
  NAND2_X1 U900 ( .A1(G116), .A2(n869), .ZN(n804) );
  NAND2_X1 U901 ( .A1(G128), .A2(n870), .ZN(n803) );
  NAND2_X1 U902 ( .A1(n804), .A2(n803), .ZN(n805) );
  XOR2_X1 U903 ( .A(KEYINPUT78), .B(n805), .Z(n806) );
  XNOR2_X1 U904 ( .A(KEYINPUT35), .B(n806), .ZN(n807) );
  NOR2_X1 U905 ( .A1(n808), .A2(n807), .ZN(n809) );
  XOR2_X1 U906 ( .A(KEYINPUT36), .B(n809), .Z(n882) );
  NAND2_X1 U907 ( .A1(n812), .A2(n882), .ZN(n810) );
  XNOR2_X1 U908 ( .A(n810), .B(KEYINPUT79), .ZN(n1026) );
  NAND2_X1 U909 ( .A1(n819), .A2(n1026), .ZN(n823) );
  NAND2_X1 U910 ( .A1(n811), .A2(n823), .ZN(n813) );
  OR2_X1 U911 ( .A1(n882), .A2(n812), .ZN(n1014) );
  NAND2_X1 U912 ( .A1(n813), .A2(n1014), .ZN(n814) );
  NAND2_X1 U913 ( .A1(n814), .A2(n819), .ZN(n818) );
  AND2_X1 U914 ( .A1(n815), .A2(n818), .ZN(n816) );
  NAND2_X1 U915 ( .A1(n817), .A2(n816), .ZN(n828) );
  INV_X1 U916 ( .A(n818), .ZN(n826) );
  XNOR2_X1 U917 ( .A(G1986), .B(G290), .ZN(n959) );
  AND2_X1 U918 ( .A1(n959), .A2(n819), .ZN(n822) );
  XOR2_X1 U919 ( .A(KEYINPUT81), .B(n820), .Z(n821) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n824) );
  AND2_X1 U921 ( .A1(n824), .A2(n823), .ZN(n825) );
  OR2_X1 U922 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n829), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U924 ( .A1(G2106), .A2(n830), .ZN(G217) );
  NAND2_X1 U925 ( .A1(G15), .A2(G2), .ZN(n831) );
  XOR2_X1 U926 ( .A(KEYINPUT96), .B(n831), .Z(n832) );
  NAND2_X1 U927 ( .A1(n832), .A2(G661), .ZN(n833) );
  XOR2_X1 U928 ( .A(KEYINPUT97), .B(n833), .Z(G259) );
  NAND2_X1 U929 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U930 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U932 ( .A(G120), .ZN(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  NOR2_X1 U935 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U936 ( .A(G325), .ZN(G261) );
  NAND2_X1 U937 ( .A1(G124), .A2(n870), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n838), .B(KEYINPUT44), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n839), .B(KEYINPUT102), .ZN(n841) );
  NAND2_X1 U940 ( .A1(G136), .A2(n875), .ZN(n840) );
  NAND2_X1 U941 ( .A1(n841), .A2(n840), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n842), .B(KEYINPUT103), .ZN(n844) );
  NAND2_X1 U943 ( .A1(G112), .A2(n869), .ZN(n843) );
  NAND2_X1 U944 ( .A1(n844), .A2(n843), .ZN(n847) );
  NAND2_X1 U945 ( .A1(n867), .A2(G100), .ZN(n845) );
  XOR2_X1 U946 ( .A(KEYINPUT104), .B(n845), .Z(n846) );
  NOR2_X1 U947 ( .A1(n847), .A2(n846), .ZN(G162) );
  XNOR2_X1 U948 ( .A(n1008), .B(G162), .ZN(n857) );
  XOR2_X1 U949 ( .A(KEYINPUT48), .B(KEYINPUT110), .Z(n849) );
  XNOR2_X1 U950 ( .A(KEYINPUT46), .B(KEYINPUT109), .ZN(n848) );
  XNOR2_X1 U951 ( .A(n849), .B(n848), .ZN(n850) );
  XNOR2_X1 U952 ( .A(n851), .B(n850), .ZN(n853) );
  XNOR2_X1 U953 ( .A(G164), .B(G160), .ZN(n852) );
  XNOR2_X1 U954 ( .A(n853), .B(n852), .ZN(n854) );
  XNOR2_X1 U955 ( .A(n855), .B(n854), .ZN(n856) );
  XNOR2_X1 U956 ( .A(n857), .B(n856), .ZN(n884) );
  NAND2_X1 U957 ( .A1(G118), .A2(n869), .ZN(n866) );
  NAND2_X1 U958 ( .A1(n870), .A2(G130), .ZN(n858) );
  XNOR2_X1 U959 ( .A(KEYINPUT105), .B(n858), .ZN(n864) );
  NAND2_X1 U960 ( .A1(G106), .A2(n867), .ZN(n860) );
  NAND2_X1 U961 ( .A1(G142), .A2(n875), .ZN(n859) );
  NAND2_X1 U962 ( .A1(n860), .A2(n859), .ZN(n861) );
  XOR2_X1 U963 ( .A(KEYINPUT45), .B(n861), .Z(n862) );
  XNOR2_X1 U964 ( .A(KEYINPUT106), .B(n862), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n880) );
  NAND2_X1 U967 ( .A1(n867), .A2(G103), .ZN(n868) );
  XNOR2_X1 U968 ( .A(KEYINPUT107), .B(n868), .ZN(n879) );
  NAND2_X1 U969 ( .A1(G115), .A2(n869), .ZN(n872) );
  NAND2_X1 U970 ( .A1(G127), .A2(n870), .ZN(n871) );
  NAND2_X1 U971 ( .A1(n872), .A2(n871), .ZN(n873) );
  XNOR2_X1 U972 ( .A(n873), .B(KEYINPUT108), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n874), .B(KEYINPUT47), .ZN(n877) );
  NAND2_X1 U974 ( .A1(n875), .A2(G139), .ZN(n876) );
  NAND2_X1 U975 ( .A1(n877), .A2(n876), .ZN(n878) );
  NOR2_X1 U976 ( .A1(n879), .A2(n878), .ZN(n1016) );
  XNOR2_X1 U977 ( .A(n880), .B(n1016), .ZN(n881) );
  XNOR2_X1 U978 ( .A(n882), .B(n881), .ZN(n883) );
  XNOR2_X1 U979 ( .A(n884), .B(n883), .ZN(n885) );
  NOR2_X1 U980 ( .A1(G37), .A2(n885), .ZN(G395) );
  XNOR2_X1 U981 ( .A(n886), .B(n949), .ZN(n888) );
  XNOR2_X1 U982 ( .A(n888), .B(n887), .ZN(n890) );
  XNOR2_X1 U983 ( .A(G286), .B(G171), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n890), .B(n889), .ZN(n891) );
  NOR2_X1 U985 ( .A1(G37), .A2(n891), .ZN(n892) );
  XOR2_X1 U986 ( .A(KEYINPUT111), .B(n892), .Z(G397) );
  XOR2_X1 U987 ( .A(KEYINPUT101), .B(G1981), .Z(n894) );
  XNOR2_X1 U988 ( .A(G1956), .B(G1971), .ZN(n893) );
  XNOR2_X1 U989 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U990 ( .A(n895), .B(KEYINPUT41), .Z(n897) );
  XNOR2_X1 U991 ( .A(G1996), .B(G1991), .ZN(n896) );
  XNOR2_X1 U992 ( .A(n897), .B(n896), .ZN(n901) );
  XOR2_X1 U993 ( .A(G1976), .B(G1961), .Z(n899) );
  XNOR2_X1 U994 ( .A(G1986), .B(G1966), .ZN(n898) );
  XNOR2_X1 U995 ( .A(n899), .B(n898), .ZN(n900) );
  XOR2_X1 U996 ( .A(n901), .B(n900), .Z(n903) );
  XNOR2_X1 U997 ( .A(KEYINPUT100), .B(G2474), .ZN(n902) );
  XNOR2_X1 U998 ( .A(n903), .B(n902), .ZN(G229) );
  XOR2_X1 U999 ( .A(KEYINPUT99), .B(KEYINPUT98), .Z(n905) );
  XNOR2_X1 U1000 ( .A(G2678), .B(KEYINPUT43), .ZN(n904) );
  XNOR2_X1 U1001 ( .A(n905), .B(n904), .ZN(n909) );
  XOR2_X1 U1002 ( .A(KEYINPUT42), .B(G2090), .Z(n907) );
  XNOR2_X1 U1003 ( .A(G2067), .B(G2072), .ZN(n906) );
  XNOR2_X1 U1004 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1005 ( .A(n909), .B(n908), .Z(n911) );
  XNOR2_X1 U1006 ( .A(G2096), .B(G2100), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n913) );
  XOR2_X1 U1008 ( .A(G2078), .B(G2084), .Z(n912) );
  XNOR2_X1 U1009 ( .A(n913), .B(n912), .ZN(G227) );
  NOR2_X1 U1010 ( .A1(G395), .A2(G397), .ZN(n914) );
  XOR2_X1 U1011 ( .A(KEYINPUT113), .B(n914), .Z(n920) );
  NOR2_X1 U1012 ( .A1(G229), .A2(G227), .ZN(n915) );
  XOR2_X1 U1013 ( .A(KEYINPUT49), .B(n915), .Z(n916) );
  NAND2_X1 U1014 ( .A1(G319), .A2(n916), .ZN(n917) );
  NOR2_X1 U1015 ( .A1(G401), .A2(n917), .ZN(n918) );
  XNOR2_X1 U1016 ( .A(KEYINPUT112), .B(n918), .ZN(n919) );
  NAND2_X1 U1017 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1018 ( .A(G225), .ZN(G308) );
  INV_X1 U1019 ( .A(G303), .ZN(G166) );
  INV_X1 U1020 ( .A(G108), .ZN(G238) );
  XNOR2_X1 U1021 ( .A(G5), .B(n921), .ZN(n932) );
  XOR2_X1 U1022 ( .A(G1971), .B(G22), .Z(n924) );
  XOR2_X1 U1023 ( .A(G24), .B(KEYINPUT126), .Z(n922) );
  XNOR2_X1 U1024 ( .A(n922), .B(G1986), .ZN(n923) );
  NAND2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1026 ( .A(KEYINPUT125), .B(G1976), .Z(n925) );
  XNOR2_X1 U1027 ( .A(G23), .B(n925), .ZN(n926) );
  NOR2_X1 U1028 ( .A1(n927), .A2(n926), .ZN(n928) );
  XOR2_X1 U1029 ( .A(KEYINPUT58), .B(n928), .Z(n930) );
  XNOR2_X1 U1030 ( .A(G1966), .B(G21), .ZN(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1032 ( .A1(n932), .A2(n931), .ZN(n943) );
  XNOR2_X1 U1033 ( .A(G1341), .B(G19), .ZN(n934) );
  XNOR2_X1 U1034 ( .A(G6), .B(G1981), .ZN(n933) );
  NOR2_X1 U1035 ( .A1(n934), .A2(n933), .ZN(n940) );
  XOR2_X1 U1036 ( .A(KEYINPUT124), .B(G4), .Z(n936) );
  XNOR2_X1 U1037 ( .A(G1348), .B(KEYINPUT59), .ZN(n935) );
  XNOR2_X1 U1038 ( .A(n936), .B(n935), .ZN(n938) );
  XNOR2_X1 U1039 ( .A(G1956), .B(G20), .ZN(n937) );
  NOR2_X1 U1040 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1041 ( .A1(n940), .A2(n939), .ZN(n941) );
  XNOR2_X1 U1042 ( .A(KEYINPUT60), .B(n941), .ZN(n942) );
  NOR2_X1 U1043 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1044 ( .A(KEYINPUT61), .B(n944), .Z(n945) );
  NOR2_X1 U1045 ( .A1(G16), .A2(n945), .ZN(n1034) );
  XNOR2_X1 U1046 ( .A(G16), .B(KEYINPUT56), .ZN(n974) );
  XOR2_X1 U1047 ( .A(G1966), .B(G168), .Z(n946) );
  NOR2_X1 U1048 ( .A1(n947), .A2(n946), .ZN(n948) );
  XOR2_X1 U1049 ( .A(KEYINPUT57), .B(n948), .Z(n972) );
  XNOR2_X1 U1050 ( .A(G1348), .B(n949), .ZN(n969) );
  XNOR2_X1 U1051 ( .A(n950), .B(G1341), .ZN(n952) );
  NAND2_X1 U1052 ( .A1(G1971), .A2(G303), .ZN(n951) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n957) );
  XNOR2_X1 U1054 ( .A(n953), .B(G1956), .ZN(n955) );
  NAND2_X1 U1055 ( .A1(n955), .A2(n954), .ZN(n956) );
  NOR2_X1 U1056 ( .A1(n957), .A2(n956), .ZN(n967) );
  XNOR2_X1 U1057 ( .A(G171), .B(G1961), .ZN(n958) );
  XNOR2_X1 U1058 ( .A(n958), .B(KEYINPUT120), .ZN(n962) );
  NOR2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n965) );
  XNOR2_X1 U1061 ( .A(KEYINPUT121), .B(n963), .ZN(n964) );
  NOR2_X1 U1062 ( .A1(n965), .A2(n964), .ZN(n966) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NOR2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n970) );
  XNOR2_X1 U1065 ( .A(KEYINPUT122), .B(n970), .ZN(n971) );
  NAND2_X1 U1066 ( .A1(n972), .A2(n971), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(n975), .B(KEYINPUT123), .ZN(n1002) );
  XOR2_X1 U1069 ( .A(G2067), .B(G26), .Z(n976) );
  NAND2_X1 U1070 ( .A1(n976), .A2(G28), .ZN(n983) );
  XNOR2_X1 U1071 ( .A(G27), .B(n977), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(G1991), .B(G25), .ZN(n979) );
  XNOR2_X1 U1073 ( .A(G33), .B(G2072), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1075 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1076 ( .A1(n983), .A2(n982), .ZN(n987) );
  XOR2_X1 U1077 ( .A(n984), .B(G32), .Z(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT117), .B(n985), .ZN(n986) );
  NAND2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1080 ( .A(KEYINPUT53), .B(n988), .ZN(n992) );
  XOR2_X1 U1081 ( .A(G34), .B(KEYINPUT118), .Z(n990) );
  XNOR2_X1 U1082 ( .A(G2084), .B(KEYINPUT54), .ZN(n989) );
  XNOR2_X1 U1083 ( .A(n990), .B(n989), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n995) );
  XNOR2_X1 U1085 ( .A(KEYINPUT116), .B(G2090), .ZN(n993) );
  XNOR2_X1 U1086 ( .A(G35), .B(n993), .ZN(n994) );
  NOR2_X1 U1087 ( .A1(n995), .A2(n994), .ZN(n996) );
  XNOR2_X1 U1088 ( .A(n996), .B(KEYINPUT55), .ZN(n998) );
  INV_X1 U1089 ( .A(G29), .ZN(n997) );
  NAND2_X1 U1090 ( .A1(n998), .A2(n997), .ZN(n999) );
  NAND2_X1 U1091 ( .A1(G11), .A2(n999), .ZN(n1000) );
  XOR2_X1 U1092 ( .A(KEYINPUT119), .B(n1000), .Z(n1001) );
  NOR2_X1 U1093 ( .A1(n1002), .A2(n1001), .ZN(n1032) );
  XOR2_X1 U1094 ( .A(G2090), .B(G162), .Z(n1003) );
  NOR2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  XOR2_X1 U1096 ( .A(KEYINPUT51), .B(n1005), .Z(n1006) );
  XNOR2_X1 U1097 ( .A(KEYINPUT114), .B(n1006), .ZN(n1024) );
  INV_X1 U1098 ( .A(n1007), .ZN(n1011) );
  NOR2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1100 ( .A1(n1011), .A2(n1010), .ZN(n1013) );
  XOR2_X1 U1101 ( .A(G160), .B(G2084), .Z(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  NAND2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1022) );
  XNOR2_X1 U1104 ( .A(G2072), .B(n1016), .ZN(n1018) );
  XNOR2_X1 U1105 ( .A(G164), .B(G2078), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XOR2_X1 U1107 ( .A(KEYINPUT115), .B(n1019), .Z(n1020) );
  XNOR2_X1 U1108 ( .A(KEYINPUT50), .B(n1020), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NOR2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(KEYINPUT52), .B(n1027), .ZN(n1029) );
  INV_X1 U1113 ( .A(KEYINPUT55), .ZN(n1028) );
  NAND2_X1 U1114 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(G29), .ZN(n1031) );
  NAND2_X1 U1116 ( .A1(n1032), .A2(n1031), .ZN(n1033) );
  NOR2_X1 U1117 ( .A1(n1034), .A2(n1033), .ZN(n1035) );
  XOR2_X1 U1118 ( .A(KEYINPUT62), .B(n1035), .Z(n1036) );
  XNOR2_X1 U1119 ( .A(KEYINPUT127), .B(n1036), .ZN(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

