

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809;

  AND2_X1 U380 ( .A1(n396), .A2(n366), .ZN(n358) );
  BUF_X1 U381 ( .A(n717), .Z(n427) );
  BUF_X1 U382 ( .A(n581), .Z(n595) );
  OR2_X1 U383 ( .A1(n758), .A2(n439), .ZN(n438) );
  XNOR2_X1 U384 ( .A(n486), .B(n485), .ZN(n540) );
  XNOR2_X1 U385 ( .A(n425), .B(G119), .ZN(n424) );
  INV_X2 U386 ( .A(G143), .ZN(n474) );
  NAND2_X1 U387 ( .A1(n358), .A2(n454), .ZN(n674) );
  XNOR2_X2 U388 ( .A(n565), .B(n564), .ZN(n631) );
  INV_X2 U389 ( .A(KEYINPUT3), .ZN(n425) );
  XNOR2_X2 U390 ( .A(n540), .B(n365), .ZN(n794) );
  XNOR2_X1 U391 ( .A(n359), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U392 ( .A1(n766), .A2(n777), .ZN(n359) );
  XNOR2_X1 U393 ( .A(G113), .B(G143), .ZN(n549) );
  XNOR2_X1 U394 ( .A(G113), .B(G116), .ZN(n423) );
  INV_X1 U395 ( .A(G953), .ZN(n797) );
  XOR2_X1 U396 ( .A(KEYINPUT24), .B(KEYINPUT92), .Z(n360) );
  AND2_X2 U397 ( .A1(n443), .A2(n442), .ZN(n441) );
  OR2_X2 U398 ( .A1(n696), .A2(n736), .ZN(n640) );
  XNOR2_X2 U399 ( .A(n786), .B(n487), .ZN(n522) );
  INV_X1 U400 ( .A(n723), .ZN(n622) );
  INV_X1 U401 ( .A(n796), .ZN(n361) );
  NAND2_X1 U402 ( .A1(n402), .A2(n405), .ZN(n404) );
  NAND2_X1 U403 ( .A1(n664), .A2(n663), .ZN(n796) );
  NAND2_X1 U404 ( .A1(n588), .A2(n620), .ZN(n692) );
  INV_X1 U405 ( .A(n595), .ZN(n384) );
  INV_X1 U406 ( .A(n620), .ZN(n719) );
  XNOR2_X1 U407 ( .A(n431), .B(n541), .ZN(n599) );
  NOR2_X1 U408 ( .A1(n769), .A2(G902), .ZN(n431) );
  XNOR2_X1 U409 ( .A(n524), .B(n490), .ZN(n758) );
  XNOR2_X1 U410 ( .A(n763), .B(n762), .ZN(n764) );
  XNOR2_X1 U411 ( .A(n449), .B(G125), .ZN(n492) );
  XNOR2_X2 U412 ( .A(n641), .B(n640), .ZN(n809) );
  NAND2_X1 U413 ( .A1(n397), .A2(n584), .ZN(n586) );
  NOR2_X2 U414 ( .A1(n754), .A2(n777), .ZN(n756) );
  XNOR2_X2 U415 ( .A(n794), .B(G146), .ZN(n524) );
  NOR2_X1 U416 ( .A1(n665), .A2(KEYINPUT81), .ZN(n405) );
  NOR2_X1 U417 ( .A1(n648), .A2(n649), .ZN(n656) );
  NAND2_X1 U418 ( .A1(n362), .A2(n441), .ZN(n437) );
  NAND2_X1 U419 ( .A1(n393), .A2(n389), .ZN(n388) );
  AND2_X1 U420 ( .A1(n390), .A2(n626), .ZN(n389) );
  NAND2_X1 U421 ( .A1(n668), .A2(KEYINPUT66), .ZN(n457) );
  AND2_X1 U422 ( .A1(n373), .A2(n406), .ZN(n403) );
  NOR2_X1 U423 ( .A1(n654), .A2(n655), .ZN(n401) );
  INV_X1 U424 ( .A(G146), .ZN(n449) );
  XNOR2_X1 U425 ( .A(n460), .B(KEYINPUT70), .ZN(n487) );
  INV_X1 U426 ( .A(G101), .ZN(n460) );
  XNOR2_X1 U427 ( .A(n461), .B(G140), .ZN(n494) );
  INV_X1 U428 ( .A(G137), .ZN(n461) );
  INV_X1 U429 ( .A(KEYINPUT39), .ZN(n421) );
  NAND2_X1 U430 ( .A1(n491), .A2(n440), .ZN(n439) );
  NAND2_X1 U431 ( .A1(G469), .A2(G902), .ZN(n442) );
  XNOR2_X1 U432 ( .A(n472), .B(n471), .ZN(n489) );
  INV_X1 U433 ( .A(G104), .ZN(n471) );
  XNOR2_X1 U434 ( .A(G110), .B(G107), .ZN(n472) );
  XNOR2_X1 U435 ( .A(n494), .B(n487), .ZN(n459) );
  XNOR2_X1 U436 ( .A(n639), .B(n432), .ZN(n736) );
  XNOR2_X1 U437 ( .A(n433), .B(KEYINPUT41), .ZN(n432) );
  INV_X1 U438 ( .A(KEYINPUT112), .ZN(n433) );
  NAND2_X1 U439 ( .A1(n708), .A2(n421), .ZN(n419) );
  INV_X1 U440 ( .A(n419), .ZN(n415) );
  NAND2_X1 U441 ( .A1(n412), .A2(n418), .ZN(n416) );
  NOR2_X1 U442 ( .A1(n708), .A2(n421), .ZN(n418) );
  INV_X1 U443 ( .A(n638), .ZN(n412) );
  NAND2_X1 U444 ( .A1(n656), .A2(n650), .ZN(n446) );
  AND2_X1 U445 ( .A1(n427), .A2(n622), .ZN(n450) );
  XNOR2_X1 U446 ( .A(n508), .B(n507), .ZN(n620) );
  XNOR2_X1 U447 ( .A(n506), .B(n470), .ZN(n507) );
  INV_X1 U448 ( .A(KEYINPUT6), .ZN(n447) );
  AND2_X1 U449 ( .A1(n680), .A2(G953), .ZN(n777) );
  NAND2_X1 U450 ( .A1(n392), .A2(n391), .ZN(n390) );
  INV_X1 U451 ( .A(KEYINPUT96), .ZN(n391) );
  XNOR2_X1 U452 ( .A(G902), .B(KEYINPUT15), .ZN(n665) );
  INV_X1 U453 ( .A(G237), .ZN(n484) );
  XNOR2_X1 U454 ( .A(n375), .B(KEYINPUT73), .ZN(n592) );
  NOR2_X1 U455 ( .A1(n717), .A2(n716), .ZN(n375) );
  XOR2_X1 U456 ( .A(G137), .B(KEYINPUT5), .Z(n520) );
  NOR2_X1 U457 ( .A1(G953), .A2(G237), .ZN(n542) );
  XOR2_X1 U458 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n479) );
  XNOR2_X1 U459 ( .A(KEYINPUT4), .B(KEYINPUT87), .ZN(n478) );
  XNOR2_X1 U460 ( .A(n492), .B(n448), .ZN(n477) );
  INV_X1 U461 ( .A(KEYINPUT89), .ZN(n448) );
  NAND2_X1 U462 ( .A1(G234), .A2(G237), .ZN(n512) );
  NOR2_X1 U463 ( .A1(n706), .A2(n708), .ZN(n714) );
  NAND2_X1 U464 ( .A1(n719), .A2(n720), .ZN(n716) );
  XNOR2_X1 U465 ( .A(KEYINPUT16), .B(G122), .ZN(n473) );
  XNOR2_X1 U466 ( .A(n498), .B(n360), .ZN(n428) );
  XOR2_X1 U467 ( .A(KEYINPUT94), .B(KEYINPUT93), .Z(n498) );
  INV_X1 U468 ( .A(G134), .ZN(n485) );
  XOR2_X1 U469 ( .A(KEYINPUT97), .B(KEYINPUT12), .Z(n544) );
  INV_X1 U470 ( .A(KEYINPUT10), .ZN(n493) );
  XOR2_X1 U471 ( .A(G122), .B(G104), .Z(n550) );
  XNOR2_X1 U472 ( .A(G131), .B(G140), .ZN(n545) );
  XOR2_X1 U473 ( .A(KEYINPUT98), .B(KEYINPUT11), .Z(n546) );
  NOR2_X1 U474 ( .A1(n671), .A2(n672), .ZN(n741) );
  XNOR2_X1 U475 ( .A(n582), .B(n371), .ZN(n397) );
  XNOR2_X1 U476 ( .A(n400), .B(KEYINPUT106), .ZN(n560) );
  OR2_X1 U477 ( .A1(n427), .A2(n719), .ZN(n400) );
  BUF_X1 U478 ( .A(n381), .Z(n773) );
  XNOR2_X1 U479 ( .A(n459), .B(n369), .ZN(n488) );
  XOR2_X1 U480 ( .A(n751), .B(n750), .Z(n752) );
  NAND2_X1 U481 ( .A1(n417), .A2(n416), .ZN(n661) );
  XNOR2_X1 U482 ( .A(n422), .B(KEYINPUT40), .ZN(n808) );
  NAND2_X1 U483 ( .A1(n413), .A2(n416), .ZN(n422) );
  NOR2_X1 U484 ( .A1(n415), .A2(n700), .ZN(n414) );
  AND2_X1 U485 ( .A1(n445), .A2(n444), .ZN(n652) );
  INV_X1 U486 ( .A(n427), .ZN(n444) );
  XNOR2_X1 U487 ( .A(n446), .B(n651), .ZN(n445) );
  AND2_X1 U488 ( .A1(n466), .A2(n467), .ZN(n465) );
  XNOR2_X1 U489 ( .A(n451), .B(n587), .ZN(n588) );
  NAND2_X1 U490 ( .A1(n382), .A2(n450), .ZN(n451) );
  INV_X1 U491 ( .A(KEYINPUT84), .ZN(n429) );
  INV_X1 U492 ( .A(KEYINPUT63), .ZN(n453) );
  AND2_X1 U493 ( .A1(n438), .A2(KEYINPUT1), .ZN(n362) );
  AND2_X1 U494 ( .A1(n526), .A2(G210), .ZN(n363) );
  XOR2_X1 U495 ( .A(n675), .B(KEYINPUT71), .Z(n364) );
  XOR2_X1 U496 ( .A(KEYINPUT4), .B(G131), .Z(n365) );
  AND2_X1 U497 ( .A1(n395), .A2(n457), .ZN(n366) );
  AND2_X1 U498 ( .A1(n374), .A2(n406), .ZN(n367) );
  AND2_X1 U499 ( .A1(n407), .A2(n403), .ZN(n368) );
  AND2_X1 U500 ( .A1(G227), .A2(n797), .ZN(n369) );
  AND2_X1 U501 ( .A1(n689), .A2(KEYINPUT96), .ZN(n370) );
  INV_X1 U502 ( .A(G902), .ZN(n440) );
  XOR2_X1 U503 ( .A(KEYINPUT34), .B(KEYINPUT75), .Z(n371) );
  XOR2_X1 U504 ( .A(n518), .B(KEYINPUT30), .Z(n372) );
  INV_X1 U505 ( .A(KEYINPUT31), .ZN(n468) );
  AND2_X1 U506 ( .A1(n669), .A2(n458), .ZN(n373) );
  NAND2_X1 U507 ( .A1(n670), .A2(KEYINPUT81), .ZN(n374) );
  NAND2_X1 U508 ( .A1(n670), .A2(KEYINPUT81), .ZN(n407) );
  XNOR2_X2 U509 ( .A(n575), .B(n574), .ZN(n382) );
  INV_X1 U510 ( .A(n689), .ZN(n392) );
  NAND2_X1 U511 ( .A1(n387), .A2(n385), .ZN(n602) );
  NAND2_X1 U512 ( .A1(n601), .A2(n719), .ZN(n683) );
  NOR2_X1 U513 ( .A1(n604), .A2(n603), .ZN(n605) );
  NAND2_X1 U514 ( .A1(n602), .A2(n683), .ZN(n603) );
  NAND2_X1 U515 ( .A1(n796), .A2(n373), .ZN(n395) );
  XNOR2_X1 U516 ( .A(n430), .B(n429), .ZN(n601) );
  BUF_X1 U517 ( .A(n735), .Z(n398) );
  NAND2_X1 U518 ( .A1(n386), .A2(n391), .ZN(n385) );
  INV_X1 U519 ( .A(n702), .ZN(n386) );
  NAND2_X1 U520 ( .A1(n702), .A2(n370), .ZN(n393) );
  NAND2_X1 U521 ( .A1(n692), .A2(n378), .ZN(n376) );
  NAND2_X1 U522 ( .A1(n376), .A2(n377), .ZN(n604) );
  OR2_X1 U523 ( .A1(n589), .A2(KEYINPUT44), .ZN(n377) );
  AND2_X1 U524 ( .A1(n608), .A2(KEYINPUT67), .ZN(n378) );
  NAND2_X1 U525 ( .A1(n692), .A2(n608), .ZN(n379) );
  XNOR2_X1 U526 ( .A(n586), .B(n585), .ZN(n380) );
  XNOR2_X1 U527 ( .A(n586), .B(n585), .ZN(n434) );
  AND2_X2 U528 ( .A1(n674), .A2(n673), .ZN(n381) );
  BUF_X1 U529 ( .A(n631), .Z(n383) );
  AND2_X1 U530 ( .A1(n595), .A2(KEYINPUT31), .ZN(n464) );
  NAND2_X1 U531 ( .A1(n384), .A2(n468), .ZN(n466) );
  NOR2_X2 U532 ( .A1(n735), .A2(n384), .ZN(n582) );
  INV_X1 U533 ( .A(n388), .ZN(n387) );
  NAND2_X2 U534 ( .A1(n465), .A2(n462), .ZN(n702) );
  NOR2_X1 U535 ( .A1(n394), .A2(n675), .ZN(n679) );
  NAND2_X1 U536 ( .A1(n674), .A2(n673), .ZN(n394) );
  NAND2_X1 U537 ( .A1(n368), .A2(n404), .ZN(n396) );
  NAND2_X1 U538 ( .A1(n381), .A2(G475), .ZN(n765) );
  XNOR2_X2 U539 ( .A(n409), .B(n613), .ZN(n670) );
  NAND2_X1 U540 ( .A1(n379), .A2(n589), .ZN(n590) );
  XNOR2_X1 U541 ( .A(n399), .B(KEYINPUT85), .ZN(n410) );
  NAND2_X1 U542 ( .A1(n605), .A2(n606), .ZN(n399) );
  NAND2_X1 U543 ( .A1(n436), .A2(n558), .ZN(n435) );
  NAND2_X1 U544 ( .A1(n749), .A2(n665), .ZN(n426) );
  XNOR2_X1 U545 ( .A(n483), .B(n482), .ZN(n749) );
  XNOR2_X1 U546 ( .A(n571), .B(n469), .ZN(n581) );
  XNOR2_X1 U547 ( .A(n401), .B(KEYINPUT48), .ZN(n664) );
  NOR2_X1 U548 ( .A1(n645), .A2(n646), .ZN(n647) );
  NAND2_X1 U549 ( .A1(n437), .A2(n435), .ZN(n717) );
  INV_X1 U550 ( .A(n670), .ZN(n402) );
  NAND2_X1 U551 ( .A1(n367), .A2(n404), .ZN(n408) );
  NAND2_X1 U552 ( .A1(n665), .A2(KEYINPUT81), .ZN(n406) );
  NAND2_X1 U553 ( .A1(n408), .A2(n455), .ZN(n454) );
  NAND2_X1 U554 ( .A1(n410), .A2(n612), .ZN(n409) );
  XNOR2_X1 U555 ( .A(n411), .B(n372), .ZN(n527) );
  NAND2_X1 U556 ( .A1(n723), .A2(n711), .ZN(n411) );
  XNOR2_X2 U557 ( .A(n525), .B(n364), .ZN(n723) );
  AND2_X1 U558 ( .A1(n420), .A2(n419), .ZN(n417) );
  AND2_X1 U559 ( .A1(n420), .A2(n414), .ZN(n413) );
  NAND2_X1 U560 ( .A1(n638), .A2(n421), .ZN(n420) );
  XNOR2_X2 U561 ( .A(n424), .B(n423), .ZN(n786) );
  INV_X1 U562 ( .A(n563), .ZN(n561) );
  XNOR2_X2 U563 ( .A(n426), .B(n363), .ZN(n563) );
  XNOR2_X2 U564 ( .A(n580), .B(KEYINPUT33), .ZN(n735) );
  XNOR2_X2 U565 ( .A(n578), .B(n577), .ZN(n608) );
  NAND2_X1 U566 ( .A1(n600), .A2(n645), .ZN(n430) );
  NOR2_X2 U567 ( .A1(n592), .A2(n645), .ZN(n580) );
  XNOR2_X1 U568 ( .A(n428), .B(n499), .ZN(n502) );
  NAND2_X1 U569 ( .A1(n434), .A2(n590), .ZN(n591) );
  NAND2_X1 U570 ( .A1(n380), .A2(n607), .ZN(n610) );
  XNOR2_X1 U571 ( .A(n380), .B(G122), .ZN(G24) );
  NAND2_X1 U572 ( .A1(n441), .A2(n438), .ZN(n436) );
  NAND2_X1 U573 ( .A1(n441), .A2(n438), .ZN(n452) );
  NAND2_X1 U574 ( .A1(n758), .A2(G469), .ZN(n443) );
  XNOR2_X2 U575 ( .A(n622), .B(n447), .ZN(n645) );
  AND2_X1 U576 ( .A1(n382), .A2(n427), .ZN(n600) );
  XNOR2_X1 U577 ( .A(n682), .B(n453), .ZN(G57) );
  NAND2_X1 U578 ( .A1(n511), .A2(n452), .ZN(n593) );
  NAND2_X1 U579 ( .A1(n625), .A2(n452), .ZN(n696) );
  AND2_X1 U580 ( .A1(n361), .A2(KEYINPUT66), .ZN(n455) );
  INV_X1 U581 ( .A(KEYINPUT66), .ZN(n458) );
  NAND2_X1 U582 ( .A1(n464), .A2(n463), .ZN(n462) );
  INV_X1 U583 ( .A(n726), .ZN(n463) );
  NAND2_X1 U584 ( .A1(n726), .A2(n468), .ZN(n467) );
  XNOR2_X1 U585 ( .A(n492), .B(n493), .ZN(n552) );
  XOR2_X1 U586 ( .A(n570), .B(KEYINPUT0), .Z(n469) );
  XOR2_X1 U587 ( .A(KEYINPUT25), .B(KEYINPUT74), .Z(n470) );
  INV_X1 U588 ( .A(G469), .ZN(n491) );
  INV_X1 U589 ( .A(n494), .ZN(n495) );
  XNOR2_X1 U590 ( .A(n489), .B(n488), .ZN(n490) );
  XNOR2_X1 U591 ( .A(n552), .B(n495), .ZN(n793) );
  INV_X1 U592 ( .A(KEYINPUT68), .ZN(n587) );
  XNOR2_X1 U593 ( .A(n769), .B(n768), .ZN(n770) );
  XNOR2_X1 U594 ( .A(n771), .B(n770), .ZN(n772) );
  XNOR2_X1 U595 ( .A(n489), .B(n473), .ZN(n785) );
  XNOR2_X1 U596 ( .A(n522), .B(n785), .ZN(n483) );
  XNOR2_X2 U597 ( .A(n474), .B(G128), .ZN(n486) );
  NAND2_X1 U598 ( .A1(G224), .A2(n797), .ZN(n475) );
  XNOR2_X1 U599 ( .A(n486), .B(n475), .ZN(n476) );
  XNOR2_X1 U600 ( .A(n476), .B(n477), .ZN(n481) );
  XNOR2_X1 U601 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U602 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U603 ( .A1(n440), .A2(n484), .ZN(n526) );
  INV_X1 U604 ( .A(n561), .ZN(n650) );
  XOR2_X1 U605 ( .A(KEYINPUT23), .B(G110), .Z(n497) );
  XNOR2_X1 U606 ( .A(G119), .B(G128), .ZN(n496) );
  XNOR2_X1 U607 ( .A(n497), .B(n496), .ZN(n499) );
  NAND2_X1 U608 ( .A1(G234), .A2(n797), .ZN(n500) );
  XOR2_X1 U609 ( .A(KEYINPUT8), .B(n500), .Z(n536) );
  NAND2_X1 U610 ( .A1(G221), .A2(n536), .ZN(n501) );
  XNOR2_X1 U611 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U612 ( .A(n503), .B(n793), .ZN(n774) );
  NOR2_X1 U613 ( .A1(n774), .A2(G902), .ZN(n508) );
  XOR2_X1 U614 ( .A(KEYINPUT95), .B(KEYINPUT20), .Z(n505) );
  NAND2_X1 U615 ( .A1(G234), .A2(n665), .ZN(n504) );
  XNOR2_X1 U616 ( .A(n505), .B(n504), .ZN(n509) );
  NAND2_X1 U617 ( .A1(G217), .A2(n509), .ZN(n506) );
  AND2_X1 U618 ( .A1(n509), .A2(G221), .ZN(n510) );
  XNOR2_X1 U619 ( .A(n510), .B(KEYINPUT21), .ZN(n720) );
  INV_X1 U620 ( .A(n716), .ZN(n511) );
  INV_X1 U621 ( .A(n593), .ZN(n529) );
  XNOR2_X1 U622 ( .A(n512), .B(KEYINPUT14), .ZN(n514) );
  NAND2_X1 U623 ( .A1(G952), .A2(n514), .ZN(n734) );
  NOR2_X1 U624 ( .A1(n734), .A2(G953), .ZN(n513) );
  XNOR2_X1 U625 ( .A(n513), .B(KEYINPUT90), .ZN(n567) );
  NAND2_X1 U626 ( .A1(n514), .A2(G902), .ZN(n515) );
  XNOR2_X1 U627 ( .A(n515), .B(KEYINPUT91), .ZN(n566) );
  NAND2_X1 U628 ( .A1(n566), .A2(G953), .ZN(n516) );
  NOR2_X1 U629 ( .A1(G900), .A2(n516), .ZN(n517) );
  NOR2_X1 U630 ( .A1(n567), .A2(n517), .ZN(n619) );
  XNOR2_X1 U631 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n518) );
  NAND2_X1 U632 ( .A1(n542), .A2(G210), .ZN(n519) );
  XNOR2_X1 U633 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U634 ( .A(n522), .B(n521), .ZN(n523) );
  XNOR2_X1 U635 ( .A(n524), .B(n523), .ZN(n677) );
  NOR2_X1 U636 ( .A1(n677), .A2(G902), .ZN(n525) );
  INV_X1 U637 ( .A(G472), .ZN(n675) );
  NAND2_X1 U638 ( .A1(n526), .A2(G214), .ZN(n711) );
  NOR2_X1 U639 ( .A1(n619), .A2(n527), .ZN(n528) );
  NAND2_X1 U640 ( .A1(n529), .A2(n528), .ZN(n638) );
  XOR2_X1 U641 ( .A(KEYINPUT101), .B(G122), .Z(n531) );
  XNOR2_X1 U642 ( .A(G116), .B(G107), .ZN(n530) );
  XNOR2_X1 U643 ( .A(n531), .B(n530), .ZN(n535) );
  XOR2_X1 U644 ( .A(KEYINPUT7), .B(KEYINPUT100), .Z(n533) );
  XNOR2_X1 U645 ( .A(KEYINPUT9), .B(KEYINPUT102), .ZN(n532) );
  XNOR2_X1 U646 ( .A(n533), .B(n532), .ZN(n534) );
  XOR2_X1 U647 ( .A(n535), .B(n534), .Z(n538) );
  NAND2_X1 U648 ( .A1(G217), .A2(n536), .ZN(n537) );
  XNOR2_X1 U649 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U650 ( .A(n540), .B(n539), .ZN(n769) );
  XNOR2_X1 U651 ( .A(KEYINPUT103), .B(G478), .ZN(n541) );
  XNOR2_X1 U652 ( .A(KEYINPUT13), .B(G475), .ZN(n556) );
  NAND2_X1 U653 ( .A1(G214), .A2(n542), .ZN(n543) );
  XNOR2_X1 U654 ( .A(n544), .B(n543), .ZN(n548) );
  XNOR2_X1 U655 ( .A(n546), .B(n545), .ZN(n547) );
  XOR2_X1 U656 ( .A(n548), .B(n547), .Z(n554) );
  XNOR2_X1 U657 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U658 ( .A(n552), .B(n551), .ZN(n553) );
  XNOR2_X1 U659 ( .A(n554), .B(n553), .ZN(n763) );
  NOR2_X1 U660 ( .A1(G902), .A2(n763), .ZN(n555) );
  XNOR2_X1 U661 ( .A(n556), .B(n555), .ZN(n596) );
  NAND2_X1 U662 ( .A1(n599), .A2(n596), .ZN(n583) );
  NOR2_X1 U663 ( .A1(n638), .A2(n583), .ZN(n557) );
  NAND2_X1 U664 ( .A1(n650), .A2(n557), .ZN(n615) );
  XNOR2_X1 U665 ( .A(n615), .B(G143), .ZN(G45) );
  INV_X1 U666 ( .A(KEYINPUT1), .ZN(n558) );
  INV_X1 U667 ( .A(n645), .ZN(n559) );
  NOR2_X1 U668 ( .A1(n560), .A2(n559), .ZN(n576) );
  INV_X1 U669 ( .A(n711), .ZN(n562) );
  NAND2_X1 U670 ( .A1(n563), .A2(n711), .ZN(n565) );
  INV_X1 U671 ( .A(KEYINPUT19), .ZN(n564) );
  NOR2_X1 U672 ( .A1(G898), .A2(n797), .ZN(n789) );
  AND2_X1 U673 ( .A1(n566), .A2(n789), .ZN(n568) );
  NOR2_X1 U674 ( .A1(n568), .A2(n567), .ZN(n569) );
  NOR2_X2 U675 ( .A1(n631), .A2(n569), .ZN(n571) );
  INV_X1 U676 ( .A(KEYINPUT86), .ZN(n570) );
  NOR2_X1 U677 ( .A1(n599), .A2(n596), .ZN(n572) );
  XNOR2_X1 U678 ( .A(n572), .B(KEYINPUT105), .ZN(n706) );
  INV_X1 U679 ( .A(n720), .ZN(n618) );
  NOR2_X1 U680 ( .A1(n706), .A2(n618), .ZN(n573) );
  NAND2_X1 U681 ( .A1(n581), .A2(n573), .ZN(n575) );
  INV_X1 U682 ( .A(KEYINPUT22), .ZN(n574) );
  NAND2_X1 U683 ( .A1(n382), .A2(n576), .ZN(n578) );
  XNOR2_X1 U684 ( .A(KEYINPUT76), .B(KEYINPUT32), .ZN(n577) );
  XOR2_X1 U685 ( .A(G119), .B(KEYINPUT127), .Z(n579) );
  XNOR2_X1 U686 ( .A(n608), .B(n579), .ZN(G21) );
  INV_X1 U687 ( .A(n583), .ZN(n584) );
  XNOR2_X1 U688 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n585) );
  INV_X1 U689 ( .A(KEYINPUT67), .ZN(n589) );
  NAND2_X1 U690 ( .A1(n591), .A2(KEYINPUT44), .ZN(n606) );
  OR2_X1 U691 ( .A1(n592), .A2(n622), .ZN(n726) );
  NOR2_X1 U692 ( .A1(n723), .A2(n593), .ZN(n594) );
  NAND2_X1 U693 ( .A1(n595), .A2(n594), .ZN(n689) );
  XNOR2_X1 U694 ( .A(n596), .B(KEYINPUT99), .ZN(n598) );
  NAND2_X1 U695 ( .A1(n598), .A2(n599), .ZN(n597) );
  XNOR2_X1 U696 ( .A(n597), .B(KEYINPUT104), .ZN(n703) );
  NOR2_X1 U697 ( .A1(n599), .A2(n598), .ZN(n644) );
  INV_X1 U698 ( .A(n644), .ZN(n700) );
  NAND2_X1 U699 ( .A1(n703), .A2(n700), .ZN(n626) );
  INV_X1 U700 ( .A(KEYINPUT44), .ZN(n607) );
  INV_X1 U701 ( .A(n608), .ZN(n609) );
  NOR2_X1 U702 ( .A1(n610), .A2(n609), .ZN(n611) );
  NAND2_X1 U703 ( .A1(n611), .A2(n692), .ZN(n612) );
  XNOR2_X1 U704 ( .A(KEYINPUT65), .B(KEYINPUT45), .ZN(n613) );
  INV_X1 U705 ( .A(n626), .ZN(n707) );
  NAND2_X1 U706 ( .A1(KEYINPUT47), .A2(n707), .ZN(n614) );
  XNOR2_X1 U707 ( .A(n614), .B(KEYINPUT78), .ZN(n616) );
  NAND2_X1 U708 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U709 ( .A(KEYINPUT77), .B(n617), .ZN(n636) );
  NOR2_X1 U710 ( .A1(n619), .A2(n618), .ZN(n621) );
  NAND2_X1 U711 ( .A1(n621), .A2(n620), .ZN(n646) );
  OR2_X1 U712 ( .A1(n622), .A2(n646), .ZN(n624) );
  XNOR2_X1 U713 ( .A(KEYINPUT28), .B(KEYINPUT111), .ZN(n623) );
  XNOR2_X1 U714 ( .A(n624), .B(n623), .ZN(n625) );
  INV_X1 U715 ( .A(n696), .ZN(n629) );
  INV_X1 U716 ( .A(KEYINPUT47), .ZN(n632) );
  NAND2_X1 U717 ( .A1(n632), .A2(n626), .ZN(n627) );
  XNOR2_X1 U718 ( .A(n627), .B(KEYINPUT72), .ZN(n628) );
  AND2_X1 U719 ( .A1(n629), .A2(n628), .ZN(n630) );
  INV_X1 U720 ( .A(n383), .ZN(n697) );
  NAND2_X1 U721 ( .A1(n630), .A2(n697), .ZN(n634) );
  OR2_X1 U722 ( .A1(n696), .A2(n383), .ZN(n693) );
  NAND2_X1 U723 ( .A1(n693), .A2(n632), .ZN(n633) );
  NAND2_X1 U724 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U725 ( .A1(n636), .A2(n635), .ZN(n655) );
  XOR2_X1 U726 ( .A(KEYINPUT64), .B(KEYINPUT46), .Z(n643) );
  INV_X1 U727 ( .A(KEYINPUT38), .ZN(n637) );
  XNOR2_X1 U728 ( .A(n561), .B(n637), .ZN(n708) );
  XOR2_X1 U729 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n641) );
  NAND2_X1 U730 ( .A1(n711), .A2(n714), .ZN(n639) );
  NAND2_X1 U731 ( .A1(n808), .A2(n809), .ZN(n642) );
  XNOR2_X1 U732 ( .A(n643), .B(n642), .ZN(n653) );
  XOR2_X1 U733 ( .A(KEYINPUT36), .B(KEYINPUT114), .Z(n651) );
  NAND2_X1 U734 ( .A1(n644), .A2(n711), .ZN(n649) );
  XNOR2_X1 U735 ( .A(n647), .B(KEYINPUT107), .ZN(n648) );
  XNOR2_X1 U736 ( .A(KEYINPUT115), .B(n652), .ZN(n806) );
  NAND2_X1 U737 ( .A1(n653), .A2(n806), .ZN(n654) );
  NAND2_X1 U738 ( .A1(n427), .A2(n656), .ZN(n657) );
  XNOR2_X1 U739 ( .A(n657), .B(KEYINPUT43), .ZN(n658) );
  AND2_X1 U740 ( .A1(n561), .A2(n658), .ZN(n660) );
  INV_X1 U741 ( .A(KEYINPUT108), .ZN(n659) );
  XNOR2_X1 U742 ( .A(n660), .B(n659), .ZN(n807) );
  NOR2_X1 U743 ( .A1(n703), .A2(n661), .ZN(n705) );
  INV_X1 U744 ( .A(n705), .ZN(n662) );
  AND2_X1 U745 ( .A1(n807), .A2(n662), .ZN(n663) );
  XOR2_X1 U746 ( .A(n665), .B(KEYINPUT82), .Z(n666) );
  NAND2_X1 U747 ( .A1(n666), .A2(KEYINPUT2), .ZN(n667) );
  XNOR2_X1 U748 ( .A(n667), .B(KEYINPUT69), .ZN(n668) );
  INV_X1 U749 ( .A(n668), .ZN(n669) );
  BUF_X1 U750 ( .A(n670), .Z(n671) );
  NAND2_X1 U751 ( .A1(n361), .A2(KEYINPUT2), .ZN(n672) );
  INV_X1 U752 ( .A(n741), .ZN(n673) );
  XOR2_X1 U753 ( .A(KEYINPUT88), .B(KEYINPUT62), .Z(n676) );
  XNOR2_X1 U754 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U755 ( .A(n679), .B(n678), .ZN(n681) );
  INV_X1 U756 ( .A(G952), .ZN(n680) );
  NOR2_X1 U757 ( .A1(n681), .A2(n777), .ZN(n682) );
  XNOR2_X1 U758 ( .A(G101), .B(KEYINPUT116), .ZN(n684) );
  XNOR2_X1 U759 ( .A(n684), .B(n683), .ZN(G3) );
  NOR2_X1 U760 ( .A1(n700), .A2(n689), .ZN(n686) );
  XNOR2_X1 U761 ( .A(G104), .B(KEYINPUT117), .ZN(n685) );
  XNOR2_X1 U762 ( .A(n686), .B(n685), .ZN(G6) );
  XOR2_X1 U763 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n688) );
  XNOR2_X1 U764 ( .A(G107), .B(KEYINPUT118), .ZN(n687) );
  XNOR2_X1 U765 ( .A(n688), .B(n687), .ZN(n691) );
  NOR2_X1 U766 ( .A1(n703), .A2(n689), .ZN(n690) );
  XOR2_X1 U767 ( .A(n691), .B(n690), .Z(G9) );
  XNOR2_X1 U768 ( .A(G110), .B(n692), .ZN(G12) );
  NOR2_X1 U769 ( .A1(n693), .A2(n703), .ZN(n695) );
  XNOR2_X1 U770 ( .A(G128), .B(KEYINPUT29), .ZN(n694) );
  XNOR2_X1 U771 ( .A(n695), .B(n694), .ZN(G30) );
  NOR2_X1 U772 ( .A1(n696), .A2(n700), .ZN(n698) );
  NAND2_X1 U773 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U774 ( .A(n699), .B(G146), .ZN(G48) );
  NOR2_X1 U775 ( .A1(n700), .A2(n702), .ZN(n701) );
  XOR2_X1 U776 ( .A(G113), .B(n701), .Z(G15) );
  NOR2_X1 U777 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U778 ( .A(G116), .B(n704), .Z(G18) );
  XOR2_X1 U779 ( .A(G134), .B(n705), .Z(G36) );
  INV_X1 U780 ( .A(n706), .ZN(n710) );
  NOR2_X1 U781 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U782 ( .A1(n710), .A2(n709), .ZN(n712) );
  NOR2_X1 U783 ( .A1(n712), .A2(n562), .ZN(n713) );
  NOR2_X1 U784 ( .A1(n714), .A2(n713), .ZN(n715) );
  NOR2_X1 U785 ( .A1(n398), .A2(n715), .ZN(n731) );
  NAND2_X1 U786 ( .A1(n427), .A2(n716), .ZN(n718) );
  XNOR2_X1 U787 ( .A(n718), .B(KEYINPUT50), .ZN(n725) );
  NOR2_X1 U788 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U789 ( .A(KEYINPUT49), .B(n721), .Z(n722) );
  NOR2_X1 U790 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U791 ( .A1(n725), .A2(n724), .ZN(n727) );
  NAND2_X1 U792 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U793 ( .A(KEYINPUT51), .B(n728), .ZN(n729) );
  NOR2_X1 U794 ( .A1(n736), .A2(n729), .ZN(n730) );
  NOR2_X1 U795 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U796 ( .A(n732), .B(KEYINPUT52), .ZN(n733) );
  NOR2_X1 U797 ( .A1(n734), .A2(n733), .ZN(n738) );
  NOR2_X1 U798 ( .A1(n736), .A2(n398), .ZN(n737) );
  NOR2_X1 U799 ( .A1(n738), .A2(n737), .ZN(n746) );
  NOR2_X1 U800 ( .A1(n361), .A2(KEYINPUT2), .ZN(n739) );
  XNOR2_X1 U801 ( .A(n739), .B(KEYINPUT80), .ZN(n740) );
  NOR2_X1 U802 ( .A1(n741), .A2(n740), .ZN(n744) );
  INV_X1 U803 ( .A(n671), .ZN(n778) );
  NOR2_X1 U804 ( .A1(n778), .A2(KEYINPUT2), .ZN(n742) );
  XNOR2_X1 U805 ( .A(n742), .B(KEYINPUT79), .ZN(n743) );
  NAND2_X1 U806 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U807 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U808 ( .A1(n747), .A2(G953), .ZN(n748) );
  XNOR2_X1 U809 ( .A(n748), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U810 ( .A1(n381), .A2(G210), .ZN(n753) );
  XOR2_X1 U811 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n751) );
  BUF_X1 U812 ( .A(n749), .Z(n750) );
  XNOR2_X1 U813 ( .A(n753), .B(n752), .ZN(n754) );
  XOR2_X1 U814 ( .A(KEYINPUT56), .B(KEYINPUT119), .Z(n755) );
  XNOR2_X1 U815 ( .A(n756), .B(n755), .ZN(G51) );
  NAND2_X1 U816 ( .A1(n773), .A2(G469), .ZN(n760) );
  XOR2_X1 U817 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n757) );
  XNOR2_X1 U818 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U819 ( .A(n760), .B(n759), .ZN(n761) );
  NOR2_X1 U820 ( .A1(n777), .A2(n761), .ZN(G54) );
  XOR2_X1 U821 ( .A(KEYINPUT120), .B(KEYINPUT59), .Z(n762) );
  XNOR2_X1 U822 ( .A(n765), .B(n764), .ZN(n766) );
  NAND2_X1 U823 ( .A1(n773), .A2(G478), .ZN(n771) );
  INV_X1 U824 ( .A(KEYINPUT121), .ZN(n768) );
  NOR2_X1 U825 ( .A1(n777), .A2(n772), .ZN(G63) );
  NAND2_X1 U826 ( .A1(n773), .A2(G217), .ZN(n775) );
  XNOR2_X1 U827 ( .A(n774), .B(n775), .ZN(n776) );
  NOR2_X1 U828 ( .A1(n777), .A2(n776), .ZN(G66) );
  NAND2_X1 U829 ( .A1(n778), .A2(n797), .ZN(n783) );
  NAND2_X1 U830 ( .A1(G224), .A2(G953), .ZN(n779) );
  XNOR2_X1 U831 ( .A(n779), .B(KEYINPUT122), .ZN(n780) );
  XNOR2_X1 U832 ( .A(KEYINPUT61), .B(n780), .ZN(n781) );
  NAND2_X1 U833 ( .A1(n781), .A2(G898), .ZN(n782) );
  NAND2_X1 U834 ( .A1(n783), .A2(n782), .ZN(n791) );
  XOR2_X1 U835 ( .A(G101), .B(KEYINPUT123), .Z(n784) );
  XNOR2_X1 U836 ( .A(n785), .B(n784), .ZN(n787) );
  XNOR2_X1 U837 ( .A(n786), .B(n787), .ZN(n788) );
  NOR2_X1 U838 ( .A1(n789), .A2(n788), .ZN(n790) );
  XNOR2_X1 U839 ( .A(n791), .B(n790), .ZN(n792) );
  XNOR2_X1 U840 ( .A(KEYINPUT124), .B(n792), .ZN(G69) );
  XNOR2_X1 U841 ( .A(n793), .B(KEYINPUT125), .ZN(n795) );
  XOR2_X1 U842 ( .A(n794), .B(n795), .Z(n800) );
  XNOR2_X1 U843 ( .A(n800), .B(n796), .ZN(n798) );
  NAND2_X1 U844 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U845 ( .A(n799), .B(KEYINPUT126), .ZN(n804) );
  XNOR2_X1 U846 ( .A(G227), .B(n800), .ZN(n801) );
  NAND2_X1 U847 ( .A1(n801), .A2(G900), .ZN(n802) );
  NAND2_X1 U848 ( .A1(n802), .A2(G953), .ZN(n803) );
  NAND2_X1 U849 ( .A1(n804), .A2(n803), .ZN(G72) );
  XOR2_X1 U850 ( .A(G125), .B(KEYINPUT37), .Z(n805) );
  XNOR2_X1 U851 ( .A(n806), .B(n805), .ZN(G27) );
  XNOR2_X1 U852 ( .A(G140), .B(n807), .ZN(G42) );
  XNOR2_X1 U853 ( .A(G131), .B(n808), .ZN(G33) );
  XNOR2_X1 U854 ( .A(G137), .B(n809), .ZN(G39) );
endmodule

