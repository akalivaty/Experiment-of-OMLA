//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 1 0 1 1 1 0 0 1 1 1 1 1 1 1 1 0 1 0 0 0 0 1 0 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 1 1 0 0 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:54 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1329, new_n1330, new_n1331,
    new_n1332, new_n1334, new_n1335, new_n1336, new_n1337, new_n1338,
    new_n1339, new_n1341, new_n1342, new_n1343, new_n1344, new_n1345,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1392, new_n1393, new_n1394, new_n1395,
    new_n1396;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT65), .ZN(new_n214));
  XNOR2_X1  g0014(.A(KEYINPUT64), .B(G20), .ZN(new_n215));
  NAND2_X1  g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n214), .A2(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n219));
  INV_X1    g0019(.A(G77), .ZN(new_n220));
  INV_X1    g0020(.A(G244), .ZN(new_n221));
  INV_X1    g0021(.A(G264), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n220), .B2(new_n221), .C1(new_n206), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n209), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n212), .B(new_n218), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  INV_X1    g0030(.A(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XOR2_X1   g0042(.A(G107), .B(G116), .Z(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  INV_X1    g0045(.A(G33), .ZN(new_n246));
  OAI21_X1  g0046(.A(KEYINPUT66), .B1(new_n209), .B2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(KEYINPUT66), .ZN(new_n248));
  NAND4_X1  g0048(.A1(new_n248), .A2(G1), .A3(G20), .A4(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G1), .ZN(new_n250));
  NAND3_X1  g0050(.A1(new_n250), .A2(G13), .A3(G20), .ZN(new_n251));
  NAND4_X1  g0051(.A1(new_n247), .A2(new_n216), .A3(new_n249), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(G20), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G50), .ZN(new_n254));
  OAI22_X1  g0054(.A1(new_n252), .A2(new_n254), .B1(G50), .B2(new_n251), .ZN(new_n255));
  XNOR2_X1  g0055(.A(KEYINPUT8), .B(G58), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(KEYINPUT67), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT67), .ZN(new_n258));
  INV_X1    g0058(.A(G58), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n259), .A3(KEYINPUT8), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n257), .A2(G33), .A3(new_n215), .A4(new_n260), .ZN(new_n261));
  NOR2_X1   g0061(.A1(G20), .A2(G33), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n247), .A2(new_n216), .A3(new_n249), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n255), .B1(new_n266), .B2(KEYINPUT68), .ZN(new_n267));
  INV_X1    g0067(.A(new_n265), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n261), .B2(new_n263), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT68), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(G33), .ZN(new_n276));
  AND2_X1   g0076(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  NOR2_X1   g0077(.A1(G222), .A2(G1698), .ZN(new_n278));
  INV_X1    g0078(.A(G1698), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G223), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n216), .B1(G33), .B2(G41), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n281), .B(new_n282), .C1(G77), .C2(new_n277), .ZN(new_n283));
  INV_X1    g0083(.A(G41), .ZN(new_n284));
  INV_X1    g0084(.A(G45), .ZN(new_n285));
  AOI21_X1  g0085(.A(G1), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(G33), .A2(G41), .ZN(new_n287));
  NAND3_X1  g0087(.A1(new_n287), .A2(G1), .A3(G13), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n286), .A2(new_n288), .A3(G274), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n285), .ZN(new_n291));
  AND2_X1   g0091(.A1(G1), .A2(G13), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n250), .A2(new_n291), .B1(new_n292), .B2(new_n287), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n290), .B1(G226), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n283), .A2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G179), .B2(new_n295), .ZN(new_n298));
  OR2_X1    g0098(.A1(new_n273), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT10), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n272), .A2(KEYINPUT9), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT9), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n267), .A2(new_n302), .A3(new_n271), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n295), .A2(G200), .ZN(new_n305));
  INV_X1    g0105(.A(G190), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n295), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n300), .B1(new_n304), .B2(new_n308), .ZN(new_n309));
  AOI211_X1 g0109(.A(KEYINPUT10), .B(new_n307), .C1(new_n301), .C2(new_n303), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n299), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT13), .ZN(new_n312));
  INV_X1    g0112(.A(G226), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n279), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n231), .A2(G1698), .ZN(new_n315));
  NAND4_X1  g0115(.A1(new_n274), .A2(new_n314), .A3(new_n276), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n318), .A2(new_n282), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n250), .B1(G41), .B2(G45), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n288), .A2(G238), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g0121(.A1(new_n289), .A2(new_n321), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n312), .B1(new_n319), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n288), .B1(new_n316), .B2(new_n317), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n289), .A2(new_n321), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n324), .A2(new_n325), .A3(KEYINPUT13), .ZN(new_n326));
  OAI21_X1  g0126(.A(G169), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n319), .A2(new_n312), .A3(new_n322), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT71), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n319), .A2(new_n322), .A3(KEYINPUT71), .A4(new_n312), .ZN(new_n332));
  OAI21_X1  g0132(.A(KEYINPUT13), .B1(new_n324), .B2(new_n325), .ZN(new_n333));
  NAND4_X1  g0133(.A1(new_n331), .A2(G179), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(new_n333), .ZN(new_n335));
  INV_X1    g0135(.A(KEYINPUT14), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n335), .A2(new_n336), .A3(G169), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n328), .A2(new_n334), .A3(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G20), .ZN(new_n339));
  OAI21_X1  g0139(.A(KEYINPUT72), .B1(new_n339), .B2(G68), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n246), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n202), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n339), .A2(KEYINPUT64), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT64), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(G20), .ZN(new_n345));
  NAND4_X1  g0145(.A1(new_n343), .A2(new_n345), .A3(G33), .A4(G77), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n262), .A2(KEYINPUT72), .A3(G50), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n342), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n348), .A2(KEYINPUT11), .A3(new_n265), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n251), .A2(G68), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT12), .ZN(new_n351));
  XNOR2_X1  g0151(.A(new_n350), .B(new_n351), .ZN(new_n352));
  AND2_X1   g0152(.A1(new_n349), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(KEYINPUT11), .B1(new_n348), .B2(new_n265), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n253), .A2(G68), .ZN(new_n355));
  NOR2_X1   g0155(.A1(new_n252), .A2(new_n355), .ZN(new_n356));
  NOR2_X1   g0156(.A1(new_n354), .A2(new_n356), .ZN(new_n357));
  AND3_X1   g0157(.A1(new_n353), .A2(new_n357), .A3(KEYINPUT73), .ZN(new_n358));
  AOI21_X1  g0158(.A(KEYINPUT73), .B1(new_n353), .B2(new_n357), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n338), .A2(new_n360), .ZN(new_n361));
  AND2_X1   g0161(.A1(new_n353), .A2(new_n357), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n331), .A2(G190), .A3(new_n332), .A4(new_n333), .ZN(new_n363));
  AND3_X1   g0163(.A1(new_n335), .A2(KEYINPUT70), .A3(G200), .ZN(new_n364));
  AOI21_X1  g0164(.A(KEYINPUT70), .B1(new_n335), .B2(G200), .ZN(new_n365));
  OAI211_X1 g0165(.A(new_n362), .B(new_n363), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n361), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n343), .A2(new_n345), .ZN(new_n369));
  XNOR2_X1  g0169(.A(KEYINPUT15), .B(G87), .ZN(new_n370));
  NOR3_X1   g0170(.A1(new_n369), .A2(new_n370), .A3(new_n246), .ZN(new_n371));
  OAI22_X1  g0171(.A1(new_n220), .A2(new_n215), .B1(new_n256), .B2(new_n341), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n265), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n268), .A2(G77), .A3(new_n251), .A4(new_n253), .ZN(new_n374));
  INV_X1    g0174(.A(new_n251), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n220), .ZN(new_n376));
  AND3_X1   g0176(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT69), .ZN(new_n378));
  INV_X1    g0178(.A(G200), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n290), .B1(G244), .B2(new_n293), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n274), .A2(new_n276), .A3(G238), .A4(G1698), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n274), .A2(new_n276), .A3(G232), .A4(new_n279), .ZN(new_n382));
  OAI211_X1 g0182(.A(new_n381), .B(new_n382), .C1(new_n277), .C2(new_n206), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n282), .ZN(new_n384));
  AND2_X1   g0184(.A1(new_n380), .A2(new_n384), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n377), .B(new_n378), .C1(new_n379), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(G190), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n379), .B1(new_n380), .B2(new_n384), .ZN(new_n388));
  NAND3_X1  g0188(.A1(new_n373), .A2(new_n374), .A3(new_n376), .ZN(new_n389));
  OAI21_X1  g0189(.A(KEYINPUT69), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n386), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G179), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n385), .A2(new_n392), .ZN(new_n393));
  OAI211_X1 g0193(.A(new_n393), .B(new_n389), .C1(G169), .C2(new_n385), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n391), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n368), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n311), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT18), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n257), .A2(new_n260), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(new_n375), .ZN(new_n400));
  NAND3_X1  g0200(.A1(new_n257), .A2(new_n260), .A3(new_n253), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n400), .B1(new_n252), .B2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(KEYINPUT75), .B1(new_n275), .B2(G33), .ZN(new_n404));
  INV_X1    g0204(.A(KEYINPUT75), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n405), .A2(new_n246), .A3(KEYINPUT3), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n404), .A2(new_n406), .A3(new_n276), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(new_n215), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT7), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n274), .A2(new_n276), .ZN(new_n410));
  NOR2_X1   g0210(.A1(KEYINPUT7), .A2(G20), .ZN(new_n411));
  AND2_X1   g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n409), .A2(G68), .A3(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(G68), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n259), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G20), .B1(new_n416), .B2(new_n201), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n262), .A2(G159), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT16), .B1(new_n414), .B2(new_n420), .ZN(new_n421));
  AND3_X1   g0221(.A1(new_n417), .A2(KEYINPUT16), .A3(new_n418), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT7), .ZN(new_n423));
  AND3_X1   g0223(.A1(new_n246), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n424));
  AOI21_X1  g0224(.A(KEYINPUT74), .B1(new_n246), .B2(KEYINPUT3), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n276), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n423), .B1(new_n426), .B2(new_n339), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n246), .A2(KEYINPUT3), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT74), .ZN(new_n429));
  OAI21_X1  g0229(.A(new_n429), .B1(new_n275), .B2(G33), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n246), .A2(KEYINPUT74), .A3(KEYINPUT3), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n428), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n343), .A2(new_n345), .A3(new_n423), .ZN(new_n433));
  OAI21_X1  g0233(.A(G68), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n422), .B1(new_n427), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n435), .A2(new_n265), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n403), .B1(new_n421), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n288), .A2(new_n320), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n289), .B1(new_n231), .B2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(G87), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n246), .A2(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n313), .A2(G1698), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G223), .B2(G1698), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n442), .B1(new_n426), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n439), .B1(new_n445), .B2(new_n282), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT76), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n446), .A2(new_n447), .A3(new_n392), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n445), .A2(new_n282), .ZN(new_n449));
  INV_X1    g0249(.A(G274), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n292), .B2(new_n287), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n293), .A2(G232), .B1(new_n451), .B2(new_n286), .ZN(new_n452));
  AOI21_X1  g0252(.A(G169), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(G223), .A2(G1698), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n454), .B1(new_n313), .B2(G1698), .ZN(new_n455));
  AOI21_X1  g0255(.A(new_n441), .B1(new_n432), .B2(new_n455), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n452), .B(new_n392), .C1(new_n456), .C2(new_n288), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(KEYINPUT76), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n448), .B1(new_n453), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n398), .B1(new_n437), .B2(new_n459), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT16), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n423), .B1(new_n407), .B2(new_n215), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n463), .A2(new_n415), .A3(new_n412), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(new_n419), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT7), .B1(new_n432), .B2(G20), .ZN(new_n466));
  INV_X1    g0266(.A(new_n433), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n426), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n466), .A2(new_n468), .A3(G68), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n268), .B1(new_n469), .B2(new_n422), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n465), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT77), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n446), .A2(new_n472), .A3(new_n306), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n452), .B(new_n306), .C1(new_n456), .C2(new_n288), .ZN(new_n474));
  OAI211_X1 g0274(.A(KEYINPUT77), .B(new_n474), .C1(new_n446), .C2(G200), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n471), .A2(new_n403), .A3(new_n473), .A4(new_n475), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT17), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n437), .A2(new_n459), .A3(new_n398), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n474), .A2(KEYINPUT77), .ZN(new_n480));
  AOI21_X1  g0280(.A(new_n472), .B1(new_n446), .B2(new_n306), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n456), .A2(new_n288), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n379), .B1(new_n482), .B2(new_n439), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n402), .B1(new_n465), .B2(new_n470), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n484), .A2(KEYINPUT17), .A3(new_n485), .ZN(new_n486));
  NAND4_X1  g0286(.A1(new_n461), .A2(new_n478), .A3(new_n479), .A4(new_n486), .ZN(new_n487));
  OR2_X1    g0287(.A1(new_n487), .A2(KEYINPUT78), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(KEYINPUT78), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n397), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  NOR2_X1   g0290(.A1(new_n251), .A2(G97), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n246), .A2(G1), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n252), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(G97), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n463), .A2(new_n206), .A3(new_n412), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT6), .ZN(new_n497));
  NOR3_X1   g0297(.A1(new_n497), .A2(new_n205), .A3(G107), .ZN(new_n498));
  XNOR2_X1  g0298(.A(G97), .B(G107), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n498), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n500), .A2(new_n215), .B1(new_n220), .B2(new_n341), .ZN(new_n501));
  OR2_X1    g0301(.A1(new_n496), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n495), .B1(new_n502), .B2(new_n265), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n274), .A2(new_n276), .A3(G250), .A4(G1698), .ZN(new_n504));
  AND2_X1   g0304(.A1(KEYINPUT4), .A2(G244), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n274), .A2(new_n276), .A3(new_n505), .A4(new_n279), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G283), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n221), .A2(G1698), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n276), .B(new_n509), .C1(new_n424), .C2(new_n425), .ZN(new_n510));
  XNOR2_X1  g0310(.A(KEYINPUT79), .B(KEYINPUT4), .ZN(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT80), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n508), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n511), .B1(new_n432), .B2(new_n509), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(KEYINPUT80), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n288), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n250), .A2(G45), .ZN(new_n519));
  OR2_X1    g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  NAND2_X1  g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n522), .A2(new_n282), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(G257), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n451), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(G200), .B1(new_n518), .B2(new_n526), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n504), .A2(new_n506), .A3(new_n507), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n516), .B2(KEYINPUT80), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n513), .A2(new_n514), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n282), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g0331(.A(new_n526), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n531), .A2(G190), .A3(new_n532), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n503), .A2(new_n527), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n296), .B1(new_n518), .B2(new_n526), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n392), .A3(new_n532), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n496), .A2(new_n501), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n494), .B1(new_n537), .B2(new_n268), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n535), .A2(new_n536), .A3(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n534), .A2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT81), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n541), .B1(new_n285), .B2(G1), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n250), .A2(KEYINPUT81), .A3(G45), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n288), .A2(new_n542), .A3(G250), .A4(new_n543), .ZN(new_n544));
  NOR2_X1   g0344(.A1(new_n285), .A2(G1), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n288), .A2(G274), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT82), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n544), .A2(KEYINPUT82), .A3(new_n546), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n221), .A2(G1698), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(G238), .B2(G1698), .ZN(new_n552));
  OR2_X1    g0352(.A1(KEYINPUT83), .A2(G116), .ZN(new_n553));
  NAND2_X1  g0353(.A1(KEYINPUT83), .A2(G116), .ZN(new_n554));
  AND2_X1   g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI22_X1  g0355(.A1(new_n426), .A2(new_n552), .B1(new_n246), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n549), .A2(new_n550), .B1(new_n556), .B2(new_n282), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT84), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n557), .A2(new_n558), .A3(new_n392), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n215), .A2(G33), .A3(G97), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT19), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n432), .A2(G68), .A3(new_n215), .ZN(new_n563));
  NAND3_X1  g0363(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n343), .A2(new_n345), .A3(KEYINPUT85), .A4(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n565), .B1(G87), .B2(new_n207), .ZN(new_n566));
  AOI21_X1  g0366(.A(KEYINPUT85), .B1(new_n215), .B2(new_n564), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n562), .B(new_n563), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(new_n265), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n370), .A2(new_n375), .ZN(new_n570));
  OR3_X1    g0370(.A1(new_n252), .A2(new_n370), .A3(new_n492), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n544), .A2(KEYINPUT82), .A3(new_n546), .ZN(new_n573));
  AOI21_X1  g0373(.A(KEYINPUT82), .B1(new_n544), .B2(new_n546), .ZN(new_n574));
  NOR2_X1   g0374(.A1(G238), .A2(G1698), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n575), .B1(new_n221), .B2(G1698), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n553), .A2(new_n554), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n432), .A2(new_n576), .B1(G33), .B2(new_n577), .ZN(new_n578));
  OAI22_X1  g0378(.A1(new_n573), .A2(new_n574), .B1(new_n578), .B2(new_n288), .ZN(new_n579));
  OAI21_X1  g0379(.A(KEYINPUT84), .B1(new_n579), .B2(G179), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n579), .A2(new_n296), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n559), .A2(new_n572), .A3(new_n580), .A4(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT86), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n579), .B2(new_n306), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n549), .A2(new_n550), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n556), .A2(new_n282), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT86), .A4(G190), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n579), .A2(G200), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n568), .A2(new_n265), .B1(new_n375), .B2(new_n370), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n493), .A2(G87), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n589), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n582), .B1(new_n588), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n540), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n523), .A2(G270), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(new_n525), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT87), .ZN(new_n597));
  INV_X1    g0397(.A(G257), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(G1698), .ZN(new_n599));
  AOI21_X1  g0399(.A(new_n597), .B1(new_n432), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n432), .A2(new_n597), .A3(new_n599), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n410), .A2(G303), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n222), .A2(new_n279), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n432), .A2(new_n604), .ZN(new_n605));
  NAND4_X1  g0405(.A1(new_n601), .A2(new_n602), .A3(new_n603), .A4(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n596), .B1(new_n606), .B2(new_n282), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n577), .A2(new_n251), .ZN(new_n608));
  INV_X1    g0408(.A(G116), .ZN(new_n609));
  NOR3_X1   g0409(.A1(new_n252), .A2(new_n609), .A3(new_n492), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n246), .A2(G97), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n215), .A2(new_n507), .A3(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n553), .A2(G20), .A3(new_n554), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n265), .A3(new_n613), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT20), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND4_X1  g0416(.A1(new_n612), .A2(new_n265), .A3(KEYINPUT20), .A4(new_n613), .ZN(new_n617));
  AOI211_X1 g0417(.A(new_n608), .B(new_n610), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n607), .B1(new_n618), .B2(new_n392), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n602), .A2(new_n603), .A3(new_n605), .ZN(new_n620));
  OAI21_X1  g0420(.A(new_n282), .B1(new_n620), .B2(new_n600), .ZN(new_n621));
  INV_X1    g0421(.A(new_n596), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(KEYINPUT21), .A2(G169), .ZN(new_n624));
  OAI21_X1  g0424(.A(new_n623), .B1(new_n618), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n619), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(KEYINPUT21), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n623), .A2(G169), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n618), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n621), .A2(G190), .A3(new_n622), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n630), .B(new_n618), .C1(new_n607), .C2(new_n379), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n626), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n521), .ZN(new_n633));
  NOR2_X1   g0433(.A1(KEYINPUT5), .A2(G41), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n545), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(G264), .A3(new_n288), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n636), .A2(new_n525), .ZN(new_n637));
  NOR2_X1   g0437(.A1(G250), .A2(G1698), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n638), .B1(new_n598), .B2(G1698), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n432), .A2(new_n639), .B1(G33), .B2(G294), .ZN(new_n640));
  OAI211_X1 g0440(.A(new_n637), .B(KEYINPUT90), .C1(new_n288), .C2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(KEYINPUT90), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n432), .A2(new_n639), .ZN(new_n643));
  NAND2_X1  g0443(.A1(G33), .A2(G294), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n288), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n636), .A2(new_n525), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n641), .A2(new_n647), .A3(G169), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n637), .B(G179), .C1(new_n288), .C2(new_n640), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n432), .A2(KEYINPUT22), .A3(G87), .A4(new_n215), .ZN(new_n651));
  INV_X1    g0451(.A(KEYINPUT22), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n343), .A2(new_n345), .A3(G87), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n652), .B1(new_n653), .B2(new_n410), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n577), .A2(new_n339), .A3(G33), .ZN(new_n655));
  NOR2_X1   g0455(.A1(KEYINPUT23), .A2(G107), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n206), .A2(G20), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n369), .A2(new_n656), .B1(KEYINPUT23), .B2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n651), .A2(new_n654), .A3(new_n655), .A4(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT24), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n658), .A2(new_n655), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n662), .A2(KEYINPUT24), .A3(new_n651), .A4(new_n654), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n661), .A2(new_n663), .A3(new_n265), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n375), .A2(new_n206), .ZN(new_n665));
  INV_X1    g0465(.A(KEYINPUT25), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n667), .A2(KEYINPUT89), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT89), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n665), .A2(new_n669), .A3(new_n666), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT88), .B1(new_n665), .B2(new_n666), .ZN(new_n671));
  OR4_X1    g0471(.A1(KEYINPUT88), .A2(new_n251), .A3(new_n666), .A4(G107), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n668), .A2(new_n670), .A3(new_n671), .A4(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n493), .A2(G107), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n664), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n650), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g0477(.A(G190), .B1(new_n641), .B2(new_n647), .ZN(new_n678));
  OAI211_X1 g0478(.A(new_n525), .B(new_n636), .C1(new_n640), .C2(new_n288), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n679), .A2(new_n379), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n664), .B(new_n675), .C1(new_n678), .C2(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n677), .A2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n632), .A2(new_n682), .ZN(new_n683));
  AND3_X1   g0483(.A1(new_n490), .A2(new_n594), .A3(new_n683), .ZN(G372));
  INV_X1    g0484(.A(new_n394), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n366), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n361), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n446), .A2(G200), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n474), .A2(KEYINPUT77), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n473), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NOR3_X1   g0490(.A1(new_n437), .A2(new_n690), .A3(new_n477), .ZN(new_n691));
  AOI21_X1  g0491(.A(KEYINPUT17), .B1(new_n484), .B2(new_n485), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n687), .A2(new_n693), .ZN(new_n694));
  AND3_X1   g0494(.A1(new_n437), .A2(new_n459), .A3(new_n398), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(new_n460), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g0497(.A1(new_n309), .A2(new_n310), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n299), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n490), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT26), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT91), .B1(new_n557), .B2(G169), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n557), .A2(new_n392), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT91), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n579), .A2(new_n706), .A3(new_n296), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n704), .A2(new_n572), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n588), .B2(new_n592), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n703), .B1(new_n709), .B2(new_n539), .ZN(new_n710));
  INV_X1    g0510(.A(new_n539), .ZN(new_n711));
  AND2_X1   g0511(.A1(new_n590), .A2(new_n591), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n584), .A2(new_n587), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n712), .A2(new_n713), .A3(new_n589), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n711), .A2(KEYINPUT26), .A3(new_n714), .A4(new_n582), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n710), .A2(new_n715), .ZN(new_n716));
  AND3_X1   g0516(.A1(new_n714), .A2(new_n681), .A3(new_n708), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n534), .A2(new_n539), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n626), .A2(new_n629), .A3(new_n677), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n717), .A2(new_n718), .A3(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n716), .A2(new_n720), .A3(new_n708), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n701), .B1(new_n702), .B2(new_n722), .ZN(G369));
  NAND2_X1  g0523(.A1(new_n626), .A2(new_n629), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n215), .A2(new_n250), .A3(G13), .ZN(new_n725));
  OR2_X1    g0525(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(KEYINPUT27), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(G213), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(G343), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n618), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(new_n632), .B2(new_n732), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n734), .A2(G330), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n677), .A2(new_n731), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT92), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n731), .B1(new_n664), .B2(new_n675), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n738), .B1(new_n682), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n736), .A2(new_n740), .ZN(new_n741));
  XOR2_X1   g0541(.A(new_n741), .B(KEYINPUT93), .Z(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n724), .A2(new_n731), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n677), .ZN(new_n746));
  AOI22_X1  g0546(.A1(new_n740), .A2(new_n745), .B1(new_n746), .B2(new_n731), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n743), .A2(new_n747), .ZN(G399));
  INV_X1    g0548(.A(new_n210), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n749), .A2(G41), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR3_X1   g0551(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n751), .A2(G1), .A3(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n214), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n753), .B1(new_n754), .B2(new_n751), .ZN(new_n755));
  XOR2_X1   g0555(.A(KEYINPUT94), .B(KEYINPUT28), .Z(new_n756));
  XNOR2_X1  g0556(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n645), .A2(new_n646), .A3(new_n392), .ZN(new_n758));
  NAND4_X1  g0558(.A1(new_n758), .A2(new_n621), .A3(new_n557), .A4(new_n595), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n531), .A2(new_n532), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT95), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n585), .A2(new_n586), .A3(new_n595), .ZN(new_n762));
  NOR2_X1   g0562(.A1(new_n762), .A2(new_n649), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n513), .A2(new_n514), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n764), .A2(new_n517), .A3(new_n528), .ZN(new_n765));
  AOI21_X1  g0565(.A(new_n526), .B1(new_n765), .B2(new_n282), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT95), .ZN(new_n767));
  NAND4_X1  g0567(.A1(new_n763), .A2(new_n766), .A3(new_n767), .A4(new_n621), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT30), .ZN(new_n769));
  AND3_X1   g0569(.A1(new_n761), .A2(new_n768), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(KEYINPUT96), .ZN(new_n771));
  AOI21_X1  g0571(.A(G179), .B1(new_n585), .B2(new_n586), .ZN(new_n772));
  NAND3_X1  g0572(.A1(new_n623), .A2(new_n679), .A3(new_n772), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n771), .B1(new_n773), .B2(new_n766), .ZN(new_n774));
  AND3_X1   g0574(.A1(new_n579), .A2(new_n392), .A3(new_n679), .ZN(new_n775));
  NAND4_X1  g0575(.A1(new_n760), .A2(new_n775), .A3(KEYINPUT96), .A4(new_n623), .ZN(new_n776));
  NAND4_X1  g0576(.A1(new_n763), .A2(new_n766), .A3(KEYINPUT30), .A4(new_n621), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n730), .B1(new_n770), .B2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(KEYINPUT31), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  NOR3_X1   g0581(.A1(new_n540), .A2(new_n593), .A3(new_n730), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(new_n683), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n731), .A2(new_n780), .ZN(new_n784));
  OAI21_X1  g0584(.A(new_n777), .B1(new_n766), .B2(new_n773), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n770), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n781), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G330), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  INV_X1    g0589(.A(KEYINPUT29), .ZN(new_n790));
  NAND3_X1  g0590(.A1(new_n721), .A2(new_n790), .A3(new_n731), .ZN(new_n791));
  INV_X1    g0591(.A(new_n708), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n714), .A2(new_n681), .A3(new_n708), .ZN(new_n793));
  NOR2_X1   g0593(.A1(new_n793), .A2(new_n540), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n792), .B1(new_n794), .B2(new_n719), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT26), .B1(new_n709), .B2(new_n539), .ZN(new_n796));
  NAND4_X1  g0596(.A1(new_n711), .A2(new_n703), .A3(new_n714), .A4(new_n582), .ZN(new_n797));
  AND2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n730), .B1(new_n795), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n791), .B1(new_n799), .B2(new_n790), .ZN(new_n800));
  OR2_X1    g0600(.A1(new_n789), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n757), .B1(new_n802), .B2(G1), .ZN(G364));
  INV_X1    g0603(.A(G13), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n369), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(G45), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(G1), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(new_n750), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n277), .A2(new_n210), .ZN(new_n809));
  INV_X1    g0609(.A(G355), .ZN(new_n810));
  OAI22_X1  g0610(.A1(new_n809), .A2(new_n810), .B1(G116), .B2(new_n210), .ZN(new_n811));
  OR2_X1    g0611(.A1(new_n241), .A2(new_n285), .ZN(new_n812));
  NOR2_X1   g0612(.A1(new_n432), .A2(new_n749), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n814), .B1(new_n285), .B2(new_n214), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n811), .B1(new_n812), .B2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(G13), .A2(G33), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(G20), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n216), .B1(G20), .B2(new_n296), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n808), .B1(new_n816), .B2(new_n822), .ZN(new_n823));
  XOR2_X1   g0623(.A(new_n823), .B(KEYINPUT97), .Z(new_n824));
  INV_X1    g0624(.A(G303), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n379), .A2(G179), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n826), .A2(G20), .A3(G190), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n369), .A2(new_n306), .A3(new_n826), .ZN(new_n828));
  INV_X1    g0628(.A(G283), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n410), .B1(new_n825), .B2(new_n827), .C1(new_n828), .C2(new_n829), .ZN(new_n830));
  NOR2_X1   g0630(.A1(G179), .A2(G200), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n215), .B1(G190), .B2(new_n831), .ZN(new_n832));
  INV_X1    g0632(.A(G294), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n369), .A2(new_n306), .A3(new_n831), .ZN(new_n834));
  INV_X1    g0634(.A(G329), .ZN(new_n835));
  OAI22_X1  g0635(.A1(new_n832), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OR3_X1    g0636(.A1(new_n215), .A2(KEYINPUT98), .A3(new_n392), .ZN(new_n837));
  OAI21_X1  g0637(.A(KEYINPUT98), .B1(new_n215), .B2(new_n392), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n839), .A2(G190), .A3(new_n379), .ZN(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n830), .B(new_n836), .C1(new_n841), .C2(G322), .ZN(new_n842));
  AOI211_X1 g0642(.A(new_n306), .B(new_n379), .C1(new_n837), .C2(new_n838), .ZN(new_n843));
  XOR2_X1   g0643(.A(KEYINPUT102), .B(G326), .Z(new_n844));
  NAND2_X1  g0644(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n839), .A2(new_n306), .A3(new_n379), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n847), .A2(G311), .ZN(new_n848));
  AOI211_X1 g0648(.A(G190), .B(new_n379), .C1(new_n837), .C2(new_n838), .ZN(new_n849));
  XNOR2_X1  g0649(.A(KEYINPUT33), .B(G317), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n842), .A2(new_n845), .A3(new_n848), .A4(new_n851), .ZN(new_n852));
  OAI22_X1  g0652(.A1(new_n259), .A2(new_n840), .B1(new_n846), .B2(new_n220), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n853), .A2(KEYINPUT99), .B1(G50), .B2(new_n843), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n854), .B1(KEYINPUT99), .B2(new_n853), .ZN(new_n855));
  XNOR2_X1  g0655(.A(new_n855), .B(KEYINPUT100), .ZN(new_n856));
  INV_X1    g0656(.A(new_n834), .ZN(new_n857));
  XOR2_X1   g0657(.A(KEYINPUT101), .B(G159), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  XOR2_X1   g0659(.A(new_n859), .B(KEYINPUT32), .Z(new_n860));
  INV_X1    g0660(.A(new_n828), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(G107), .ZN(new_n862));
  INV_X1    g0662(.A(new_n827), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n863), .A2(G87), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n277), .A3(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n832), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n865), .B1(G97), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n849), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n860), .B(new_n867), .C1(new_n415), .C2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n852), .B1(new_n856), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n824), .B1(new_n870), .B2(new_n820), .ZN(new_n871));
  INV_X1    g0671(.A(new_n819), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n871), .B1(new_n734), .B2(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n736), .A2(new_n808), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(G330), .B2(new_n734), .ZN(new_n875));
  AND2_X1   g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(G396));
  NOR2_X1   g0677(.A1(new_n394), .A2(new_n730), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n730), .A2(new_n389), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n391), .A2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n878), .B1(new_n880), .B2(new_n394), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n881), .B(KEYINPUT103), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n722), .B2(new_n730), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n395), .A2(new_n731), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n721), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n883), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n789), .ZN(new_n888));
  INV_X1    g0688(.A(new_n808), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n883), .A2(new_n788), .A3(new_n886), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(G294), .A2(new_n841), .B1(new_n847), .B2(new_n577), .ZN(new_n892));
  OAI21_X1  g0692(.A(new_n892), .B1(new_n829), .B2(new_n868), .ZN(new_n893));
  INV_X1    g0693(.A(new_n843), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n894), .A2(new_n825), .ZN(new_n895));
  OAI221_X1 g0695(.A(new_n410), .B1(new_n206), .B2(new_n827), .C1(new_n832), .C2(new_n205), .ZN(new_n896));
  INV_X1    g0696(.A(G311), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n440), .A2(new_n828), .B1(new_n834), .B2(new_n897), .ZN(new_n898));
  NOR4_X1   g0698(.A1(new_n893), .A2(new_n895), .A3(new_n896), .A4(new_n898), .ZN(new_n899));
  AOI22_X1  g0699(.A1(G143), .A2(new_n841), .B1(new_n847), .B2(new_n858), .ZN(new_n900));
  INV_X1    g0700(.A(G137), .ZN(new_n901));
  INV_X1    g0701(.A(G150), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n900), .B1(new_n901), .B2(new_n894), .C1(new_n902), .C2(new_n868), .ZN(new_n903));
  XNOR2_X1  g0703(.A(new_n903), .B(KEYINPUT34), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n828), .A2(new_n415), .ZN(new_n905));
  OAI221_X1 g0705(.A(new_n432), .B1(new_n202), .B2(new_n827), .C1(new_n832), .C2(new_n259), .ZN(new_n906));
  AOI211_X1 g0706(.A(new_n905), .B(new_n906), .C1(G132), .C2(new_n857), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n899), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(new_n820), .ZN(new_n909));
  NOR2_X1   g0709(.A1(new_n820), .A2(new_n817), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  OAI22_X1  g0711(.A1(new_n908), .A2(new_n909), .B1(G77), .B2(new_n911), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n881), .A2(new_n818), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n808), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n891), .A2(new_n914), .ZN(new_n915));
  AND2_X1   g0715(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n916));
  NOR2_X1   g0716(.A1(new_n915), .A2(KEYINPUT104), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  INV_X1    g0718(.A(new_n918), .ZN(G384));
  NOR2_X1   g0719(.A1(new_n805), .A2(new_n250), .ZN(new_n920));
  INV_X1    g0720(.A(new_n728), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n415), .B1(new_n426), .B2(new_n467), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n419), .B1(new_n922), .B2(new_n466), .ZN(new_n923));
  OAI211_X1 g0723(.A(new_n265), .B(new_n435), .C1(new_n923), .C2(KEYINPUT16), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n403), .ZN(new_n925));
  AOI21_X1  g0725(.A(KEYINPUT106), .B1(new_n924), .B2(new_n403), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n487), .A2(new_n921), .A3(new_n927), .ZN(new_n928));
  INV_X1    g0728(.A(KEYINPUT37), .ZN(new_n929));
  INV_X1    g0729(.A(new_n476), .ZN(new_n930));
  AOI21_X1  g0730(.A(new_n930), .B1(new_n927), .B2(new_n459), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT16), .B1(new_n469), .B2(new_n420), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n403), .B1(new_n436), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(KEYINPUT106), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n924), .A2(KEYINPUT106), .A3(new_n403), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n921), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n929), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n437), .A2(new_n459), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n437), .A2(new_n921), .ZN(new_n940));
  AND4_X1   g0740(.A1(new_n929), .A2(new_n939), .A3(new_n940), .A4(new_n476), .ZN(new_n941));
  OAI211_X1 g0741(.A(KEYINPUT38), .B(new_n928), .C1(new_n938), .C2(new_n941), .ZN(new_n942));
  XOR2_X1   g0742(.A(KEYINPUT108), .B(KEYINPUT39), .Z(new_n943));
  NAND3_X1  g0743(.A1(new_n939), .A2(new_n940), .A3(new_n476), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(KEYINPUT37), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT107), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n939), .A2(new_n940), .A3(new_n476), .A4(new_n929), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n946), .B1(new_n945), .B2(new_n947), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n940), .B1(new_n693), .B2(new_n696), .ZN(new_n950));
  NOR3_X1   g0750(.A1(new_n948), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  OAI211_X1 g0751(.A(new_n942), .B(new_n943), .C1(new_n951), .C2(KEYINPUT38), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n935), .A2(new_n459), .A3(new_n936), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n937), .A2(new_n953), .A3(new_n476), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n954), .A2(KEYINPUT37), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n947), .ZN(new_n956));
  AOI21_X1  g0756(.A(KEYINPUT38), .B1(new_n956), .B2(new_n928), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n941), .B1(new_n954), .B2(KEYINPUT37), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n937), .B1(new_n693), .B2(new_n696), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT38), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n958), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT39), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n952), .A2(new_n962), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n361), .A2(new_n730), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n960), .B1(new_n958), .B2(new_n959), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n942), .A2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n358), .ZN(new_n968));
  INV_X1    g0768(.A(new_n359), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n968), .A2(new_n969), .A3(new_n730), .ZN(new_n970));
  AND3_X1   g0770(.A1(new_n361), .A2(new_n366), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n970), .B1(new_n361), .B2(new_n366), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT105), .ZN(new_n975));
  INV_X1    g0775(.A(new_n878), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n975), .B1(new_n886), .B2(new_n976), .ZN(new_n977));
  AOI211_X1 g0777(.A(KEYINPUT105), .B(new_n878), .C1(new_n721), .C2(new_n885), .ZN(new_n978));
  OAI211_X1 g0778(.A(new_n967), .B(new_n974), .C1(new_n977), .C2(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n728), .B1(new_n695), .B2(new_n460), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n965), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n700), .B1(new_n800), .B2(new_n490), .ZN(new_n982));
  XNOR2_X1  g0782(.A(new_n981), .B(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(G330), .ZN(new_n984));
  INV_X1    g0784(.A(KEYINPUT109), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n945), .A2(new_n947), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT107), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n945), .A2(new_n946), .A3(new_n947), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n487), .A2(new_n437), .A3(new_n921), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n987), .A2(new_n988), .A3(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n961), .B1(new_n960), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n881), .B1(new_n971), .B2(new_n972), .ZN(new_n992));
  INV_X1    g0792(.A(new_n992), .ZN(new_n993));
  AND2_X1   g0793(.A1(new_n777), .A2(new_n776), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n761), .A2(new_n768), .A3(new_n769), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n994), .A2(new_n995), .A3(new_n774), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n996), .A2(new_n784), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n783), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g0798(.A(KEYINPUT31), .B1(new_n996), .B2(new_n730), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n993), .B(KEYINPUT40), .C1(new_n998), .C2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n985), .B1(new_n991), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n942), .B1(new_n951), .B2(KEYINPUT38), .ZN(new_n1002));
  INV_X1    g0802(.A(KEYINPUT40), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n782), .A2(new_n683), .B1(new_n996), .B2(new_n784), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n1003), .B(new_n992), .C1(new_n1004), .C2(new_n781), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1002), .A2(new_n1005), .A3(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n781), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1007), .B(new_n993), .C1(new_n957), .C2(new_n961), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n1001), .A2(new_n1006), .B1(new_n1003), .B2(new_n1008), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n490), .A2(new_n1007), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n984), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n1011), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n920), .B1(new_n983), .B2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1013), .B1(new_n983), .B2(new_n1012), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n500), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT35), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(KEYINPUT35), .ZN(new_n1017));
  NAND4_X1  g0817(.A1(new_n1016), .A2(G116), .A3(new_n217), .A4(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT36), .ZN(new_n1019));
  NOR3_X1   g0819(.A1(new_n754), .A2(new_n220), .A3(new_n416), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n415), .A2(G50), .ZN(new_n1021));
  OAI211_X1 g0821(.A(G1), .B(new_n804), .C1(new_n1020), .C2(new_n1021), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1014), .A2(new_n1019), .A3(new_n1022), .ZN(G367));
  NOR2_X1   g0823(.A1(new_n712), .A2(new_n731), .ZN(new_n1024));
  MUX2_X1   g0824(.A(new_n709), .B(new_n708), .S(new_n1024), .Z(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT110), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n819), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n277), .B1(new_n259), .B2(new_n827), .C1(new_n832), .C2(new_n415), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n861), .A2(G77), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n901), .B2(new_n834), .ZN(new_n1030));
  AOI211_X1 g0830(.A(new_n1028), .B(new_n1030), .C1(new_n849), .C2(new_n858), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G50), .A2(new_n847), .B1(new_n841), .B2(G150), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n843), .A2(G143), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n849), .A2(G294), .ZN(new_n1035));
  AND3_X1   g0835(.A1(new_n863), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1036));
  AOI21_X1  g0836(.A(KEYINPUT46), .B1(new_n863), .B2(new_n577), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1036), .A2(new_n1037), .A3(new_n432), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n861), .A2(G97), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(new_n866), .A2(G107), .B1(new_n857), .B2(G317), .ZN(new_n1040));
  NAND4_X1  g0840(.A1(new_n1035), .A2(new_n1038), .A3(new_n1039), .A4(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n841), .A2(G303), .B1(G311), .B2(new_n843), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n829), .B2(new_n846), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1034), .B1(new_n1041), .B2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g0844(.A(new_n1044), .B(KEYINPUT47), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1045), .A2(new_n820), .ZN(new_n1046));
  OAI221_X1 g0846(.A(new_n821), .B1(new_n210), .B2(new_n370), .C1(new_n237), .C2(new_n814), .ZN(new_n1047));
  NAND4_X1  g0847(.A1(new_n1027), .A2(new_n808), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT114), .ZN(new_n1049));
  INV_X1    g0849(.A(KEYINPUT43), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1026), .A2(new_n1050), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1026), .A2(new_n1050), .ZN(new_n1052));
  OAI21_X1  g0852(.A(new_n718), .B1(new_n503), .B2(new_n731), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n539), .B2(new_n731), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT111), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n740), .A2(new_n745), .ZN(new_n1056));
  INV_X1    g0856(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT42), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1055), .A2(new_n746), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n730), .B1(new_n1060), .B2(new_n539), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n1051), .B(new_n1052), .C1(new_n1059), .C2(new_n1061), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT42), .ZN(new_n1063));
  XNOR2_X1  g0863(.A(new_n1058), .B(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1061), .ZN(new_n1065));
  NAND4_X1  g0865(.A1(new_n1064), .A2(new_n1050), .A3(new_n1026), .A4(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  XOR2_X1   g0867(.A(new_n1054), .B(KEYINPUT111), .Z(new_n1068));
  NOR2_X1   g0868(.A1(new_n743), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1067), .A2(new_n1070), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1062), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n750), .B(KEYINPUT41), .Z(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n740), .A2(new_n745), .ZN(new_n1077));
  OR2_X1    g0877(.A1(new_n1057), .A2(new_n1077), .ZN(new_n1078));
  XOR2_X1   g0878(.A(new_n735), .B(KEYINPUT113), .Z(new_n1079));
  OR2_X1    g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1078), .B1(KEYINPUT113), .B2(new_n735), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n802), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1055), .A2(new_n747), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT45), .ZN(new_n1084));
  XNOR2_X1  g0884(.A(new_n1083), .B(new_n1084), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n747), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n1087));
  OR2_X1    g0887(.A1(KEYINPUT112), .A2(KEYINPUT44), .ZN(new_n1088));
  NAND4_X1  g0888(.A1(new_n1086), .A2(new_n1068), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1089));
  OAI211_X1 g0889(.A(KEYINPUT112), .B(KEYINPUT44), .C1(new_n1055), .C2(new_n747), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1085), .A2(new_n742), .A3(new_n1089), .A4(new_n1090), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT45), .B1(new_n1055), .B2(new_n747), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1089), .B(new_n1090), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n743), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1082), .B1(new_n1091), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1076), .B1(new_n1096), .B2(new_n801), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n807), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1049), .B1(new_n1074), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(G387));
  NAND2_X1  g0901(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1102), .A2(new_n801), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1103), .A2(new_n750), .A3(new_n1082), .ZN(new_n1104));
  OAI22_X1  g0904(.A1(new_n809), .A2(new_n752), .B1(G107), .B2(new_n210), .ZN(new_n1105));
  OR2_X1    g0905(.A1(new_n234), .A2(new_n285), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n752), .ZN(new_n1107));
  AOI211_X1 g0907(.A(G45), .B(new_n1107), .C1(G68), .C2(G77), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n256), .A2(G50), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1109), .B(KEYINPUT50), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n814), .B1(new_n1108), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1105), .B1(new_n1106), .B2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n808), .B1(new_n1112), .B2(new_n822), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G303), .A2(new_n847), .B1(new_n841), .B2(G317), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1114), .A2(KEYINPUT116), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(G311), .A2(new_n849), .B1(new_n843), .B2(G322), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT48), .ZN(new_n1119));
  OR2_X1    g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1121));
  AOI22_X1  g0921(.A1(new_n866), .A2(G283), .B1(new_n863), .B2(G294), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(KEYINPUT49), .ZN(new_n1124));
  OR2_X1    g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1126));
  OAI21_X1  g0926(.A(new_n426), .B1(new_n828), .B2(new_n555), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n857), .B2(new_n844), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1125), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n426), .B1(G77), .B2(new_n863), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1039), .A2(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n832), .A2(new_n370), .B1(new_n834), .B2(new_n902), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1131), .B(new_n1132), .C1(new_n847), .C2(G68), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n841), .A2(G50), .B1(G159), .B2(new_n843), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1133), .B(new_n1134), .C1(new_n399), .C2(new_n868), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1113), .B1(new_n1136), .B2(new_n820), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT117), .ZN(new_n1138));
  OR2_X1    g0938(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1137), .A2(new_n1138), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1139), .B(new_n1140), .C1(new_n740), .C2(new_n872), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1102), .A2(new_n1098), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1142), .A2(KEYINPUT115), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT115), .ZN(new_n1144));
  NOR3_X1   g0944(.A1(new_n1102), .A2(new_n1144), .A3(new_n1098), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1104), .B(new_n1141), .C1(new_n1143), .C2(new_n1145), .ZN(G393));
  INV_X1    g0946(.A(new_n1096), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1091), .A2(new_n1095), .A3(new_n1082), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1147), .A2(new_n750), .A3(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n832), .A2(new_n555), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n862), .B(new_n410), .C1(new_n829), .C2(new_n827), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G322), .C2(new_n857), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1152), .B1(new_n833), .B2(new_n846), .C1(new_n825), .C2(new_n868), .ZN(new_n1153));
  AOI22_X1  g0953(.A1(new_n841), .A2(G311), .B1(G317), .B2(new_n843), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(new_n1154), .B(KEYINPUT52), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n841), .A2(G159), .B1(G150), .B2(new_n843), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1156), .B(KEYINPUT51), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n832), .A2(new_n220), .ZN(new_n1158));
  OAI221_X1 g0958(.A(new_n432), .B1(new_n415), .B2(new_n827), .C1(new_n828), .C2(new_n440), .ZN(new_n1159));
  AOI211_X1 g0959(.A(new_n1158), .B(new_n1159), .C1(G143), .C2(new_n857), .ZN(new_n1160));
  OAI221_X1 g0960(.A(new_n1160), .B1(new_n202), .B2(new_n868), .C1(new_n256), .C2(new_n846), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1153), .A2(new_n1155), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1162), .A2(new_n820), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n244), .A2(new_n813), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1164), .B(new_n821), .C1(new_n205), .C2(new_n210), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1163), .A2(new_n808), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(new_n1068), .B2(new_n819), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1091), .A2(new_n1095), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1167), .B1(new_n1168), .B2(new_n807), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1149), .A2(new_n1169), .ZN(G390));
  AOI21_X1  g0970(.A(new_n984), .B1(new_n1004), .B2(new_n781), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n964), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n963), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  NAND4_X1  g0974(.A1(new_n720), .A2(new_n708), .A3(new_n796), .A4(new_n797), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n880), .A2(new_n394), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(new_n731), .A3(new_n1176), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n973), .B1(new_n1177), .B2(new_n976), .ZN(new_n1178));
  NOR3_X1   g0978(.A1(new_n1178), .A2(new_n991), .A3(new_n964), .ZN(new_n1179));
  OAI211_X1 g0979(.A(new_n993), .B(new_n1171), .C1(new_n1174), .C2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n878), .B1(new_n799), .B2(new_n1176), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1173), .B(new_n1002), .C1(new_n1181), .C2(new_n973), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n787), .A2(G330), .A3(new_n881), .A4(new_n974), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n884), .B1(new_n795), .B2(new_n716), .ZN(new_n1184));
  OAI21_X1  g0984(.A(KEYINPUT105), .B1(new_n1184), .B2(new_n878), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n886), .A2(new_n975), .A3(new_n976), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1185), .A2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n964), .B1(new_n1187), .B2(new_n974), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1182), .B(new_n1183), .C1(new_n1188), .C2(new_n963), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n1180), .A2(new_n807), .A3(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n889), .B1(new_n399), .B2(new_n910), .ZN(new_n1191));
  XOR2_X1   g0991(.A(new_n1191), .B(KEYINPUT119), .Z(new_n1192));
  XNOR2_X1  g0992(.A(KEYINPUT54), .B(G143), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n847), .A2(new_n1194), .B1(G128), .B2(new_n843), .ZN(new_n1195));
  INV_X1    g0995(.A(G132), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1195), .B1(new_n1196), .B2(new_n840), .C1(new_n901), .C2(new_n868), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n410), .B1(new_n861), .B2(G50), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n1198), .A2(KEYINPUT120), .ZN(new_n1199));
  AND2_X1   g0999(.A1(new_n1198), .A2(KEYINPUT120), .ZN(new_n1200));
  NOR2_X1   g1000(.A1(new_n827), .A2(new_n902), .ZN(new_n1201));
  XNOR2_X1  g1001(.A(new_n1201), .B(KEYINPUT53), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n857), .A2(G125), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n866), .A2(G159), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1202), .A2(new_n1203), .A3(new_n1204), .ZN(new_n1205));
  NOR4_X1   g1005(.A1(new_n1197), .A2(new_n1199), .A3(new_n1200), .A4(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT121), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n905), .B1(G294), .B2(new_n857), .ZN(new_n1208));
  INV_X1    g1008(.A(new_n1208), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n1209), .A2(KEYINPUT122), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n864), .A2(new_n410), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1210), .A2(new_n1158), .A3(new_n1211), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1209), .A2(KEYINPUT122), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n841), .A2(G116), .B1(G107), .B2(new_n849), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n847), .A2(G97), .B1(G283), .B2(new_n843), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1212), .A2(new_n1213), .A3(new_n1214), .A4(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1207), .A2(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(KEYINPUT121), .B2(new_n1206), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1192), .B1(new_n909), .B2(new_n1218), .C1(new_n963), .C2(new_n818), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1190), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT118), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n791), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n790), .B1(new_n1175), .B2(new_n731), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n490), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n490), .A2(new_n1171), .ZN(new_n1225));
  AND4_X1   g1025(.A1(new_n1221), .A2(new_n1224), .A3(new_n701), .A4(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1221), .B1(new_n982), .B2(new_n1225), .ZN(new_n1227));
  NOR2_X1   g1027(.A1(new_n1226), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1007), .A2(G330), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n973), .B1(new_n1229), .B2(new_n882), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1230), .A2(new_n1181), .A3(new_n1183), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n787), .A2(G330), .A3(new_n881), .ZN(new_n1232));
  AOI22_X1  g1032(.A1(new_n1232), .A2(new_n973), .B1(new_n993), .B2(new_n1171), .ZN(new_n1233));
  NOR2_X1   g1033(.A1(new_n977), .A2(new_n978), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1231), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1180), .A2(new_n1228), .A3(new_n1189), .A4(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n963), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1179), .B1(new_n1237), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1171), .A2(new_n993), .ZN(new_n1240));
  OAI21_X1  g1040(.A(new_n1189), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n982), .A2(new_n1225), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1242), .A2(KEYINPUT118), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n982), .A2(new_n1221), .A3(new_n1225), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1243), .A2(new_n1235), .A3(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n751), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1220), .B1(new_n1236), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(G378));
  OAI21_X1  g1048(.A(new_n1228), .B1(new_n1241), .B2(new_n1245), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n965), .A2(new_n979), .A3(new_n980), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n984), .B1(new_n1008), .B2(new_n1003), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n273), .A2(new_n728), .ZN(new_n1252));
  OR2_X1    g1052(.A1(new_n311), .A2(new_n1252), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n311), .A2(new_n1252), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  XNOR2_X1  g1055(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1255), .A2(new_n1257), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(new_n1254), .A3(new_n1256), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1260));
  NOR3_X1   g1060(.A1(new_n991), .A2(new_n1000), .A3(new_n985), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT109), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1251), .B(new_n1260), .C1(new_n1261), .C2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1001), .A2(new_n1006), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1260), .B1(new_n1265), .B2(new_n1251), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1250), .B1(new_n1264), .B2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1251), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1260), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1270), .A2(new_n981), .A3(new_n1263), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1249), .A2(KEYINPUT57), .A3(new_n1272), .ZN(new_n1273));
  AOI22_X1  g1073(.A1(new_n1236), .A2(new_n1228), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n750), .C1(KEYINPUT57), .C2(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1264), .A2(new_n1266), .A3(new_n1250), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n981), .B1(new_n1270), .B2(new_n1263), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n807), .B1(new_n1276), .B2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT123), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1269), .A2(new_n817), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n808), .B1(G50), .B2(new_n911), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n432), .A2(G41), .ZN(new_n1282));
  AOI211_X1 g1082(.A(G50), .B(new_n1282), .C1(new_n246), .C2(new_n284), .ZN(new_n1283));
  AOI22_X1  g1083(.A1(new_n866), .A2(G68), .B1(new_n863), .B2(G77), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n857), .A2(G283), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n861), .A2(G58), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1284), .A2(new_n1285), .A3(new_n1282), .A4(new_n1286), .ZN(new_n1287));
  AOI21_X1  g1087(.A(new_n1287), .B1(G107), .B2(new_n841), .ZN(new_n1288));
  AOI22_X1  g1088(.A1(G97), .A2(new_n849), .B1(new_n843), .B2(G116), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1288), .B(new_n1289), .C1(new_n370), .C2(new_n846), .ZN(new_n1290));
  INV_X1    g1090(.A(KEYINPUT58), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1283), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  OAI22_X1  g1092(.A1(new_n832), .A2(new_n902), .B1(new_n827), .B2(new_n1193), .ZN(new_n1293));
  AOI22_X1  g1093(.A1(new_n841), .A2(G128), .B1(G125), .B2(new_n843), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1294), .B1(new_n901), .B2(new_n846), .ZN(new_n1295));
  AOI211_X1 g1095(.A(new_n1293), .B(new_n1295), .C1(G132), .C2(new_n849), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NOR2_X1   g1097(.A1(new_n1297), .A2(KEYINPUT59), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n857), .A2(G124), .ZN(new_n1299));
  AOI211_X1 g1099(.A(G33), .B(G41), .C1(new_n861), .C2(new_n858), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT59), .ZN(new_n1301));
  OAI211_X1 g1101(.A(new_n1299), .B(new_n1300), .C1(new_n1296), .C2(new_n1301), .ZN(new_n1302));
  OAI221_X1 g1102(.A(new_n1292), .B1(new_n1291), .B2(new_n1290), .C1(new_n1298), .C2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1281), .B1(new_n1303), .B2(new_n820), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1280), .A2(new_n1304), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1278), .A2(new_n1279), .A3(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1098), .B1(new_n1267), .B2(new_n1271), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1305), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT123), .B1(new_n1307), .B2(new_n1308), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1275), .A2(new_n1310), .ZN(G375));
  NAND2_X1  g1111(.A1(new_n973), .A2(new_n817), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n808), .B1(G68), .B2(new_n911), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n841), .A2(G283), .B1(G294), .B2(new_n843), .ZN(new_n1314));
  OAI221_X1 g1114(.A(new_n1314), .B1(new_n206), .B2(new_n846), .C1(new_n555), .C2(new_n868), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1029), .A2(new_n410), .ZN(new_n1316));
  OR2_X1    g1116(.A1(new_n1316), .A2(KEYINPUT124), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1316), .A2(KEYINPUT124), .ZN(new_n1318));
  OAI22_X1  g1118(.A1(new_n832), .A2(new_n370), .B1(new_n205), .B2(new_n827), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(G303), .B2(new_n857), .ZN(new_n1320));
  NAND3_X1  g1120(.A1(new_n1317), .A2(new_n1318), .A3(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n843), .A2(G132), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n426), .B1(G159), .B2(new_n863), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n866), .A2(G50), .B1(new_n857), .B2(G128), .ZN(new_n1324));
  NAND4_X1  g1124(.A1(new_n1322), .A2(new_n1286), .A3(new_n1323), .A4(new_n1324), .ZN(new_n1325));
  AOI22_X1  g1125(.A1(new_n847), .A2(G150), .B1(new_n849), .B2(new_n1194), .ZN(new_n1326));
  OAI21_X1  g1126(.A(new_n1326), .B1(new_n901), .B2(new_n840), .ZN(new_n1327));
  OAI22_X1  g1127(.A1(new_n1315), .A2(new_n1321), .B1(new_n1325), .B2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(new_n1313), .B1(new_n1328), .B2(new_n820), .ZN(new_n1329));
  AOI22_X1  g1129(.A1(new_n1235), .A2(new_n807), .B1(new_n1312), .B2(new_n1329), .ZN(new_n1330));
  NAND2_X1  g1130(.A1(new_n1245), .A2(new_n1076), .ZN(new_n1331));
  AOI21_X1  g1131(.A(new_n1235), .B1(new_n1243), .B2(new_n1244), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(new_n1331), .B2(new_n1332), .ZN(G381));
  NOR4_X1   g1133(.A1(G390), .A2(G396), .A3(G393), .A4(G384), .ZN(new_n1334));
  INV_X1    g1134(.A(G381), .ZN(new_n1335));
  AND4_X1   g1135(.A1(new_n1100), .A2(new_n1334), .A3(new_n1247), .A4(new_n1335), .ZN(new_n1336));
  XNOR2_X1  g1136(.A(G375), .B(KEYINPUT125), .ZN(new_n1337));
  AND3_X1   g1137(.A1(new_n1336), .A2(new_n1337), .A3(KEYINPUT126), .ZN(new_n1338));
  AOI21_X1  g1138(.A(KEYINPUT126), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1339));
  OR2_X1    g1139(.A1(new_n1338), .A2(new_n1339), .ZN(G407));
  INV_X1    g1140(.A(G213), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1341), .A2(G343), .ZN(new_n1342));
  INV_X1    g1142(.A(new_n1342), .ZN(new_n1343));
  NOR2_X1   g1143(.A1(G378), .A2(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1341), .B1(new_n1337), .B2(new_n1344), .ZN(new_n1345));
  OAI21_X1  g1145(.A(new_n1345), .B1(new_n1338), .B2(new_n1339), .ZN(G409));
  INV_X1    g1146(.A(KEYINPUT61), .ZN(new_n1347));
  NAND3_X1  g1147(.A1(new_n1275), .A2(new_n1310), .A3(G378), .ZN(new_n1348));
  AND2_X1   g1148(.A1(new_n1274), .A2(new_n1076), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1278), .A2(new_n1305), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1247), .B1(new_n1349), .B2(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1342), .B1(new_n1348), .B2(new_n1351), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1342), .A2(G2897), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1245), .A2(KEYINPUT60), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1354), .B1(new_n1228), .B2(new_n1235), .ZN(new_n1355));
  INV_X1    g1155(.A(new_n1235), .ZN(new_n1356));
  OAI211_X1 g1156(.A(new_n1356), .B(KEYINPUT60), .C1(new_n1226), .C2(new_n1227), .ZN(new_n1357));
  NAND3_X1  g1157(.A1(new_n1355), .A2(new_n750), .A3(new_n1357), .ZN(new_n1358));
  AOI21_X1  g1158(.A(new_n918), .B1(new_n1358), .B2(new_n1330), .ZN(new_n1359));
  AOI21_X1  g1159(.A(new_n1332), .B1(KEYINPUT60), .B2(new_n1245), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1357), .A2(new_n750), .ZN(new_n1361));
  OAI211_X1 g1161(.A(new_n918), .B(new_n1330), .C1(new_n1360), .C2(new_n1361), .ZN(new_n1362));
  INV_X1    g1162(.A(new_n1362), .ZN(new_n1363));
  OAI21_X1  g1163(.A(new_n1353), .B1(new_n1359), .B2(new_n1363), .ZN(new_n1364));
  OAI21_X1  g1164(.A(new_n1330), .B1(new_n1360), .B2(new_n1361), .ZN(new_n1365));
  NAND2_X1  g1165(.A1(new_n1365), .A2(G384), .ZN(new_n1366));
  NAND4_X1  g1166(.A1(new_n1366), .A2(G2897), .A3(new_n1342), .A4(new_n1362), .ZN(new_n1367));
  NAND2_X1  g1167(.A1(new_n1364), .A2(new_n1367), .ZN(new_n1368));
  OAI21_X1  g1168(.A(new_n1347), .B1(new_n1352), .B2(new_n1368), .ZN(new_n1369));
  INV_X1    g1169(.A(new_n1369), .ZN(new_n1370));
  XOR2_X1   g1170(.A(KEYINPUT127), .B(KEYINPUT63), .Z(new_n1371));
  NAND2_X1  g1171(.A1(new_n1348), .A2(new_n1351), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1372), .A2(new_n1343), .ZN(new_n1373));
  NOR2_X1   g1173(.A1(new_n1359), .A2(new_n1363), .ZN(new_n1374));
  OAI21_X1  g1174(.A(new_n1371), .B1(new_n1373), .B2(new_n1374), .ZN(new_n1375));
  NAND2_X1  g1175(.A1(new_n1100), .A2(G390), .ZN(new_n1376));
  INV_X1    g1176(.A(G390), .ZN(new_n1377));
  AOI21_X1  g1177(.A(new_n1073), .B1(new_n1098), .B2(new_n1097), .ZN(new_n1378));
  OAI21_X1  g1178(.A(new_n1377), .B1(new_n1378), .B2(new_n1049), .ZN(new_n1379));
  XNOR2_X1  g1179(.A(G393), .B(new_n876), .ZN(new_n1380));
  AND3_X1   g1180(.A1(new_n1376), .A2(new_n1379), .A3(new_n1380), .ZN(new_n1381));
  AOI21_X1  g1181(.A(new_n1380), .B1(new_n1376), .B2(new_n1379), .ZN(new_n1382));
  NOR2_X1   g1182(.A1(new_n1381), .A2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(new_n1374), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1352), .A2(KEYINPUT63), .A3(new_n1384), .ZN(new_n1385));
  NAND4_X1  g1185(.A1(new_n1370), .A2(new_n1375), .A3(new_n1383), .A4(new_n1385), .ZN(new_n1386));
  INV_X1    g1186(.A(KEYINPUT62), .ZN(new_n1387));
  AND3_X1   g1187(.A1(new_n1352), .A2(new_n1387), .A3(new_n1384), .ZN(new_n1388));
  AOI21_X1  g1188(.A(new_n1387), .B1(new_n1352), .B2(new_n1384), .ZN(new_n1389));
  NOR3_X1   g1189(.A1(new_n1388), .A2(new_n1369), .A3(new_n1389), .ZN(new_n1390));
  OAI21_X1  g1190(.A(new_n1386), .B1(new_n1390), .B2(new_n1383), .ZN(G405));
  NAND2_X1  g1191(.A1(G375), .A2(new_n1247), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1392), .A2(new_n1348), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1393), .A2(new_n1374), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1384), .A2(new_n1392), .A3(new_n1348), .ZN(new_n1395));
  NAND2_X1  g1195(.A1(new_n1394), .A2(new_n1395), .ZN(new_n1396));
  XNOR2_X1  g1196(.A(new_n1396), .B(new_n1383), .ZN(G402));
endmodule


