//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 0 1 1 1 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 0 0 0 1 0 0 1 0 0 1 1 1 1 0 1 0 1 1 1 1 0 1 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:28:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989;
  XNOR2_X1  g000(.A(KEYINPUT22), .B(G137), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND3_X1   g002(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n189));
  XOR2_X1   g003(.A(new_n187), .B(new_n189), .Z(new_n190));
  XNOR2_X1  g004(.A(G125), .B(G140), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT16), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT75), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(G140), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n193), .A2(new_n194), .A3(new_n195), .A4(G125), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(G125), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT75), .B1(new_n197), .B2(KEYINPUT16), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n192), .A2(new_n196), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n192), .A2(G146), .A3(new_n196), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT23), .ZN(new_n204));
  INV_X1    g018(.A(G119), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n204), .B1(new_n205), .B2(G128), .ZN(new_n206));
  INV_X1    g020(.A(G128), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(KEYINPUT23), .A3(G119), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(G128), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n206), .A2(new_n208), .A3(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G110), .ZN(new_n211));
  XOR2_X1   g025(.A(KEYINPUT24), .B(G110), .Z(new_n212));
  XNOR2_X1  g026(.A(G119), .B(G128), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n203), .A2(new_n216), .ZN(new_n217));
  OAI22_X1  g031(.A1(new_n210), .A2(G110), .B1(new_n212), .B2(new_n213), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n191), .A2(new_n200), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n202), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT76), .B1(new_n217), .B2(new_n221), .ZN(new_n222));
  AOI21_X1  g036(.A(new_n215), .B1(new_n201), .B2(new_n202), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT76), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n223), .A2(new_n220), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n190), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G902), .ZN(new_n227));
  INV_X1    g041(.A(new_n190), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n217), .A2(new_n221), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n228), .B1(new_n229), .B2(new_n224), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT25), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT25), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n226), .A2(new_n233), .A3(new_n227), .A4(new_n230), .ZN(new_n234));
  INV_X1    g048(.A(G217), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n235), .B1(G234), .B2(new_n227), .ZN(new_n236));
  XNOR2_X1  g050(.A(new_n236), .B(KEYINPUT74), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n232), .A2(new_n234), .A3(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT77), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n232), .A2(KEYINPUT77), .A3(new_n234), .A4(new_n237), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n236), .A2(G902), .ZN(new_n242));
  XNOR2_X1  g056(.A(new_n242), .B(KEYINPUT78), .ZN(new_n243));
  INV_X1    g057(.A(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n226), .A2(new_n230), .A3(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n240), .A2(new_n241), .A3(new_n245), .ZN(new_n246));
  NOR2_X1   g060(.A1(G472), .A2(G902), .ZN(new_n247));
  INV_X1    g061(.A(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n205), .A2(G116), .ZN(new_n249));
  INV_X1    g063(.A(G116), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n250), .A2(G119), .ZN(new_n251));
  INV_X1    g065(.A(G113), .ZN(new_n252));
  AND2_X1   g066(.A1(new_n252), .A2(KEYINPUT2), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(KEYINPUT2), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n249), .B(new_n251), .C1(new_n253), .C2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n249), .A2(new_n251), .ZN(new_n256));
  XNOR2_X1  g070(.A(KEYINPUT2), .B(G113), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT69), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n255), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n256), .A2(new_n257), .A3(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n200), .A2(G143), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT65), .ZN(new_n265));
  INV_X1    g079(.A(G143), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n265), .B1(new_n266), .B2(G146), .ZN(new_n267));
  NOR3_X1   g081(.A1(new_n200), .A2(KEYINPUT65), .A3(G143), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n264), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT0), .A2(G128), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n266), .A2(G146), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT64), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n272), .B1(new_n200), .B2(G143), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n266), .A2(KEYINPUT64), .A3(G146), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  XNOR2_X1  g089(.A(KEYINPUT0), .B(G128), .ZN(new_n276));
  OAI22_X1  g090(.A1(new_n269), .A2(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  AND2_X1   g091(.A1(KEYINPUT68), .A2(G137), .ZN(new_n278));
  NOR2_X1   g092(.A1(KEYINPUT68), .A2(G137), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT11), .ZN(new_n281));
  INV_X1    g095(.A(G134), .ZN(new_n282));
  NOR2_X1   g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n280), .A2(new_n283), .B1(new_n282), .B2(G137), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n285));
  XNOR2_X1  g099(.A(KEYINPUT66), .B(KEYINPUT11), .ZN(new_n286));
  INV_X1    g100(.A(G137), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n287), .A2(G134), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n281), .A2(KEYINPUT66), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT66), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n291), .A2(KEYINPUT11), .ZN(new_n292));
  AND4_X1   g106(.A1(new_n285), .A2(new_n288), .A3(new_n290), .A4(new_n292), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n284), .B1(new_n289), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n294), .A2(G131), .ZN(new_n295));
  INV_X1    g109(.A(G131), .ZN(new_n296));
  OAI211_X1 g110(.A(new_n284), .B(new_n296), .C1(new_n289), .C2(new_n293), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n277), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT1), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n207), .B1(new_n264), .B2(KEYINPUT1), .ZN(new_n301));
  OAI22_X1  g115(.A1(new_n269), .A2(new_n300), .B1(new_n275), .B2(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n288), .B1(new_n280), .B2(G134), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G131), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n297), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  NOR3_X1   g119(.A1(new_n298), .A2(new_n305), .A3(KEYINPUT30), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT30), .ZN(new_n307));
  INV_X1    g121(.A(new_n277), .ZN(new_n308));
  INV_X1    g122(.A(new_n297), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n288), .A2(new_n290), .A3(new_n292), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT67), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n286), .A2(new_n285), .A3(new_n288), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g127(.A(new_n296), .B1(new_n313), .B2(new_n284), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n308), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n297), .A2(new_n302), .A3(new_n304), .ZN(new_n316));
  AOI21_X1  g130(.A(new_n307), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n263), .B1(new_n306), .B2(new_n317), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n260), .A2(KEYINPUT70), .A3(new_n261), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT70), .B1(new_n260), .B2(new_n261), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n315), .A2(new_n321), .A3(new_n316), .ZN(new_n322));
  XOR2_X1   g136(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n323));
  NOR2_X1   g137(.A1(G237), .A2(G953), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G210), .ZN(new_n325));
  XNOR2_X1  g139(.A(new_n323), .B(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(KEYINPUT26), .B(G101), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n326), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n318), .A2(new_n322), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT31), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(new_n322), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT30), .B1(new_n298), .B2(new_n305), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n315), .A2(new_n307), .A3(new_n316), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n333), .B1(new_n336), .B2(new_n263), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(KEYINPUT31), .A3(new_n329), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n262), .B1(new_n315), .B2(new_n316), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT28), .B1(new_n333), .B2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT28), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n322), .A2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT72), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n322), .A2(KEYINPUT72), .A3(new_n342), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n341), .A2(new_n345), .A3(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n328), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n248), .B1(new_n339), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT73), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n337), .B2(new_n329), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT29), .ZN(new_n352));
  NAND4_X1  g166(.A1(new_n341), .A2(new_n345), .A3(new_n346), .A4(new_n329), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n262), .B1(new_n334), .B2(new_n335), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT73), .B(new_n328), .C1(new_n354), .C2(new_n333), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n351), .A2(new_n352), .A3(new_n353), .A4(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n346), .ZN(new_n357));
  OAI22_X1  g171(.A1(new_n298), .A2(new_n305), .B1(new_n319), .B2(new_n320), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n342), .B1(new_n358), .B2(new_n322), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT72), .B1(new_n322), .B2(new_n342), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n357), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n328), .A2(new_n352), .ZN(new_n362));
  AOI21_X1  g176(.A(G902), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n356), .A2(new_n363), .ZN(new_n364));
  AOI22_X1  g178(.A1(KEYINPUT32), .A2(new_n349), .B1(new_n364), .B2(G472), .ZN(new_n365));
  INV_X1    g179(.A(KEYINPUT32), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n332), .A2(new_n338), .B1(new_n347), .B2(new_n328), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n366), .B1(new_n367), .B2(new_n248), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n246), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(G221), .ZN(new_n370));
  XNOR2_X1  g184(.A(KEYINPUT9), .B(G234), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n370), .B1(new_n372), .B2(new_n227), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n374));
  INV_X1    g188(.A(new_n301), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n269), .A2(new_n375), .A3(KEYINPUT79), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT79), .ZN(new_n377));
  OAI21_X1  g191(.A(KEYINPUT65), .B1(new_n200), .B2(G143), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n265), .A2(new_n266), .A3(G146), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n271), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  OAI21_X1  g194(.A(new_n377), .B1(new_n380), .B2(new_n301), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(new_n299), .A3(G128), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n376), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G104), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(G107), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n384), .A2(G107), .ZN(new_n387));
  OAI21_X1  g201(.A(G101), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g202(.A(KEYINPUT3), .B1(new_n384), .B2(G107), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n390), .A2(new_n391), .A3(G104), .ZN(new_n392));
  INV_X1    g206(.A(G101), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n389), .A2(new_n392), .A3(new_n393), .A4(new_n385), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n383), .A2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT80), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n398), .B1(new_n302), .B2(new_n396), .ZN(new_n399));
  OR2_X1    g213(.A1(new_n275), .A2(new_n301), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n400), .A2(KEYINPUT80), .A3(new_n382), .A4(new_n395), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n397), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n295), .A2(new_n297), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT12), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT81), .ZN(new_n405));
  AOI21_X1  g219(.A(KEYINPUT12), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  NOR2_X1   g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n402), .A2(new_n403), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT81), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT12), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n408), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n302), .A2(new_n396), .A3(KEYINPUT10), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n389), .A2(new_n392), .A3(new_n385), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT4), .A3(new_n394), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n413), .A2(new_n416), .A3(G101), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n412), .B1(new_n418), .B2(new_n277), .ZN(new_n419));
  AOI21_X1  g233(.A(KEYINPUT10), .B1(new_n383), .B2(new_n396), .ZN(new_n420));
  NOR3_X1   g234(.A1(new_n419), .A2(new_n420), .A3(new_n403), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n411), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n374), .B1(new_n407), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G110), .B(G140), .ZN(new_n425));
  INV_X1    g239(.A(G227), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(G953), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n425), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n408), .A2(new_n410), .ZN(new_n429));
  NAND3_X1  g243(.A1(new_n429), .A2(KEYINPUT81), .A3(new_n404), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT82), .A3(new_n411), .A4(new_n422), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n424), .A2(new_n428), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n428), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n403), .B1(new_n419), .B2(new_n420), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n422), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n432), .A2(G469), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G469), .ZN(new_n437));
  NOR2_X1   g251(.A1(new_n437), .A2(new_n227), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n433), .B1(new_n422), .B2(new_n434), .ZN(new_n442));
  NAND4_X1  g256(.A1(new_n430), .A2(new_n433), .A3(new_n411), .A4(new_n422), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT83), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n423), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n446), .A2(KEYINPUT83), .A3(new_n433), .A4(new_n430), .ZN(new_n447));
  AOI21_X1  g261(.A(G902), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n437), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n373), .B1(new_n441), .B2(new_n449), .ZN(new_n450));
  INV_X1    g264(.A(G122), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G116), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n250), .A2(G122), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT92), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT92), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n452), .A2(new_n453), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n458), .A2(new_n391), .ZN(new_n459));
  AOI21_X1  g273(.A(G107), .B1(new_n455), .B2(new_n457), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT93), .ZN(new_n461));
  OAI22_X1  g275(.A1(new_n461), .A2(KEYINPUT13), .B1(new_n266), .B2(G128), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n461), .A2(KEYINPUT13), .ZN(new_n463));
  OAI21_X1  g277(.A(G134), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(G128), .B(G143), .Z(new_n465));
  AND2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(new_n464), .A2(new_n465), .ZN(new_n467));
  OAI22_X1  g281(.A1(new_n459), .A2(new_n460), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n460), .ZN(new_n469));
  XNOR2_X1  g283(.A(new_n465), .B(G134), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n250), .A2(KEYINPUT14), .A3(G122), .ZN(new_n471));
  OAI211_X1 g285(.A(G107), .B(new_n471), .C1(new_n454), .C2(KEYINPUT14), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n469), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n371), .A2(new_n235), .A3(G953), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n468), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n468), .B2(new_n473), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n227), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT15), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(G478), .ZN(new_n479));
  INV_X1    g293(.A(G478), .ZN(new_n480));
  OAI221_X1 g294(.A(new_n227), .B1(KEYINPUT15), .B2(new_n480), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n479), .A2(new_n481), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n482), .B(KEYINPUT94), .Z(new_n483));
  NAND3_X1  g297(.A1(new_n324), .A2(G143), .A3(G214), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(G143), .B1(new_n324), .B2(G214), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(KEYINPUT18), .A2(G131), .ZN(new_n488));
  OR2_X1    g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(new_n488), .ZN(new_n490));
  INV_X1    g304(.A(G125), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G140), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n197), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(G146), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n219), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n489), .A2(new_n490), .A3(new_n495), .ZN(new_n496));
  OAI21_X1  g310(.A(G131), .B1(new_n485), .B2(new_n486), .ZN(new_n497));
  INV_X1    g311(.A(new_n486), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n498), .A2(new_n296), .A3(new_n484), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g314(.A1(new_n191), .A2(KEYINPUT19), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n191), .A2(KEYINPUT19), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n200), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AND2_X1   g317(.A1(new_n503), .A2(new_n202), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT89), .ZN(new_n505));
  OAI21_X1  g319(.A(new_n500), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n503), .A2(new_n505), .A3(new_n202), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n496), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  XNOR2_X1  g322(.A(G113), .B(G122), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n509), .B(new_n384), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT17), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n497), .A2(new_n499), .A3(new_n512), .ZN(new_n513));
  OAI211_X1 g327(.A(KEYINPUT17), .B(G131), .C1(new_n485), .C2(new_n486), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n513), .A2(new_n201), .A3(new_n202), .A4(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n515), .A2(new_n496), .A3(new_n510), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(KEYINPUT90), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT90), .ZN(new_n518));
  NAND4_X1  g332(.A1(new_n515), .A2(new_n496), .A3(new_n518), .A4(new_n510), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n508), .A2(new_n511), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(KEYINPUT20), .B1(new_n520), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n517), .A2(new_n519), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n505), .B1(new_n503), .B2(new_n202), .ZN(new_n525));
  INV_X1    g339(.A(new_n500), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n507), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  INV_X1    g341(.A(new_n496), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n511), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT20), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n530), .A2(new_n531), .A3(new_n521), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n523), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g347(.A1(new_n515), .A2(new_n496), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n524), .B1(new_n510), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(new_n227), .ZN(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT91), .B(G475), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND2_X1   g352(.A1(new_n533), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(G234), .A2(G237), .ZN(new_n540));
  AND3_X1   g354(.A1(new_n540), .A2(G952), .A3(new_n188), .ZN(new_n541));
  XNOR2_X1  g355(.A(KEYINPUT21), .B(G898), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT95), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  AND3_X1   g358(.A1(new_n540), .A2(G902), .A3(G953), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n483), .A2(new_n539), .A3(new_n547), .ZN(new_n548));
  OAI21_X1  g362(.A(G214), .B1(G237), .B2(G902), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n250), .A2(G119), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT5), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n552), .B(G113), .C1(new_n256), .C2(new_n551), .ZN(new_n553));
  AND2_X1   g367(.A1(new_n553), .A2(new_n255), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n554), .A2(KEYINPUT86), .A3(new_n396), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT86), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n255), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n395), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n555), .B(new_n558), .C1(new_n396), .C2(new_n554), .ZN(new_n559));
  XNOR2_X1  g373(.A(G110), .B(G122), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT85), .B(KEYINPUT8), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT87), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n559), .A2(KEYINPUT87), .A3(new_n562), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n277), .A2(G125), .ZN(new_n568));
  OAI21_X1  g382(.A(new_n568), .B1(G125), .B2(new_n302), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n188), .A2(G224), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT7), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n571), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n568), .B(new_n573), .C1(G125), .C2(new_n302), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n415), .A2(new_n261), .A3(new_n260), .A4(new_n417), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n554), .A2(new_n396), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT84), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .A4(new_n560), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n577), .A3(new_n560), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(KEYINPUT84), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n575), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g396(.A(G902), .B1(new_n567), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n560), .B1(new_n576), .B2(new_n577), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n584), .A2(KEYINPUT6), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT6), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n586), .B1(new_n581), .B2(new_n579), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n585), .B1(new_n587), .B2(new_n584), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n569), .B(new_n570), .Z(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(G210), .B1(G237), .B2(G902), .ZN(new_n591));
  AND3_X1   g405(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n583), .B2(new_n590), .ZN(new_n593));
  OAI21_X1  g407(.A(new_n549), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n594), .A2(KEYINPUT88), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n583), .A2(new_n590), .ZN(new_n596));
  INV_X1    g410(.A(new_n591), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n583), .A2(new_n590), .A3(new_n591), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT88), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n600), .A2(new_n601), .A3(new_n549), .ZN(new_n602));
  AOI21_X1  g416(.A(new_n548), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n369), .A2(new_n450), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G101), .ZN(G3));
  OAI21_X1  g419(.A(G472), .B1(new_n367), .B2(G902), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n367), .B2(new_n248), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n607), .A2(new_n246), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n450), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n549), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n610), .B1(new_n592), .B2(KEYINPUT96), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n598), .A2(new_n612), .A3(new_n599), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n611), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(KEYINPUT97), .B(KEYINPUT33), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n475), .B2(new_n476), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n480), .A2(G902), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT99), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n468), .A2(new_n473), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n618), .B1(new_n619), .B2(KEYINPUT98), .ZN(new_n620));
  INV_X1    g434(.A(new_n474), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT98), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n622), .B1(new_n621), .B2(KEYINPUT99), .ZN(new_n623));
  AOI22_X1  g437(.A1(new_n620), .A2(new_n621), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT33), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n616), .B(new_n617), .C1(new_n624), .C2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n477), .A2(new_n480), .ZN(new_n627));
  AOI22_X1  g441(.A1(new_n533), .A2(new_n538), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n629), .A2(new_n546), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n609), .A2(new_n614), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  AND2_X1   g447(.A1(new_n536), .A2(new_n537), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n483), .A2(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT100), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n531), .B1(new_n530), .B2(new_n521), .ZN(new_n637));
  AOI211_X1 g451(.A(KEYINPUT20), .B(new_n522), .C1(new_n524), .C2(new_n529), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n523), .A2(new_n532), .A3(KEYINPUT100), .ZN(new_n640));
  AND2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g455(.A1(new_n635), .A2(new_n547), .A3(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n609), .A2(new_n614), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G107), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n644), .B(new_n645), .ZN(G9));
  NOR2_X1   g460(.A1(new_n228), .A2(KEYINPUT36), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n229), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n244), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n240), .A2(new_n241), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n607), .A2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n450), .A2(new_n603), .A3(new_n652), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT37), .B(G110), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(new_n373), .ZN(new_n656));
  AOI211_X1 g470(.A(G469), .B(G902), .C1(new_n445), .C2(new_n447), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n656), .B(new_n650), .C1(new_n657), .C2(new_n440), .ZN(new_n658));
  INV_X1    g472(.A(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n541), .B1(new_n545), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  AND3_X1   g476(.A1(new_n635), .A2(new_n641), .A3(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n611), .A2(new_n613), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n664), .B1(new_n365), .B2(new_n368), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n659), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G128), .ZN(G30));
  XOR2_X1   g481(.A(new_n661), .B(KEYINPUT39), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n450), .A2(new_n668), .ZN(new_n669));
  OR2_X1    g483(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n670));
  XOR2_X1   g484(.A(KEYINPUT102), .B(KEYINPUT38), .Z(new_n671));
  XNOR2_X1  g485(.A(new_n600), .B(new_n671), .ZN(new_n672));
  NOR4_X1   g486(.A1(new_n650), .A2(new_n483), .A3(new_n539), .A4(new_n610), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n349), .A2(KEYINPUT32), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n337), .A2(new_n328), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n358), .A2(new_n322), .A3(new_n328), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n227), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n675), .B2(new_n677), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n674), .A2(new_n368), .A3(new_n678), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n672), .A2(new_n673), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n669), .A2(KEYINPUT40), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n670), .A2(new_n680), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  NOR2_X1   g497(.A1(new_n629), .A2(new_n661), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n659), .A2(new_n665), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G146), .ZN(G48));
  NAND2_X1  g500(.A1(new_n443), .A2(new_n444), .ZN(new_n687));
  INV_X1    g501(.A(new_n442), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n687), .A2(new_n447), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n437), .B1(new_n689), .B2(new_n227), .ZN(new_n690));
  NOR3_X1   g504(.A1(new_n657), .A2(new_n690), .A3(new_n373), .ZN(new_n691));
  NAND4_X1  g505(.A1(new_n369), .A2(new_n614), .A3(new_n691), .A4(new_n630), .ZN(new_n692));
  XNOR2_X1  g506(.A(KEYINPUT41), .B(G113), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT103), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n692), .B(new_n694), .ZN(G15));
  NAND4_X1  g509(.A1(new_n369), .A2(new_n642), .A3(new_n691), .A4(new_n614), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G116), .ZN(G18));
  NOR2_X1   g511(.A1(new_n548), .A2(new_n651), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n364), .A2(G472), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n674), .A2(new_n699), .A3(new_n368), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n691), .A2(new_n698), .A3(new_n700), .A4(new_n614), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G119), .ZN(G21));
  NOR3_X1   g516(.A1(new_n664), .A2(new_n539), .A3(new_n483), .ZN(new_n703));
  INV_X1    g517(.A(new_n246), .ZN(new_n704));
  AOI21_X1  g518(.A(KEYINPUT31), .B1(new_n337), .B2(new_n329), .ZN(new_n705));
  NOR4_X1   g519(.A1(new_n354), .A2(new_n333), .A3(new_n331), .A4(new_n328), .ZN(new_n706));
  OAI22_X1  g520(.A1(new_n705), .A2(new_n706), .B1(new_n361), .B2(new_n329), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(new_n247), .ZN(new_n708));
  AND4_X1   g522(.A1(new_n704), .A2(new_n606), .A3(new_n547), .A4(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n703), .A2(new_n709), .A3(new_n691), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G122), .ZN(G24));
  INV_X1    g525(.A(new_n684), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n606), .A2(new_n650), .A3(new_n708), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT104), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n606), .A2(new_n650), .A3(new_n715), .A4(new_n708), .ZN(new_n716));
  AOI21_X1  g530(.A(new_n712), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  NOR4_X1   g531(.A1(new_n664), .A2(new_n657), .A3(new_n690), .A4(new_n373), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(G125), .ZN(G27));
  INV_X1    g534(.A(KEYINPUT108), .ZN(new_n721));
  OAI21_X1  g535(.A(new_n721), .B1(new_n349), .B2(KEYINPUT32), .ZN(new_n722));
  OAI211_X1 g536(.A(KEYINPUT108), .B(new_n366), .C1(new_n367), .C2(new_n248), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n722), .A2(new_n674), .A3(new_n699), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n724), .A2(new_n704), .A3(new_n684), .ZN(new_n725));
  INV_X1    g539(.A(KEYINPUT106), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n432), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n424), .A2(new_n431), .A3(KEYINPUT106), .A4(new_n428), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n435), .B(KEYINPUT107), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n727), .A2(G469), .A3(new_n728), .A4(new_n729), .ZN(new_n730));
  XOR2_X1   g544(.A(new_n438), .B(KEYINPUT105), .Z(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n730), .A2(new_n449), .A3(new_n732), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n592), .A2(new_n593), .A3(new_n610), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n656), .A3(new_n734), .ZN(new_n735));
  OAI21_X1  g549(.A(KEYINPUT42), .B1(new_n725), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n598), .A2(new_n549), .A3(new_n599), .ZN(new_n737));
  AOI21_X1  g551(.A(new_n731), .B1(new_n448), .B2(new_n437), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n373), .B(new_n737), .C1(new_n738), .C2(new_n730), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n712), .A2(KEYINPUT42), .ZN(new_n740));
  NAND3_X1  g554(.A1(new_n739), .A2(new_n369), .A3(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n736), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT109), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT109), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n736), .A2(new_n744), .A3(new_n741), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND3_X1  g561(.A1(new_n739), .A2(new_n369), .A3(new_n663), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G134), .ZN(G36));
  AOI21_X1  g563(.A(KEYINPUT43), .B1(new_n539), .B2(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n626), .A2(new_n627), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n539), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n750), .B(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n753), .A2(KEYINPUT44), .A3(new_n607), .A4(new_n650), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(KEYINPUT111), .ZN(new_n755));
  AND3_X1   g569(.A1(new_n753), .A2(new_n607), .A3(new_n650), .ZN(new_n756));
  OAI211_X1 g570(.A(new_n755), .B(new_n734), .C1(KEYINPUT44), .C2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(KEYINPUT45), .B1(new_n432), .B2(new_n435), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n758), .A2(new_n437), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n727), .A2(KEYINPUT45), .A3(new_n728), .A4(new_n729), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n731), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n657), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n373), .B1(new_n764), .B2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n668), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n757), .A2(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(new_n287), .ZN(G39));
  XNOR2_X1  g583(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n770));
  OR2_X1    g584(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT47), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n766), .B1(KEYINPUT112), .B2(new_n772), .ZN(new_n773));
  NOR4_X1   g587(.A1(new_n712), .A2(new_n700), .A3(new_n704), .A4(new_n737), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n771), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT113), .ZN(new_n776));
  XNOR2_X1  g590(.A(new_n776), .B(G140), .ZN(G42));
  NOR2_X1   g591(.A1(new_n657), .A2(new_n690), .ZN(new_n778));
  XOR2_X1   g592(.A(new_n778), .B(KEYINPUT114), .Z(new_n779));
  XNOR2_X1  g593(.A(new_n779), .B(KEYINPUT49), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n679), .A2(new_n246), .ZN(new_n781));
  OR4_X1    g595(.A1(new_n373), .A2(new_n672), .A3(new_n610), .A4(new_n752), .ZN(new_n782));
  OR3_X1    g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT121), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n771), .A2(new_n773), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n779), .A2(new_n656), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT119), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n606), .A2(new_n708), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n753), .A2(new_n704), .A3(new_n541), .A4(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n791), .A2(new_n737), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n789), .A2(new_n792), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n672), .A2(new_n549), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(new_n691), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(KEYINPUT50), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT50), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n798), .B1(new_n791), .B2(new_n795), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n714), .A2(new_n716), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n753), .A2(new_n541), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n691), .A2(new_n734), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n541), .ZN(new_n805));
  NOR3_X1   g619(.A1(new_n803), .A2(new_n781), .A3(new_n805), .ZN(new_n806));
  AOI211_X1 g620(.A(new_n751), .B(new_n634), .C1(new_n523), .C2(new_n532), .ZN(new_n807));
  AOI22_X1  g621(.A1(new_n801), .A2(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n800), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(KEYINPUT51), .B1(new_n793), .B2(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n786), .B1(new_n771), .B2(new_n773), .ZN(new_n811));
  INV_X1    g625(.A(new_n792), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n809), .B(KEYINPUT51), .C1(new_n811), .C2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n718), .ZN(new_n814));
  OAI211_X1 g628(.A(G952), .B(new_n188), .C1(new_n791), .C2(new_n814), .ZN(new_n815));
  NOR4_X1   g629(.A1(new_n803), .A2(new_n781), .A3(new_n805), .A4(new_n629), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT48), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n724), .A2(new_n704), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n804), .A2(new_n818), .A3(new_n819), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n818), .B1(new_n804), .B2(new_n819), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n817), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT120), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI211_X1 g638(.A(new_n817), .B(KEYINPUT120), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n813), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g641(.A(new_n784), .B1(new_n810), .B2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT51), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n812), .B1(new_n785), .B2(new_n788), .ZN(new_n830));
  INV_X1    g644(.A(new_n809), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n829), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT121), .A3(new_n826), .A4(new_n813), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n828), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n717), .A2(new_n739), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n482), .B1(new_n536), .B2(new_n537), .ZN(new_n836));
  AND4_X1   g650(.A1(new_n640), .A2(new_n639), .A3(new_n662), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n837), .A2(new_n734), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n838), .B1(new_n368), .B2(new_n365), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n659), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n748), .A2(new_n835), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AOI22_X1  g657(.A1(new_n717), .A2(new_n739), .B1(new_n659), .B2(new_n839), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .A3(new_n748), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n700), .A2(new_n614), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(new_n658), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n663), .A2(new_n848), .B1(new_n717), .B2(new_n718), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n373), .B1(new_n738), .B2(new_n730), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n650), .A2(new_n661), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n703), .A2(new_n850), .A3(new_n679), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n849), .A2(KEYINPUT52), .A3(new_n685), .A4(new_n852), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n719), .A2(new_n666), .A3(new_n685), .A4(new_n852), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT52), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n692), .A2(new_n696), .A3(new_n604), .A4(new_n710), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n595), .A2(new_n602), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n628), .B1(new_n539), .B2(new_n482), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n860), .A2(new_n546), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n450), .A2(new_n608), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n862), .A2(new_n653), .A3(new_n701), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n858), .A2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n746), .A2(new_n846), .A3(new_n857), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT53), .ZN(new_n866));
  OAI21_X1  g680(.A(KEYINPUT117), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n746), .A2(new_n846), .A3(new_n864), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n853), .A2(new_n856), .A3(KEYINPUT116), .ZN(new_n869));
  OR3_X1    g683(.A1(new_n854), .A2(KEYINPUT116), .A3(new_n855), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n866), .B1(new_n868), .B2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n864), .A2(new_n743), .A3(new_n745), .ZN(new_n873));
  AND4_X1   g687(.A1(KEYINPUT115), .A2(new_n748), .A3(new_n835), .A4(new_n840), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT115), .B1(new_n844), .B2(new_n748), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n873), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT117), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(KEYINPUT53), .A4(new_n857), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n867), .A2(new_n872), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT54), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n865), .A2(new_n866), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT54), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n742), .A2(new_n866), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n884), .A2(new_n864), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n885), .A2(new_n869), .A3(new_n846), .A4(new_n870), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n882), .A2(new_n883), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n881), .A2(KEYINPUT118), .A3(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT118), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n880), .A2(new_n889), .A3(KEYINPUT54), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n834), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(G952), .A2(G953), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n783), .B1(new_n891), .B2(new_n892), .ZN(G75));
  NAND2_X1  g707(.A1(new_n882), .A2(new_n886), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(G210), .A3(G902), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT56), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n588), .B(new_n589), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n898), .B(KEYINPUT55), .Z(new_n899));
  NAND4_X1  g713(.A1(new_n895), .A2(new_n896), .A3(new_n897), .A4(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n188), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n895), .A2(new_n897), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n895), .A2(KEYINPUT122), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n905), .A2(new_n899), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(G51));
  AND4_X1   g721(.A1(G902), .A2(new_n894), .A3(new_n760), .A4(new_n759), .ZN(new_n908));
  INV_X1    g722(.A(new_n689), .ZN(new_n909));
  AOI21_X1  g723(.A(KEYINPUT53), .B1(new_n877), .B2(new_n857), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n846), .A2(new_n864), .A3(new_n884), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n871), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g726(.A(KEYINPUT54), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n887), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n731), .B(KEYINPUT57), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n909), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n908), .B1(new_n916), .B2(KEYINPUT123), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT123), .ZN(new_n918));
  INV_X1    g732(.A(new_n915), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n919), .B1(new_n913), .B2(new_n887), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n918), .B1(new_n920), .B2(new_n909), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n901), .B1(new_n917), .B2(new_n921), .ZN(G54));
  NAND4_X1  g736(.A1(new_n894), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n923));
  AND2_X1   g737(.A1(new_n923), .A2(new_n520), .ZN(new_n924));
  NOR2_X1   g738(.A1(new_n923), .A2(new_n520), .ZN(new_n925));
  NOR3_X1   g739(.A1(new_n924), .A2(new_n925), .A3(new_n901), .ZN(G60));
  INV_X1    g740(.A(new_n914), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n616), .B1(new_n624), .B2(new_n625), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT124), .Z(new_n929));
  NAND2_X1  g743(.A1(G478), .A2(G902), .ZN(new_n930));
  XOR2_X1   g744(.A(new_n930), .B(KEYINPUT59), .Z(new_n931));
  OR2_X1    g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n902), .B1(new_n927), .B2(new_n932), .ZN(new_n933));
  INV_X1    g747(.A(new_n931), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n888), .A2(new_n890), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n933), .B1(new_n935), .B2(new_n929), .ZN(G63));
  NAND2_X1  g750(.A1(G217), .A2(G902), .ZN(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT60), .Z(new_n938));
  NAND3_X1  g752(.A1(new_n894), .A2(new_n648), .A3(new_n938), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n894), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n226), .A2(new_n230), .ZN(new_n941));
  XOR2_X1   g755(.A(new_n941), .B(KEYINPUT125), .Z(new_n942));
  OAI211_X1 g756(.A(new_n902), .B(new_n939), .C1(new_n940), .C2(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT61), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G66));
  INV_X1    g759(.A(G224), .ZN(new_n946));
  OAI21_X1  g760(.A(G953), .B1(new_n544), .B2(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n947), .B1(new_n864), .B2(G953), .ZN(new_n948));
  INV_X1    g762(.A(new_n588), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(G898), .B2(new_n188), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n948), .B(new_n950), .ZN(G69));
  OAI21_X1  g765(.A(G953), .B1(new_n426), .B2(new_n660), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT126), .Z(new_n953));
  NOR2_X1   g767(.A1(new_n501), .A2(new_n502), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n336), .B(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  INV_X1    g770(.A(new_n369), .ZN(new_n957));
  NOR4_X1   g771(.A1(new_n669), .A2(new_n957), .A3(new_n737), .A4(new_n860), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n768), .A2(new_n958), .ZN(new_n959));
  AND3_X1   g773(.A1(new_n719), .A2(new_n666), .A3(new_n685), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n682), .A2(new_n960), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT62), .Z(new_n962));
  NAND3_X1  g776(.A1(new_n776), .A2(new_n959), .A3(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n956), .B1(new_n963), .B2(new_n188), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n819), .A2(new_n703), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n767), .B1(new_n757), .B2(new_n966), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n746), .A2(new_n748), .A3(new_n960), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g783(.A1(new_n776), .A2(new_n969), .A3(new_n188), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n955), .B1(G900), .B2(G953), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n953), .B1(new_n965), .B2(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(new_n972), .ZN(new_n974));
  INV_X1    g788(.A(new_n953), .ZN(new_n975));
  NOR3_X1   g789(.A1(new_n974), .A2(new_n964), .A3(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n973), .A2(new_n976), .ZN(G72));
  NAND3_X1  g791(.A1(new_n776), .A2(new_n969), .A3(new_n864), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT127), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n978), .A2(new_n981), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n354), .A2(new_n333), .A3(new_n329), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n901), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n864), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n981), .B1(new_n963), .B2(new_n985), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n986), .A2(new_n675), .ZN(new_n987));
  NAND3_X1  g801(.A1(new_n351), .A2(new_n330), .A3(new_n355), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n880), .A2(new_n980), .A3(new_n988), .ZN(new_n989));
  AND3_X1   g803(.A1(new_n984), .A2(new_n987), .A3(new_n989), .ZN(G57));
endmodule


