//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 0 0 0 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:14:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n707, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n810, new_n811, new_n812, new_n813,
    new_n815, new_n816, new_n817, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n954, new_n955, new_n956;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT25), .ZN(new_n203));
  INV_X1    g002(.A(G183gat), .ZN(new_n204));
  INV_X1    g003(.A(G190gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(G183gat), .A2(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT24), .A3(new_n207), .ZN(new_n208));
  OAI21_X1  g007(.A(new_n208), .B1(KEYINPUT24), .B2(new_n207), .ZN(new_n209));
  NOR2_X1   g008(.A1(G169gat), .A2(G176gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT23), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT23), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n211), .A2(new_n212), .A3(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n203), .B1(new_n209), .B2(new_n215), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n203), .ZN(new_n217));
  NOR2_X1   g016(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n218));
  OR2_X1    g017(.A1(new_n218), .A2(new_n207), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n207), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n219), .A2(new_n206), .A3(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n217), .A2(new_n221), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT65), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(KEYINPUT27), .B(G183gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n205), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT66), .B(KEYINPUT28), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n210), .B(KEYINPUT26), .ZN(new_n230));
  AOI22_X1  g029(.A1(new_n230), .A2(new_n212), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n225), .A2(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(G127gat), .B(G134gat), .Z(new_n234));
  INV_X1    g033(.A(G113gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n235), .A2(KEYINPUT68), .A3(G120gat), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT68), .ZN(new_n237));
  INV_X1    g036(.A(G120gat), .ZN(new_n238));
  AOI21_X1  g037(.A(new_n237), .B1(G113gat), .B2(new_n238), .ZN(new_n239));
  NOR2_X1   g038(.A1(new_n238), .A2(G113gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n236), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AOI211_X1 g040(.A(KEYINPUT1), .B(new_n234), .C1(new_n241), .C2(KEYINPUT69), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n242), .B1(KEYINPUT69), .B2(new_n241), .ZN(new_n243));
  XNOR2_X1  g042(.A(G113gat), .B(G120gat), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n234), .B1(KEYINPUT1), .B2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n248), .ZN(new_n249));
  AND2_X1   g048(.A1(new_n243), .A2(new_n247), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n225), .A2(new_n250), .A3(new_n232), .ZN(new_n251));
  AOI21_X1  g050(.A(new_n202), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT32), .ZN(new_n253));
  OR3_X1    g052(.A1(new_n252), .A2(new_n253), .A3(KEYINPUT34), .ZN(new_n254));
  OAI21_X1  g053(.A(KEYINPUT34), .B1(new_n252), .B2(new_n253), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n249), .A2(new_n202), .A3(new_n251), .ZN(new_n257));
  XNOR2_X1  g056(.A(G15gat), .B(G99gat), .ZN(new_n258));
  INV_X1    g057(.A(G43gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(KEYINPUT70), .B(G71gat), .ZN(new_n261));
  XOR2_X1   g060(.A(new_n260), .B(new_n261), .Z(new_n262));
  OAI211_X1 g061(.A(new_n257), .B(new_n262), .C1(new_n252), .C2(KEYINPUT33), .ZN(new_n263));
  AND2_X1   g062(.A1(new_n249), .A2(new_n251), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT33), .ZN(new_n265));
  INV_X1    g064(.A(new_n262), .ZN(new_n266));
  OAI211_X1 g065(.A(new_n264), .B(new_n202), .C1(new_n265), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n256), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g068(.A1(new_n254), .A2(new_n263), .A3(new_n267), .A4(new_n255), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n269), .A2(KEYINPUT36), .A3(new_n270), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT36), .B1(new_n269), .B2(new_n270), .ZN(new_n272));
  NOR2_X1   g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(G211gat), .B(G218gat), .ZN(new_n274));
  OR2_X1    g073(.A1(new_n274), .A2(KEYINPUT71), .ZN(new_n275));
  XOR2_X1   g074(.A(G197gat), .B(G204gat), .Z(new_n276));
  AOI21_X1  g075(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n275), .B(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND2_X1  g079(.A1(G226gat), .A2(G233gat), .ZN(new_n281));
  XOR2_X1   g080(.A(new_n281), .B(KEYINPUT72), .Z(new_n282));
  XNOR2_X1  g081(.A(KEYINPUT73), .B(KEYINPUT29), .ZN(new_n283));
  INV_X1    g082(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n282), .B1(new_n233), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n232), .A2(new_n223), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n286), .A2(new_n282), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT74), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n280), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n282), .B1(new_n286), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g090(.A(new_n291), .B1(new_n233), .B2(new_n282), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n279), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n289), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT30), .ZN(new_n296));
  XNOR2_X1  g095(.A(G8gat), .B(G36gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G64gat), .B(G92gat), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n297), .B(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n295), .A2(new_n296), .A3(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT40), .ZN(new_n302));
  XNOR2_X1  g101(.A(G141gat), .B(G148gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT2), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n304), .B1(G155gat), .B2(G162gat), .ZN(new_n305));
  INV_X1    g104(.A(G155gat), .ZN(new_n306));
  INV_X1    g105(.A(G162gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  OAI22_X1  g107(.A1(new_n303), .A2(new_n305), .B1(KEYINPUT75), .B2(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(G155gat), .B(G162gat), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n250), .A2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n314));
  NOR2_X1   g113(.A1(new_n248), .A2(new_n311), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(KEYINPUT76), .B(KEYINPUT3), .ZN(new_n318));
  NOR2_X1   g117(.A1(new_n311), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n319), .B1(KEYINPUT3), .B2(new_n311), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n314), .A2(new_n317), .B1(new_n320), .B2(new_n248), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT39), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  XOR2_X1   g124(.A(G57gat), .B(G85gat), .Z(new_n326));
  XNOR2_X1  g125(.A(G1gat), .B(G29gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(new_n326), .B(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT77), .B(KEYINPUT0), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  NAND2_X1  g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n248), .A2(new_n311), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n313), .A2(new_n322), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n324), .B1(new_n333), .B2(KEYINPUT84), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n334), .B1(KEYINPUT84), .B2(new_n333), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n335), .A2(new_n323), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n302), .B1(new_n331), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n296), .B1(new_n294), .B2(new_n299), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n338), .B1(new_n294), .B2(new_n299), .ZN(new_n339));
  INV_X1    g138(.A(new_n330), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n340), .B1(new_n323), .B2(new_n324), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n341), .B(KEYINPUT40), .C1(new_n323), .C2(new_n335), .ZN(new_n342));
  AND4_X1   g141(.A1(new_n301), .A2(new_n337), .A3(new_n339), .A4(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT5), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n320), .A2(new_n248), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n313), .A2(KEYINPUT4), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n315), .A2(new_n316), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n322), .B(new_n345), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(new_n322), .B1(new_n313), .B2(new_n332), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT5), .B1(new_n321), .B2(new_n322), .ZN(new_n352));
  NOR2_X1   g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n353), .A2(KEYINPUT85), .A3(new_n340), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n348), .A2(new_n344), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n349), .B1(new_n321), .B2(new_n322), .ZN(new_n356));
  OAI211_X1 g155(.A(new_n355), .B(new_n340), .C1(new_n356), .C2(new_n344), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT85), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(G78gat), .B(G106gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT79), .B(G22gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(G50gat), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n280), .B1(new_n319), .B2(new_n283), .ZN(new_n365));
  INV_X1    g164(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g165(.A(KEYINPUT3), .B1(new_n279), .B2(new_n290), .ZN(new_n367));
  NOR2_X1   g166(.A1(new_n367), .A2(new_n312), .ZN(new_n368));
  NAND2_X1  g167(.A1(G228gat), .A2(G233gat), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n366), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  OR3_X1    g170(.A1(new_n278), .A2(KEYINPUT81), .A3(new_n274), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT81), .B1(new_n278), .B2(new_n274), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n278), .A2(new_n274), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n372), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n318), .B1(new_n375), .B2(new_n284), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT82), .ZN(new_n377));
  OR3_X1    g176(.A1(new_n376), .A2(new_n377), .A3(new_n312), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n377), .B1(new_n376), .B2(new_n312), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n378), .A2(new_n365), .A3(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT83), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n369), .B(KEYINPUT80), .Z(new_n382));
  AND3_X1   g181(.A1(new_n380), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n371), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT31), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT31), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n387), .B(new_n371), .C1(new_n383), .C2(new_n384), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n364), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n386), .A2(new_n388), .A3(new_n364), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n343), .A2(new_n360), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n355), .B1(new_n356), .B2(new_n344), .ZN(new_n393));
  AOI21_X1  g192(.A(KEYINPUT6), .B1(new_n393), .B2(new_n330), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n360), .A2(new_n394), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n299), .B1(new_n294), .B2(KEYINPUT37), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n396), .A2(KEYINPUT38), .ZN(new_n397));
  OR2_X1    g196(.A1(new_n285), .A2(new_n288), .ZN(new_n398));
  OR2_X1    g197(.A1(new_n292), .A2(new_n279), .ZN(new_n399));
  OAI22_X1  g198(.A1(new_n280), .A2(new_n398), .B1(new_n399), .B2(KEYINPUT86), .ZN(new_n400));
  AND2_X1   g199(.A1(new_n399), .A2(KEYINPUT86), .ZN(new_n401));
  OAI21_X1  g200(.A(KEYINPUT37), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n397), .A2(new_n402), .B1(new_n295), .B2(new_n300), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n340), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n294), .A2(KEYINPUT37), .ZN(new_n405));
  OAI21_X1  g204(.A(KEYINPUT38), .B1(new_n405), .B2(new_n396), .ZN(new_n406));
  NAND4_X1  g205(.A1(new_n395), .A2(new_n403), .A3(new_n404), .A4(new_n406), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n273), .B1(new_n392), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n339), .A2(new_n301), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT78), .B1(new_n394), .B2(new_n357), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n330), .B1(new_n351), .B2(new_n352), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n411), .A2(new_n357), .A3(KEYINPUT78), .A4(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n404), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n409), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  INV_X1    g214(.A(new_n391), .ZN(new_n416));
  NOR2_X1   g215(.A1(new_n416), .A2(new_n389), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n269), .A2(new_n270), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(new_n420), .B1(new_n416), .B2(new_n389), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT35), .B1(new_n421), .B2(new_n415), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n390), .A2(new_n391), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n269), .A2(KEYINPUT87), .A3(new_n270), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT87), .B1(new_n269), .B2(new_n270), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  AND2_X1   g225(.A1(new_n339), .A2(new_n301), .ZN(new_n427));
  XOR2_X1   g226(.A(KEYINPUT88), .B(KEYINPUT35), .Z(new_n428));
  NOR2_X1   g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n395), .A2(new_n404), .ZN(new_n430));
  NAND4_X1  g229(.A1(new_n423), .A2(new_n426), .A3(new_n429), .A4(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n408), .A2(new_n418), .B1(new_n422), .B2(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT92), .ZN(new_n433));
  INV_X1    g232(.A(G8gat), .ZN(new_n434));
  AND2_X1   g233(.A1(G15gat), .A2(G22gat), .ZN(new_n435));
  NOR2_X1   g234(.A1(G15gat), .A2(G22gat), .ZN(new_n436));
  OAI21_X1  g235(.A(KEYINPUT91), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(G15gat), .ZN(new_n438));
  INV_X1    g237(.A(G22gat), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT91), .ZN(new_n441));
  NAND2_X1  g240(.A1(G15gat), .A2(G22gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(G1gat), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n444), .A2(KEYINPUT16), .ZN(new_n445));
  AND3_X1   g244(.A1(new_n437), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  AOI21_X1  g245(.A(G1gat), .B1(new_n437), .B2(new_n443), .ZN(new_n447));
  OAI211_X1 g246(.A(new_n433), .B(new_n434), .C1(new_n446), .C2(new_n447), .ZN(new_n448));
  NOR3_X1   g247(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT91), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n444), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n437), .A2(new_n443), .A3(new_n445), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n434), .ZN(new_n453));
  NAND2_X1  g252(.A1(KEYINPUT92), .A2(G8gat), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n451), .A2(new_n452), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n448), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(G29gat), .A2(G36gat), .ZN(new_n457));
  OAI21_X1  g256(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  AOI21_X1  g260(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n462));
  XNOR2_X1  g261(.A(KEYINPUT90), .B(G50gat), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n462), .B1(new_n463), .B2(G43gat), .ZN(new_n464));
  XNOR2_X1  g263(.A(G43gat), .B(G50gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n465), .A2(KEYINPUT15), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n461), .A2(new_n466), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT17), .B1(new_n467), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT17), .ZN(new_n471));
  AND2_X1   g270(.A1(new_n464), .A2(new_n466), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n471), .B(new_n468), .C1(new_n472), .C2(new_n461), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n456), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n448), .A2(KEYINPUT93), .A3(new_n455), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT93), .B1(new_n448), .B2(new_n455), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n467), .A2(new_n469), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(G229gat), .A2(G233gat), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n479), .A2(KEYINPUT95), .A3(KEYINPUT18), .A4(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT93), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n448), .A2(KEYINPUT93), .A3(new_n455), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n456), .A2(new_n473), .A3(new_n470), .ZN(new_n486));
  NAND4_X1  g285(.A1(new_n485), .A2(KEYINPUT18), .A3(new_n480), .A4(new_n486), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT95), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI22_X1  g288(.A1(new_n475), .A2(new_n476), .B1(new_n467), .B2(new_n469), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(new_n485), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n480), .B(KEYINPUT13), .ZN(new_n492));
  INV_X1    g291(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n491), .A2(new_n493), .ZN(new_n494));
  AND3_X1   g293(.A1(new_n481), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n485), .A2(new_n480), .A3(new_n486), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT18), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT94), .ZN(new_n499));
  XNOR2_X1  g298(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n500));
  XNOR2_X1  g299(.A(G113gat), .B(G141gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(G169gat), .B(G197gat), .Z(new_n503));
  XNOR2_X1  g302(.A(new_n502), .B(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(new_n504), .B(KEYINPUT12), .ZN(new_n505));
  OAI211_X1 g304(.A(new_n495), .B(new_n498), .C1(new_n499), .C2(new_n505), .ZN(new_n506));
  NAND4_X1  g305(.A1(new_n481), .A2(new_n498), .A3(new_n489), .A4(new_n494), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n481), .A2(new_n499), .A3(new_n489), .A4(new_n494), .ZN(new_n508));
  INV_X1    g307(.A(new_n505), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n506), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  AND2_X1   g311(.A1(G71gat), .A2(G78gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(G71gat), .A2(G78gat), .ZN(new_n514));
  NOR2_X1   g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G57gat), .B(G64gat), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n515), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(G57gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G64gat), .ZN(new_n520));
  INV_X1    g319(.A(G64gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n521), .A2(G57gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  XNOR2_X1  g322(.A(G71gat), .B(G78gat), .ZN(new_n524));
  INV_X1    g323(.A(new_n517), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n518), .A2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(KEYINPUT96), .B(KEYINPUT21), .Z(new_n528));
  OAI21_X1  g327(.A(new_n477), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  XNOR2_X1  g328(.A(KEYINPUT98), .B(KEYINPUT19), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n527), .A2(KEYINPUT21), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n531), .B1(new_n527), .B2(new_n528), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n532), .B1(new_n475), .B2(new_n476), .ZN(new_n533));
  AND3_X1   g332(.A1(new_n529), .A2(new_n530), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n530), .B1(new_n529), .B2(new_n533), .ZN(new_n535));
  XOR2_X1   g334(.A(G127gat), .B(G155gat), .Z(new_n536));
  OR3_X1    g335(.A1(new_n534), .A2(new_n535), .A3(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n536), .B1(new_n534), .B2(new_n535), .ZN(new_n538));
  NAND2_X1  g337(.A1(G231gat), .A2(G233gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n204), .ZN(new_n540));
  INV_X1    g339(.A(G211gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT97), .B(KEYINPUT20), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n537), .A2(new_n538), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n544), .B1(new_n537), .B2(new_n538), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT100), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT99), .ZN(new_n549));
  NAND2_X1  g348(.A1(G99gat), .A2(G106gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n550), .A2(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g350(.A1(G85gat), .A2(G92gat), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT7), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(G85gat), .ZN(new_n555));
  INV_X1    g354(.A(G92gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n551), .A2(new_n554), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(G99gat), .B(G106gat), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n559), .A2(new_n561), .ZN(new_n562));
  AND3_X1   g361(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT7), .B1(G85gat), .B2(G92gat), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI22_X1  g364(.A1(KEYINPUT8), .A2(new_n550), .B1(new_n555), .B2(new_n556), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g366(.A(new_n549), .B1(new_n562), .B2(new_n567), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n565), .A2(new_n560), .A3(new_n566), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT99), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n548), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n559), .A2(new_n561), .ZN(new_n572));
  AOI21_X1  g371(.A(KEYINPUT99), .B1(new_n572), .B2(new_n569), .ZN(new_n573));
  AND4_X1   g372(.A1(new_n551), .A2(new_n554), .A3(new_n557), .A4(new_n558), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n549), .B1(new_n574), .B2(new_n560), .ZN(new_n575));
  NOR3_X1   g374(.A1(new_n573), .A2(new_n575), .A3(KEYINPUT100), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n478), .B1(new_n571), .B2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n568), .A2(new_n548), .A3(new_n570), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT100), .B1(new_n573), .B2(new_n575), .ZN(new_n579));
  NAND4_X1  g378(.A1(new_n578), .A2(new_n579), .A3(new_n470), .A4(new_n473), .ZN(new_n580));
  NAND3_X1  g379(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n577), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G134gat), .B(G162gat), .Z(new_n583));
  OR2_X1    g382(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G190gat), .B(G218gat), .ZN(new_n585));
  AOI21_X1  g384(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n582), .A2(new_n583), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n584), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n587), .B1(new_n584), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n547), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g393(.A1(G230gat), .A2(G233gat), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  NOR3_X1   g395(.A1(new_n573), .A2(new_n527), .A3(new_n575), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n518), .A2(new_n526), .ZN(new_n598));
  AOI21_X1  g397(.A(new_n598), .B1(new_n569), .B2(new_n572), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n596), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(new_n598), .A2(new_n596), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  AOI21_X1  g401(.A(new_n602), .B1(new_n578), .B2(new_n579), .ZN(new_n603));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  AOI211_X1 g404(.A(KEYINPUT101), .B(new_n602), .C1(new_n578), .C2(new_n579), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n595), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(new_n599), .ZN(new_n608));
  NAND3_X1  g407(.A1(new_n568), .A2(new_n598), .A3(new_n570), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n607), .B1(new_n595), .B2(new_n610), .ZN(new_n611));
  XNOR2_X1  g410(.A(G176gat), .B(G204gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n612), .B(KEYINPUT103), .ZN(new_n613));
  XNOR2_X1  g412(.A(G120gat), .B(G148gat), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n613), .B(new_n614), .Z(new_n615));
  INV_X1    g414(.A(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(new_n605), .B2(new_n606), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n601), .B1(new_n571), .B2(new_n576), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n619), .A2(KEYINPUT101), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n604), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n620), .A2(new_n621), .A3(KEYINPUT102), .A4(new_n600), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n595), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n610), .ZN(new_n624));
  INV_X1    g423(.A(new_n595), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n616), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  AOI22_X1  g425(.A1(new_n611), .A2(new_n616), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n594), .A2(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n432), .A2(new_n512), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n410), .A2(new_n414), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(new_n631), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g431(.A1(new_n629), .A2(new_n427), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(G8gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n634), .A2(KEYINPUT42), .ZN(new_n635));
  XNOR2_X1  g434(.A(KEYINPUT16), .B(G8gat), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  MUX2_X1   g436(.A(new_n635), .B(KEYINPUT42), .S(new_n637), .Z(G1325gat));
  AOI21_X1  g437(.A(G15gat), .B1(new_n629), .B2(new_n426), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n273), .A2(G15gat), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n640), .B(KEYINPUT104), .Z(new_n641));
  AOI21_X1  g440(.A(new_n639), .B1(new_n629), .B2(new_n641), .ZN(G1326gat));
  NAND2_X1  g441(.A1(new_n629), .A2(new_n417), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(G22gat), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n629), .A2(new_n439), .A3(new_n417), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(G1327gat));
  NOR2_X1   g447(.A1(new_n432), .A2(new_n512), .ZN(new_n649));
  INV_X1    g448(.A(new_n547), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n650), .A2(new_n591), .A3(new_n627), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT106), .Z(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(new_n630), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n653), .A2(G29gat), .A3(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT45), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT44), .B1(new_n432), .B2(new_n592), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n422), .A2(new_n431), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n427), .A2(new_n360), .A3(new_n342), .A4(new_n337), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n407), .A2(new_n660), .A3(new_n423), .ZN(new_n661));
  INV_X1    g460(.A(new_n273), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n661), .A2(new_n418), .A3(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n592), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT44), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n658), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n611), .A2(new_n616), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n623), .A2(new_n626), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NOR3_X1   g469(.A1(new_n547), .A2(new_n512), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(G29gat), .B1(new_n672), .B2(new_n654), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n673), .ZN(G1328gat));
  NOR3_X1   g473(.A1(new_n653), .A2(G36gat), .A3(new_n409), .ZN(new_n675));
  XNOR2_X1  g474(.A(new_n675), .B(KEYINPUT46), .ZN(new_n676));
  OAI21_X1  g475(.A(G36gat), .B1(new_n672), .B2(new_n409), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n676), .A2(new_n677), .ZN(G1329gat));
  NAND3_X1  g477(.A1(new_n649), .A2(new_n426), .A3(new_n652), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT107), .ZN(new_n680));
  AOI22_X1  g479(.A1(new_n679), .A2(new_n259), .B1(new_n680), .B2(KEYINPUT47), .ZN(new_n681));
  NAND4_X1  g480(.A1(new_n667), .A2(G43gat), .A3(new_n273), .A4(new_n671), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n680), .A2(KEYINPUT47), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(G1330gat));
  NOR3_X1   g484(.A1(new_n432), .A2(KEYINPUT44), .A3(new_n592), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n664), .A2(new_n665), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n417), .B(new_n671), .C1(new_n686), .C2(new_n687), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n649), .A2(new_n652), .ZN(new_n689));
  NOR2_X1   g488(.A1(new_n423), .A2(new_n463), .ZN(new_n690));
  AOI22_X1  g489(.A1(new_n688), .A2(new_n463), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g491(.A1(new_n659), .A2(new_n663), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n693), .A2(new_n512), .A3(new_n594), .A4(new_n670), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n694), .A2(new_n654), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(new_n519), .ZN(G1332gat));
  XNOR2_X1  g495(.A(new_n427), .B(KEYINPUT108), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g498(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n700));
  AND2_X1   g499(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n699), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n702), .B1(new_n699), .B2(new_n700), .ZN(G1333gat));
  INV_X1    g502(.A(new_n426), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n694), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n273), .A2(G71gat), .ZN(new_n706));
  OAI22_X1  g505(.A1(new_n705), .A2(G71gat), .B1(new_n694), .B2(new_n706), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n707), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g507(.A1(new_n694), .A2(new_n423), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n709), .B(G78gat), .Z(G1335gat));
  NOR2_X1   g509(.A1(new_n547), .A2(new_n511), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n670), .ZN(new_n712));
  XNOR2_X1  g511(.A(new_n712), .B(KEYINPUT109), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n714), .B1(new_n658), .B2(new_n666), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G85gat), .B1(new_n716), .B2(new_n654), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n664), .A2(KEYINPUT51), .A3(new_n711), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT51), .B1(new_n664), .B2(new_n711), .ZN(new_n719));
  OR3_X1    g518(.A1(new_n718), .A2(new_n719), .A3(KEYINPUT110), .ZN(new_n720));
  OAI21_X1  g519(.A(KEYINPUT110), .B1(new_n718), .B2(new_n719), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n720), .A2(new_n670), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n630), .A2(new_n555), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n717), .B1(new_n722), .B2(new_n723), .ZN(G1336gat));
  NAND2_X1  g523(.A1(new_n697), .A2(new_n556), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(new_n670), .B(new_n726), .C1(new_n718), .C2(new_n719), .ZN(new_n727));
  INV_X1    g526(.A(KEYINPUT52), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n556), .B1(new_n715), .B2(new_n697), .ZN(new_n730));
  OAI21_X1  g529(.A(KEYINPUT111), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n667), .A2(new_n697), .A3(new_n713), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G92gat), .ZN(new_n733));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n734));
  NAND4_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n728), .A4(new_n727), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n556), .B1(new_n715), .B2(new_n427), .ZN(new_n736));
  NAND3_X1  g535(.A1(new_n693), .A2(new_n591), .A3(new_n711), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT51), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n737), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n664), .A2(KEYINPUT51), .A3(new_n711), .ZN(new_n740));
  AOI211_X1 g539(.A(new_n627), .B(new_n725), .C1(new_n739), .C2(new_n740), .ZN(new_n741));
  OAI21_X1  g540(.A(KEYINPUT52), .B1(new_n736), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n731), .A2(new_n735), .A3(new_n742), .ZN(G1337gat));
  OAI21_X1  g542(.A(G99gat), .B1(new_n716), .B2(new_n662), .ZN(new_n744));
  OR2_X1    g543(.A1(new_n704), .A2(G99gat), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n744), .B1(new_n722), .B2(new_n745), .ZN(G1338gat));
  OAI211_X1 g545(.A(new_n417), .B(new_n713), .C1(new_n686), .C2(new_n687), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G106gat), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n423), .A2(G106gat), .ZN(new_n749));
  OAI211_X1 g548(.A(new_n670), .B(new_n749), .C1(new_n718), .C2(new_n719), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT53), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT53), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n748), .A2(new_n753), .A3(new_n750), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n752), .A2(new_n754), .ZN(G1339gat));
  INV_X1    g554(.A(new_n669), .ZN(new_n756));
  AOI22_X1  g555(.A1(new_n619), .A2(KEYINPUT101), .B1(new_n610), .B2(new_n596), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n625), .B1(new_n757), .B2(new_n621), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT54), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n615), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  NAND4_X1  g559(.A1(new_n620), .A2(new_n621), .A3(new_n625), .A4(new_n600), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n757), .A2(KEYINPUT112), .A3(new_n625), .A4(new_n621), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(new_n764), .A3(KEYINPUT54), .ZN(new_n765));
  AND3_X1   g564(.A1(new_n618), .A2(new_n595), .A3(new_n622), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n760), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT55), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n756), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI211_X1 g568(.A(KEYINPUT55), .B(new_n760), .C1(new_n765), .C2(new_n766), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT113), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n623), .A2(KEYINPUT54), .A3(new_n764), .A4(new_n763), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n773), .A2(KEYINPUT113), .A3(KEYINPUT55), .A4(new_n760), .ZN(new_n774));
  NAND4_X1  g573(.A1(new_n769), .A2(new_n511), .A3(new_n772), .A4(new_n774), .ZN(new_n775));
  AND2_X1   g574(.A1(new_n489), .A2(new_n494), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n776), .A2(new_n498), .A3(new_n481), .A4(new_n505), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n490), .A2(new_n485), .A3(new_n492), .ZN(new_n778));
  OAI22_X1  g577(.A1(new_n778), .A2(KEYINPUT114), .B1(new_n479), .B2(new_n480), .ZN(new_n779));
  AND2_X1   g578(.A1(new_n778), .A2(KEYINPUT114), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n504), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n670), .A2(new_n777), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n775), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT116), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n775), .A2(KEYINPUT116), .A3(new_n782), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n592), .A3(new_n786), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n769), .A2(new_n772), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT115), .ZN(new_n789));
  AND3_X1   g588(.A1(new_n591), .A2(new_n777), .A3(new_n781), .ZN(new_n790));
  NAND4_X1  g589(.A1(new_n788), .A2(new_n789), .A3(new_n774), .A4(new_n790), .ZN(new_n791));
  NAND4_X1  g590(.A1(new_n790), .A2(new_n769), .A3(new_n774), .A4(new_n772), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT115), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n547), .B1(new_n787), .B2(new_n794), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n628), .A2(new_n511), .ZN(new_n796));
  NOR2_X1   g595(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n423), .A2(new_n426), .ZN(new_n798));
  NOR2_X1   g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NOR2_X1   g598(.A1(new_n697), .A2(new_n654), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G113gat), .B1(new_n801), .B2(new_n512), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n797), .A2(new_n654), .ZN(new_n803));
  INV_X1    g602(.A(new_n421), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n698), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n511), .A2(new_n235), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n802), .B1(new_n807), .B2(new_n808), .ZN(G1340gat));
  OAI21_X1  g608(.A(G120gat), .B1(new_n801), .B2(new_n627), .ZN(new_n810));
  NOR2_X1   g609(.A1(new_n627), .A2(G120gat), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n803), .A2(new_n804), .A3(new_n698), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(new_n813), .B(KEYINPUT117), .ZN(G1341gat));
  INV_X1    g613(.A(G127gat), .ZN(new_n815));
  NOR3_X1   g614(.A1(new_n801), .A2(new_n815), .A3(new_n650), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n806), .A2(new_n547), .A3(new_n698), .ZN(new_n817));
  AOI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n815), .ZN(G1342gat));
  NOR2_X1   g617(.A1(new_n427), .A2(new_n592), .ZN(new_n819));
  INV_X1    g618(.A(new_n819), .ZN(new_n820));
  OR4_X1    g619(.A1(KEYINPUT56), .A2(new_n805), .A3(G134gat), .A4(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(G134gat), .B1(new_n801), .B2(new_n592), .ZN(new_n822));
  OR2_X1    g621(.A1(new_n820), .A2(G134gat), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT56), .B1(new_n805), .B2(new_n823), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n821), .A2(new_n822), .A3(new_n824), .ZN(G1343gat));
  NOR2_X1   g624(.A1(new_n423), .A2(new_n273), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n512), .A2(G141gat), .ZN(new_n827));
  AND4_X1   g626(.A1(new_n698), .A2(new_n803), .A3(new_n826), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT120), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT57), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n831), .B(new_n417), .C1(new_n795), .C2(new_n796), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n781), .B1(new_n507), .B2(new_n509), .ZN(new_n833));
  OAI21_X1  g632(.A(KEYINPUT118), .B1(new_n833), .B2(new_n627), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT118), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n670), .A2(new_n777), .A3(new_n835), .A4(new_n781), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n775), .A2(new_n834), .A3(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(new_n592), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n794), .A2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n796), .B1(new_n839), .B2(new_n650), .ZN(new_n840));
  OAI21_X1  g639(.A(KEYINPUT57), .B1(new_n840), .B2(new_n423), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n697), .A2(new_n654), .A3(new_n273), .ZN(new_n842));
  NAND4_X1  g641(.A1(new_n832), .A2(new_n841), .A3(new_n511), .A4(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(KEYINPUT58), .B1(new_n843), .B2(G141gat), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n803), .A2(new_n698), .A3(new_n826), .ZN(new_n845));
  INV_X1    g644(.A(new_n827), .ZN(new_n846));
  OAI21_X1  g645(.A(KEYINPUT120), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n830), .A2(new_n844), .A3(new_n847), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  AND3_X1   g648(.A1(new_n843), .A2(new_n849), .A3(G141gat), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n849), .B1(new_n843), .B2(G141gat), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n850), .A2(new_n851), .A3(new_n828), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT58), .ZN(new_n853));
  OAI21_X1  g652(.A(new_n848), .B1(new_n852), .B2(new_n853), .ZN(G1344gat));
  INV_X1    g653(.A(G148gat), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n670), .A2(new_n855), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n845), .A2(KEYINPUT121), .A3(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(KEYINPUT121), .B1(new_n845), .B2(new_n856), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n860));
  INV_X1    g659(.A(new_n796), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n591), .B1(new_n783), .B2(new_n784), .ZN(new_n862));
  AOI22_X1  g661(.A1(new_n862), .A2(new_n786), .B1(new_n793), .B2(new_n791), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n861), .B1(new_n863), .B2(new_n547), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n831), .B1(new_n864), .B2(new_n417), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n838), .A2(new_n792), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n650), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n861), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n831), .A3(new_n417), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n866), .A2(new_n670), .A3(new_n842), .A4(new_n870), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n860), .B1(new_n871), .B2(G148gat), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n832), .A2(new_n841), .A3(new_n842), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  AOI211_X1 g673(.A(KEYINPUT59), .B(new_n855), .C1(new_n874), .C2(new_n670), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n859), .B1(new_n872), .B2(new_n875), .ZN(G1345gat));
  NOR3_X1   g675(.A1(new_n873), .A2(new_n306), .A3(new_n650), .ZN(new_n877));
  OR2_X1    g676(.A1(new_n845), .A2(new_n650), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n878), .B2(new_n306), .ZN(G1346gat));
  OAI21_X1  g678(.A(G162gat), .B1(new_n873), .B2(new_n592), .ZN(new_n880));
  NAND4_X1  g679(.A1(new_n803), .A2(new_n307), .A3(new_n819), .A4(new_n826), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g681(.A(new_n882), .B(KEYINPUT122), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n630), .A2(new_n409), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n799), .A2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G169gat), .B1(new_n885), .B2(new_n512), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n797), .A2(new_n630), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n698), .A2(new_n421), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n512), .A2(G169gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n889), .B2(new_n890), .ZN(G1348gat));
  INV_X1    g690(.A(G176gat), .ZN(new_n892));
  NOR3_X1   g691(.A1(new_n885), .A2(new_n892), .A3(new_n627), .ZN(new_n893));
  INV_X1    g692(.A(new_n889), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(new_n670), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n893), .B1(new_n892), .B2(new_n895), .ZN(G1349gat));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n226), .A3(new_n547), .ZN(new_n897));
  OAI21_X1  g696(.A(G183gat), .B1(new_n885), .B2(new_n650), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(KEYINPUT60), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT60), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(new_n901), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(G1350gat));
  NAND3_X1  g702(.A1(new_n799), .A2(new_n591), .A3(new_n884), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G190gat), .ZN(new_n905));
  OAI21_X1  g704(.A(KEYINPUT123), .B1(new_n905), .B2(KEYINPUT61), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(KEYINPUT61), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT123), .ZN(new_n908));
  INV_X1    g707(.A(KEYINPUT61), .ZN(new_n909));
  NAND4_X1  g708(.A1(new_n904), .A2(new_n908), .A3(new_n909), .A4(G190gat), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n894), .A2(new_n205), .A3(new_n591), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(G1351gat));
  AND2_X1   g712(.A1(new_n826), .A2(new_n697), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n887), .A2(new_n914), .ZN(new_n915));
  OR3_X1    g714(.A1(new_n915), .A2(G197gat), .A3(new_n512), .ZN(new_n916));
  AOI211_X1 g715(.A(KEYINPUT57), .B(new_n423), .C1(new_n868), .C2(new_n861), .ZN(new_n917));
  OAI21_X1  g716(.A(KEYINPUT124), .B1(new_n865), .B2(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT124), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n775), .A2(KEYINPUT116), .A3(new_n782), .ZN(new_n920));
  AOI21_X1  g719(.A(KEYINPUT116), .B1(new_n775), .B2(new_n782), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n920), .A2(new_n921), .A3(new_n591), .ZN(new_n922));
  INV_X1    g721(.A(new_n794), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n650), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n423), .B1(new_n924), .B2(new_n861), .ZN(new_n925));
  OAI211_X1 g724(.A(new_n919), .B(new_n870), .C1(new_n925), .C2(new_n831), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n884), .A2(new_n662), .ZN(new_n927));
  INV_X1    g726(.A(new_n927), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n918), .A2(new_n511), .A3(new_n926), .A4(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT125), .ZN(new_n930));
  AND2_X1   g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G197gat), .B1(new_n929), .B2(new_n930), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n916), .B1(new_n931), .B2(new_n932), .ZN(G1352gat));
  INV_X1    g732(.A(KEYINPUT126), .ZN(new_n934));
  INV_X1    g733(.A(new_n915), .ZN(new_n935));
  NOR2_X1   g734(.A1(new_n627), .A2(G204gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n934), .B1(new_n937), .B2(KEYINPUT62), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n918), .A2(new_n926), .A3(new_n928), .ZN(new_n939));
  OAI21_X1  g738(.A(G204gat), .B1(new_n939), .B2(new_n627), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n935), .A2(KEYINPUT126), .A3(new_n941), .A4(new_n936), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n937), .A2(KEYINPUT62), .ZN(new_n943));
  NAND4_X1  g742(.A1(new_n938), .A2(new_n940), .A3(new_n942), .A4(new_n943), .ZN(G1353gat));
  NAND3_X1  g743(.A1(new_n935), .A2(new_n541), .A3(new_n547), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n927), .A2(new_n650), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n870), .B(new_n946), .C1(new_n925), .C2(new_n831), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n541), .B1(new_n947), .B2(KEYINPUT127), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT127), .ZN(new_n949));
  NAND4_X1  g748(.A1(new_n866), .A2(new_n949), .A3(new_n870), .A4(new_n946), .ZN(new_n950));
  AND3_X1   g749(.A1(new_n948), .A2(KEYINPUT63), .A3(new_n950), .ZN(new_n951));
  AOI21_X1  g750(.A(KEYINPUT63), .B1(new_n948), .B2(new_n950), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n945), .B1(new_n951), .B2(new_n952), .ZN(G1354gat));
  INV_X1    g752(.A(G218gat), .ZN(new_n954));
  NOR3_X1   g753(.A1(new_n939), .A2(new_n954), .A3(new_n592), .ZN(new_n955));
  AOI21_X1  g754(.A(G218gat), .B1(new_n935), .B2(new_n591), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n955), .A2(new_n956), .ZN(G1355gat));
endmodule


