

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750;

  XNOR2_X1 U367 ( .A(KEYINPUT66), .B(G131), .ZN(n509) );
  XNOR2_X2 U368 ( .A(n460), .B(n434), .ZN(n657) );
  INV_X1 U369 ( .A(G953), .ZN(n744) );
  AND2_X2 U370 ( .A1(n616), .A2(n356), .ZN(n344) );
  NOR2_X1 U371 ( .A1(n654), .A2(G902), .ZN(n399) );
  INV_X2 U372 ( .A(n622), .ZN(n616) );
  NOR2_X1 U373 ( .A1(n740), .A2(n404), .ZN(n403) );
  XNOR2_X1 U374 ( .A(n570), .B(KEYINPUT39), .ZN(n607) );
  NOR2_X1 U375 ( .A1(n588), .A2(n587), .ZN(n631) );
  NAND2_X1 U376 ( .A1(n585), .A2(n705), .ZN(n570) );
  XNOR2_X1 U377 ( .A(n397), .B(KEYINPUT1), .ZN(n522) );
  XNOR2_X1 U378 ( .A(n399), .B(n350), .ZN(n521) );
  NOR2_X1 U379 ( .A1(n416), .A2(G953), .ZN(n415) );
  XNOR2_X1 U380 ( .A(n488), .B(KEYINPUT4), .ZN(n470) );
  XNOR2_X1 U381 ( .A(G122), .B(G104), .ZN(n507) );
  XOR2_X1 U382 ( .A(KEYINPUT77), .B(KEYINPUT34), .Z(n486) );
  XNOR2_X1 U383 ( .A(KEYINPUT82), .B(KEYINPUT8), .ZN(n417) );
  NOR2_X2 U384 ( .A1(n374), .A2(n375), .ZN(n656) );
  NAND2_X2 U385 ( .A1(n405), .A2(n401), .ZN(n374) );
  XNOR2_X1 U386 ( .A(n477), .B(n476), .ZN(n569) );
  NAND2_X1 U387 ( .A1(n419), .A2(n353), .ZN(n418) );
  NOR2_X2 U388 ( .A1(n727), .A2(n623), .ZN(n375) );
  AND2_X1 U389 ( .A1(n606), .A2(n605), .ZN(n413) );
  INV_X1 U390 ( .A(G237), .ZN(n475) );
  XNOR2_X1 U391 ( .A(n415), .B(n417), .ZN(n398) );
  INV_X1 U392 ( .A(G234), .ZN(n416) );
  INV_X1 U393 ( .A(n419), .ZN(n404) );
  XNOR2_X1 U394 ( .A(n387), .B(n386), .ZN(n709) );
  INV_X1 U395 ( .A(KEYINPUT103), .ZN(n386) );
  INV_X1 U396 ( .A(KEYINPUT19), .ZN(n377) );
  NAND2_X1 U397 ( .A1(n381), .A2(KEYINPUT19), .ZN(n380) );
  XOR2_X1 U398 ( .A(KEYINPUT81), .B(G110), .Z(n439) );
  XNOR2_X1 U399 ( .A(n392), .B(n732), .ZN(n649) );
  NAND2_X1 U400 ( .A1(n371), .A2(n373), .ZN(n364) );
  NOR2_X1 U401 ( .A1(n375), .A2(n372), .ZN(n371) );
  INV_X1 U402 ( .A(G475), .ZN(n372) );
  NAND2_X1 U403 ( .A1(n368), .A2(n370), .ZN(n360) );
  NOR2_X1 U404 ( .A1(n375), .A2(n369), .ZN(n368) );
  INV_X1 U405 ( .A(G210), .ZN(n369) );
  NOR2_X1 U406 ( .A1(G953), .A2(G237), .ZN(n500) );
  INV_X1 U407 ( .A(KEYINPUT64), .ZN(n423) );
  XNOR2_X1 U408 ( .A(G902), .B(KEYINPUT15), .ZN(n618) );
  XOR2_X1 U409 ( .A(KEYINPUT72), .B(KEYINPUT5), .Z(n454) );
  XOR2_X1 U410 ( .A(G137), .B(G116), .Z(n455) );
  XNOR2_X1 U411 ( .A(G113), .B(KEYINPUT3), .ZN(n458) );
  XOR2_X1 U412 ( .A(KEYINPUT11), .B(KEYINPUT96), .Z(n502) );
  INV_X1 U413 ( .A(n507), .ZN(n508) );
  XNOR2_X1 U414 ( .A(G113), .B(G143), .ZN(n503) );
  XOR2_X1 U415 ( .A(KEYINPUT12), .B(G140), .Z(n504) );
  XNOR2_X1 U416 ( .A(n429), .B(G110), .ZN(n469) );
  INV_X1 U417 ( .A(KEYINPUT67), .ZN(n429) );
  NAND2_X1 U418 ( .A1(n422), .A2(n420), .ZN(n419) );
  NAND2_X1 U419 ( .A1(n618), .A2(n423), .ZN(n422) );
  NAND2_X1 U420 ( .A1(n619), .A2(n421), .ZN(n420) );
  NAND2_X1 U421 ( .A1(KEYINPUT2), .A2(n423), .ZN(n421) );
  XNOR2_X1 U422 ( .A(KEYINPUT88), .B(KEYINPUT17), .ZN(n472) );
  XNOR2_X1 U423 ( .A(KEYINPUT18), .B(KEYINPUT76), .ZN(n471) );
  NAND2_X1 U424 ( .A1(G234), .A2(G237), .ZN(n480) );
  INV_X1 U425 ( .A(KEYINPUT48), .ZN(n411) );
  XNOR2_X1 U426 ( .A(n388), .B(n346), .ZN(n532) );
  INV_X1 U427 ( .A(G902), .ZN(n514) );
  XNOR2_X1 U428 ( .A(n390), .B(n467), .ZN(n732) );
  XNOR2_X1 U429 ( .A(n391), .B(n495), .ZN(n390) );
  XNOR2_X1 U430 ( .A(n507), .B(KEYINPUT16), .ZN(n391) );
  XNOR2_X1 U431 ( .A(G134), .B(G122), .ZN(n492) );
  XOR2_X1 U432 ( .A(G116), .B(G107), .Z(n495) );
  NAND2_X1 U433 ( .A1(n744), .A2(G227), .ZN(n426) );
  XNOR2_X1 U434 ( .A(KEYINPUT74), .B(G107), .ZN(n430) );
  NAND2_X1 U435 ( .A1(n378), .A2(n349), .ZN(n376) );
  BUF_X1 U436 ( .A(n522), .Z(n689) );
  XNOR2_X1 U437 ( .A(n520), .B(KEYINPUT92), .ZN(n389) );
  XNOR2_X1 U438 ( .A(n692), .B(n464), .ZN(n595) );
  XNOR2_X1 U439 ( .A(n383), .B(n352), .ZN(n544) );
  XNOR2_X1 U440 ( .A(n519), .B(KEYINPUT104), .ZN(n384) );
  NAND2_X1 U441 ( .A1(n367), .A2(n365), .ZN(n643) );
  NOR2_X1 U442 ( .A1(n375), .A2(n366), .ZN(n365) );
  INV_X1 U443 ( .A(G472), .ZN(n366) );
  XNOR2_X1 U444 ( .A(n443), .B(n738), .ZN(n654) );
  NOR2_X1 U445 ( .A1(n345), .A2(n375), .ZN(n685) );
  INV_X1 U446 ( .A(G140), .ZN(n635) );
  INV_X1 U447 ( .A(G134), .ZN(n637) );
  INV_X1 U448 ( .A(KEYINPUT60), .ZN(n361) );
  XNOR2_X1 U449 ( .A(n364), .B(n354), .ZN(n363) );
  INV_X1 U450 ( .A(KEYINPUT56), .ZN(n357) );
  XNOR2_X1 U451 ( .A(n360), .B(n355), .ZN(n359) );
  AND2_X1 U452 ( .A1(n424), .A2(n617), .ZN(n345) );
  XOR2_X1 U453 ( .A(n516), .B(n515), .Z(n346) );
  XOR2_X1 U454 ( .A(G101), .B(G119), .Z(n347) );
  NOR2_X1 U455 ( .A1(n744), .A2(n561), .ZN(n348) );
  AND2_X1 U456 ( .A1(n706), .A2(n377), .ZN(n349) );
  XNOR2_X1 U457 ( .A(n447), .B(n446), .ZN(n350) );
  AND2_X1 U458 ( .A1(n664), .A2(n538), .ZN(n351) );
  XNOR2_X1 U459 ( .A(KEYINPUT65), .B(KEYINPUT22), .ZN(n352) );
  INV_X1 U460 ( .A(n706), .ZN(n381) );
  NAND2_X1 U461 ( .A1(n617), .A2(KEYINPUT64), .ZN(n353) );
  XOR2_X1 U462 ( .A(n651), .B(n650), .Z(n354) );
  XOR2_X1 U463 ( .A(n649), .B(n648), .Z(n355) );
  AND2_X1 U464 ( .A1(n619), .A2(n423), .ZN(n356) );
  XNOR2_X1 U465 ( .A(n358), .B(n357), .ZN(G51) );
  NAND2_X1 U466 ( .A1(n359), .A2(n644), .ZN(n358) );
  XNOR2_X1 U467 ( .A(n362), .B(n361), .ZN(G60) );
  NAND2_X1 U468 ( .A1(n363), .A2(n644), .ZN(n362) );
  INV_X1 U469 ( .A(n374), .ZN(n367) );
  INV_X1 U470 ( .A(n374), .ZN(n370) );
  INV_X1 U471 ( .A(n374), .ZN(n373) );
  XNOR2_X1 U472 ( .A(n394), .B(n474), .ZN(n393) );
  NAND2_X1 U473 ( .A1(n344), .A2(n400), .ZN(n405) );
  NAND2_X1 U474 ( .A1(n402), .A2(n418), .ZN(n401) );
  NAND2_X1 U475 ( .A1(n379), .A2(n376), .ZN(n590) );
  INV_X1 U476 ( .A(n569), .ZN(n378) );
  AND2_X1 U477 ( .A1(n382), .A2(n380), .ZN(n379) );
  NAND2_X1 U478 ( .A1(n569), .A2(KEYINPUT19), .ZN(n382) );
  NAND2_X1 U479 ( .A1(n590), .A2(n484), .ZN(n485) );
  NAND2_X1 U480 ( .A1(n544), .A2(n543), .ZN(n546) );
  NAND2_X1 U481 ( .A1(n385), .A2(n384), .ZN(n383) );
  INV_X1 U482 ( .A(n520), .ZN(n385) );
  NAND2_X1 U483 ( .A1(n536), .A2(n532), .ZN(n387) );
  AND2_X1 U484 ( .A1(n651), .A2(n514), .ZN(n388) );
  OR2_X1 U485 ( .A1(n389), .A2(n531), .ZN(n669) );
  NOR2_X2 U486 ( .A1(n712), .A2(n389), .ZN(n487) );
  XNOR2_X1 U487 ( .A(n395), .B(n393), .ZN(n392) );
  XNOR2_X1 U488 ( .A(n469), .B(KEYINPUT75), .ZN(n394) );
  XNOR2_X1 U489 ( .A(n470), .B(n396), .ZN(n395) );
  XNOR2_X1 U490 ( .A(n473), .B(n468), .ZN(n396) );
  NAND2_X1 U491 ( .A1(n529), .A2(n397), .ZN(n530) );
  XNOR2_X1 U492 ( .A(n397), .B(n580), .ZN(n581) );
  XNOR2_X2 U493 ( .A(n435), .B(G469), .ZN(n397) );
  NAND2_X1 U494 ( .A1(n398), .A2(G221), .ZN(n437) );
  AND2_X1 U495 ( .A1(n398), .A2(G217), .ZN(n491) );
  NOR2_X2 U496 ( .A1(n521), .A2(n686), .ZN(n529) );
  XNOR2_X2 U497 ( .A(n620), .B(n615), .ZN(n740) );
  NAND2_X2 U498 ( .A1(n410), .A2(n614), .ZN(n620) );
  NAND2_X1 U499 ( .A1(n400), .A2(n616), .ZN(n424) );
  INV_X1 U500 ( .A(n740), .ZN(n400) );
  NAND2_X1 U501 ( .A1(n403), .A2(n616), .ZN(n402) );
  NAND2_X1 U502 ( .A1(n406), .A2(n547), .ZN(n548) );
  XNOR2_X1 U503 ( .A(n408), .B(n407), .ZN(n406) );
  INV_X1 U504 ( .A(KEYINPUT86), .ZN(n407) );
  NAND2_X1 U505 ( .A1(n409), .A2(n351), .ZN(n408) );
  NAND2_X1 U506 ( .A1(n550), .A2(KEYINPUT44), .ZN(n409) );
  XNOR2_X2 U507 ( .A(n412), .B(n411), .ZN(n410) );
  NAND2_X1 U508 ( .A1(n414), .A2(n413), .ZN(n412) );
  XNOR2_X1 U509 ( .A(n584), .B(KEYINPUT46), .ZN(n414) );
  BUF_X1 U510 ( .A(n622), .Z(n727) );
  INV_X1 U511 ( .A(KEYINPUT80), .ZN(n589) );
  XNOR2_X1 U512 ( .A(n455), .B(KEYINPUT71), .ZN(n456) );
  INV_X1 U513 ( .A(KEYINPUT2), .ZN(n617) );
  XNOR2_X1 U514 ( .A(n457), .B(n456), .ZN(n459) );
  XNOR2_X1 U515 ( .A(n572), .B(n571), .ZN(n652) );
  XNOR2_X2 U516 ( .A(G143), .B(G128), .ZN(n488) );
  XNOR2_X1 U517 ( .A(n509), .B(n637), .ZN(n425) );
  XNOR2_X2 U518 ( .A(n470), .B(n425), .ZN(n739) );
  XNOR2_X2 U519 ( .A(n739), .B(G146), .ZN(n460) );
  XNOR2_X1 U520 ( .A(G104), .B(G101), .ZN(n427) );
  XNOR2_X1 U521 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U522 ( .A(n635), .B(G137), .ZN(n442) );
  XNOR2_X1 U523 ( .A(n428), .B(n442), .ZN(n433) );
  INV_X1 U524 ( .A(n469), .ZN(n431) );
  XNOR2_X1 U525 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U526 ( .A(n433), .B(n432), .ZN(n434) );
  OR2_X2 U527 ( .A1(n657), .A2(G902), .ZN(n435) );
  XOR2_X1 U528 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n436) );
  XNOR2_X1 U529 ( .A(n437), .B(n436), .ZN(n441) );
  XNOR2_X1 U530 ( .A(G119), .B(G128), .ZN(n438) );
  XNOR2_X1 U531 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U532 ( .A(n441), .B(n440), .ZN(n443) );
  XNOR2_X1 U533 ( .A(G146), .B(G125), .ZN(n468) );
  XNOR2_X1 U534 ( .A(n468), .B(KEYINPUT10), .ZN(n511) );
  XNOR2_X1 U535 ( .A(n511), .B(n442), .ZN(n738) );
  XOR2_X1 U536 ( .A(KEYINPUT93), .B(KEYINPUT20), .Z(n445) );
  NAND2_X1 U537 ( .A1(G234), .A2(n618), .ZN(n444) );
  XNOR2_X1 U538 ( .A(n445), .B(n444), .ZN(n448) );
  NAND2_X1 U539 ( .A1(G217), .A2(n448), .ZN(n447) );
  INV_X1 U540 ( .A(KEYINPUT25), .ZN(n446) );
  NAND2_X1 U541 ( .A1(n448), .A2(G221), .ZN(n449) );
  XNOR2_X1 U542 ( .A(n449), .B(KEYINPUT21), .ZN(n450) );
  XNOR2_X1 U543 ( .A(n450), .B(KEYINPUT94), .ZN(n686) );
  NAND2_X1 U544 ( .A1(n522), .A2(n529), .ZN(n452) );
  INV_X1 U545 ( .A(KEYINPUT70), .ZN(n451) );
  XNOR2_X2 U546 ( .A(n452), .B(n451), .ZN(n526) );
  NAND2_X1 U547 ( .A1(n500), .A2(G210), .ZN(n453) );
  XNOR2_X1 U548 ( .A(n454), .B(n453), .ZN(n457) );
  XNOR2_X1 U549 ( .A(n347), .B(n458), .ZN(n467) );
  XNOR2_X1 U550 ( .A(n459), .B(n467), .ZN(n461) );
  XNOR2_X1 U551 ( .A(n460), .B(n461), .ZN(n641) );
  NAND2_X1 U552 ( .A1(n641), .A2(n514), .ZN(n462) );
  XNOR2_X2 U553 ( .A(n462), .B(G472), .ZN(n692) );
  INV_X1 U554 ( .A(KEYINPUT102), .ZN(n463) );
  XNOR2_X1 U555 ( .A(n463), .B(KEYINPUT6), .ZN(n464) );
  NAND2_X1 U556 ( .A1(n526), .A2(n595), .ZN(n466) );
  XNOR2_X1 U557 ( .A(KEYINPUT107), .B(KEYINPUT33), .ZN(n465) );
  XNOR2_X1 U558 ( .A(n466), .B(n465), .ZN(n712) );
  XNOR2_X1 U559 ( .A(n472), .B(n471), .ZN(n474) );
  NAND2_X1 U560 ( .A1(n744), .A2(G224), .ZN(n473) );
  NAND2_X1 U561 ( .A1(n649), .A2(n618), .ZN(n477) );
  NAND2_X1 U562 ( .A1(n514), .A2(n475), .ZN(n478) );
  NAND2_X1 U563 ( .A1(n478), .A2(G210), .ZN(n476) );
  NAND2_X1 U564 ( .A1(n478), .A2(G214), .ZN(n706) );
  NOR2_X1 U565 ( .A1(G898), .A2(n744), .ZN(n479) );
  XNOR2_X1 U566 ( .A(KEYINPUT91), .B(n479), .ZN(n734) );
  XOR2_X1 U567 ( .A(KEYINPUT69), .B(KEYINPUT14), .Z(n481) );
  XNOR2_X1 U568 ( .A(n481), .B(n480), .ZN(n482) );
  NAND2_X1 U569 ( .A1(G902), .A2(n482), .ZN(n561) );
  OR2_X1 U570 ( .A1(n734), .A2(n561), .ZN(n483) );
  NAND2_X1 U571 ( .A1(G952), .A2(n482), .ZN(n718) );
  OR2_X1 U572 ( .A1(n718), .A2(G953), .ZN(n564) );
  NAND2_X1 U573 ( .A1(n483), .A2(n564), .ZN(n484) );
  XNOR2_X2 U574 ( .A(n485), .B(KEYINPUT0), .ZN(n520) );
  XNOR2_X1 U575 ( .A(n487), .B(n486), .ZN(n517) );
  XOR2_X1 U576 ( .A(KEYINPUT100), .B(KEYINPUT99), .Z(n489) );
  XNOR2_X1 U577 ( .A(n488), .B(n489), .ZN(n490) );
  XNOR2_X1 U578 ( .A(n491), .B(n490), .ZN(n497) );
  XOR2_X1 U579 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n493) );
  XNOR2_X1 U580 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U581 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U582 ( .A(n497), .B(n496), .ZN(n624) );
  NAND2_X1 U583 ( .A1(n624), .A2(n514), .ZN(n499) );
  INV_X1 U584 ( .A(G478), .ZN(n498) );
  XNOR2_X1 U585 ( .A(n499), .B(n498), .ZN(n536) );
  NAND2_X1 U586 ( .A1(G214), .A2(n500), .ZN(n501) );
  XNOR2_X1 U587 ( .A(n502), .B(n501), .ZN(n506) );
  XNOR2_X1 U588 ( .A(n504), .B(n503), .ZN(n505) );
  XOR2_X1 U589 ( .A(n506), .B(n505), .Z(n513) );
  XNOR2_X1 U590 ( .A(n509), .B(n508), .ZN(n510) );
  XNOR2_X1 U591 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U592 ( .A(n513), .B(n512), .ZN(n651) );
  XOR2_X1 U593 ( .A(KEYINPUT98), .B(KEYINPUT13), .Z(n516) );
  XNOR2_X1 U594 ( .A(KEYINPUT97), .B(G475), .ZN(n515) );
  NOR2_X1 U595 ( .A1(n536), .A2(n532), .ZN(n586) );
  NAND2_X1 U596 ( .A1(n517), .A2(n586), .ZN(n518) );
  XNOR2_X1 U597 ( .A(n518), .B(KEYINPUT35), .ZN(n550) );
  NOR2_X1 U598 ( .A1(n709), .A2(n686), .ZN(n519) );
  BUF_X1 U599 ( .A(n521), .Z(n577) );
  XOR2_X1 U600 ( .A(KEYINPUT105), .B(n577), .Z(n687) );
  INV_X1 U601 ( .A(n687), .ZN(n523) );
  INV_X1 U602 ( .A(n689), .ZN(n601) );
  NAND2_X1 U603 ( .A1(n523), .A2(n601), .ZN(n524) );
  NOR2_X1 U604 ( .A1(n524), .A2(n595), .ZN(n525) );
  NAND2_X1 U605 ( .A1(n544), .A2(n525), .ZN(n664) );
  BUF_X1 U606 ( .A(n526), .Z(n527) );
  NAND2_X1 U607 ( .A1(n527), .A2(n692), .ZN(n696) );
  NOR2_X1 U608 ( .A1(n696), .A2(n520), .ZN(n528) );
  XNOR2_X1 U609 ( .A(n528), .B(KEYINPUT31), .ZN(n632) );
  XNOR2_X2 U610 ( .A(n530), .B(KEYINPUT95), .ZN(n559) );
  INV_X1 U611 ( .A(n692), .ZN(n578) );
  NAND2_X1 U612 ( .A1(n559), .A2(n578), .ZN(n531) );
  NAND2_X1 U613 ( .A1(n632), .A2(n669), .ZN(n537) );
  INV_X1 U614 ( .A(n532), .ZN(n535) );
  NAND2_X1 U615 ( .A1(n536), .A2(n535), .ZN(n534) );
  INV_X1 U616 ( .A(KEYINPUT101), .ZN(n533) );
  XNOR2_X1 U617 ( .A(n534), .B(n533), .ZN(n666) );
  OR2_X1 U618 ( .A1(n536), .A2(n535), .ZN(n675) );
  NAND2_X1 U619 ( .A1(n666), .A2(n675), .ZN(n701) );
  NAND2_X1 U620 ( .A1(n537), .A2(n701), .ZN(n538) );
  NAND2_X1 U621 ( .A1(n578), .A2(n577), .ZN(n539) );
  NOR2_X1 U622 ( .A1(n689), .A2(n539), .ZN(n540) );
  NAND2_X1 U623 ( .A1(n544), .A2(n540), .ZN(n541) );
  XNOR2_X1 U624 ( .A(n541), .B(KEYINPUT106), .ZN(n749) );
  NAND2_X1 U625 ( .A1(n687), .A2(n689), .ZN(n542) );
  NOR2_X1 U626 ( .A1(n542), .A2(n595), .ZN(n543) );
  XNOR2_X1 U627 ( .A(KEYINPUT78), .B(KEYINPUT32), .ZN(n545) );
  XNOR2_X1 U628 ( .A(n546), .B(n545), .ZN(n634) );
  NAND2_X1 U629 ( .A1(n749), .A2(n634), .ZN(n549) );
  NAND2_X1 U630 ( .A1(n549), .A2(KEYINPUT44), .ZN(n547) );
  XNOR2_X1 U631 ( .A(n548), .B(KEYINPUT85), .ZN(n556) );
  NOR2_X1 U632 ( .A1(n549), .A2(KEYINPUT44), .ZN(n553) );
  BUF_X1 U633 ( .A(n550), .Z(n551) );
  INV_X1 U634 ( .A(n551), .ZN(n552) );
  NAND2_X1 U635 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U636 ( .A(n554), .B(KEYINPUT68), .ZN(n555) );
  NAND2_X1 U637 ( .A1(n556), .A2(n555), .ZN(n558) );
  XOR2_X1 U638 ( .A(KEYINPUT84), .B(KEYINPUT45), .Z(n557) );
  XNOR2_X1 U639 ( .A(n558), .B(n557), .ZN(n622) );
  INV_X1 U640 ( .A(KEYINPUT83), .ZN(n615) );
  XNOR2_X1 U641 ( .A(n559), .B(KEYINPUT110), .ZN(n567) );
  NAND2_X1 U642 ( .A1(n692), .A2(n706), .ZN(n560) );
  XNOR2_X1 U643 ( .A(n560), .B(KEYINPUT30), .ZN(n565) );
  INV_X1 U644 ( .A(G900), .ZN(n562) );
  NAND2_X1 U645 ( .A1(n562), .A2(n348), .ZN(n563) );
  AND2_X1 U646 ( .A1(n564), .A2(n563), .ZN(n575) );
  NOR2_X1 U647 ( .A1(n565), .A2(n575), .ZN(n566) );
  NAND2_X1 U648 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X2 U649 ( .A(n568), .B(KEYINPUT73), .ZN(n585) );
  BUF_X1 U650 ( .A(n569), .Z(n599) );
  XNOR2_X1 U651 ( .A(n599), .B(KEYINPUT38), .ZN(n705) );
  INV_X1 U652 ( .A(n666), .ZN(n679) );
  NAND2_X1 U653 ( .A1(n607), .A2(n679), .ZN(n572) );
  XOR2_X1 U654 ( .A(KEYINPUT112), .B(KEYINPUT40), .Z(n571) );
  NOR2_X1 U655 ( .A1(n709), .A2(n381), .ZN(n573) );
  NAND2_X1 U656 ( .A1(n573), .A2(n705), .ZN(n574) );
  XNOR2_X1 U657 ( .A(n574), .B(KEYINPUT41), .ZN(n699) );
  NOR2_X1 U658 ( .A1(n575), .A2(n686), .ZN(n576) );
  NAND2_X1 U659 ( .A1(n577), .A2(n576), .ZN(n598) );
  NOR2_X1 U660 ( .A1(n578), .A2(n598), .ZN(n579) );
  XNOR2_X1 U661 ( .A(n579), .B(KEYINPUT28), .ZN(n582) );
  INV_X1 U662 ( .A(KEYINPUT111), .ZN(n580) );
  AND2_X1 U663 ( .A1(n582), .A2(n581), .ZN(n591) );
  NAND2_X1 U664 ( .A1(n699), .A2(n591), .ZN(n583) );
  XOR2_X1 U665 ( .A(n583), .B(KEYINPUT42), .Z(n750) );
  NOR2_X1 U666 ( .A1(n652), .A2(n750), .ZN(n584) );
  INV_X1 U667 ( .A(n585), .ZN(n588) );
  NAND2_X1 U668 ( .A1(n586), .A2(n378), .ZN(n587) );
  XNOR2_X1 U669 ( .A(n631), .B(n589), .ZN(n593) );
  AND2_X1 U670 ( .A1(n590), .A2(n591), .ZN(n680) );
  NAND2_X1 U671 ( .A1(n680), .A2(n701), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n603), .A2(KEYINPUT47), .ZN(n592) );
  NAND2_X1 U673 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U674 ( .A(n594), .B(KEYINPUT79), .ZN(n606) );
  AND2_X1 U675 ( .A1(n595), .A2(n679), .ZN(n596) );
  NAND2_X1 U676 ( .A1(n596), .A2(n706), .ZN(n597) );
  OR2_X1 U677 ( .A1(n598), .A2(n597), .ZN(n609) );
  NOR2_X1 U678 ( .A1(n609), .A2(n599), .ZN(n600) );
  XOR2_X1 U679 ( .A(n600), .B(KEYINPUT36), .Z(n602) );
  NOR2_X1 U680 ( .A1(n602), .A2(n601), .ZN(n683) );
  NOR2_X1 U681 ( .A1(n603), .A2(KEYINPUT47), .ZN(n604) );
  NOR2_X1 U682 ( .A1(n683), .A2(n604), .ZN(n605) );
  INV_X1 U683 ( .A(n607), .ZN(n608) );
  NOR2_X1 U684 ( .A1(n608), .A2(n675), .ZN(n638) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT108), .ZN(n610) );
  NOR2_X1 U686 ( .A1(n610), .A2(n689), .ZN(n612) );
  XOR2_X1 U687 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n611) );
  XNOR2_X1 U688 ( .A(n612), .B(n611), .ZN(n613) );
  NOR2_X1 U689 ( .A1(n613), .A2(n378), .ZN(n636) );
  NOR2_X1 U690 ( .A1(n638), .A2(n636), .ZN(n614) );
  INV_X1 U691 ( .A(n618), .ZN(n619) );
  INV_X1 U692 ( .A(n620), .ZN(n621) );
  NAND2_X1 U693 ( .A1(n621), .A2(KEYINPUT2), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n656), .A2(G478), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(n624), .ZN(n628) );
  INV_X1 U696 ( .A(G952), .ZN(n626) );
  NAND2_X1 U697 ( .A1(n626), .A2(G953), .ZN(n627) );
  XNOR2_X1 U698 ( .A(n627), .B(KEYINPUT90), .ZN(n644) );
  INV_X1 U699 ( .A(n644), .ZN(n662) );
  AND2_X1 U700 ( .A1(n628), .A2(n644), .ZN(G63) );
  NOR2_X1 U701 ( .A1(n632), .A2(n675), .ZN(n630) );
  XNOR2_X1 U702 ( .A(G116), .B(KEYINPUT119), .ZN(n629) );
  XNOR2_X1 U703 ( .A(n630), .B(n629), .ZN(G18) );
  XOR2_X1 U704 ( .A(G143), .B(n631), .Z(G45) );
  NOR2_X1 U705 ( .A1(n632), .A2(n666), .ZN(n633) );
  XOR2_X1 U706 ( .A(G113), .B(n633), .Z(G15) );
  XNOR2_X1 U707 ( .A(n634), .B(G119), .ZN(G21) );
  XNOR2_X1 U708 ( .A(n636), .B(n635), .ZN(G42) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(G36) );
  XOR2_X1 U710 ( .A(n551), .B(G122), .Z(G24) );
  XNOR2_X1 U711 ( .A(KEYINPUT89), .B(KEYINPUT113), .ZN(n639) );
  XNOR2_X1 U712 ( .A(n639), .B(KEYINPUT62), .ZN(n640) );
  XNOR2_X1 U713 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n643), .B(n642), .ZN(n645) );
  NAND2_X1 U715 ( .A1(n645), .A2(n644), .ZN(n647) );
  XOR2_X1 U716 ( .A(KEYINPUT87), .B(KEYINPUT63), .Z(n646) );
  XNOR2_X1 U717 ( .A(n647), .B(n646), .ZN(G57) );
  XNOR2_X1 U718 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n648) );
  XNOR2_X1 U719 ( .A(KEYINPUT124), .B(KEYINPUT59), .ZN(n650) );
  XOR2_X1 U720 ( .A(n652), .B(G131), .Z(G33) );
  NAND2_X1 U721 ( .A1(n656), .A2(G217), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n654), .B(n653), .ZN(n655) );
  NOR2_X1 U723 ( .A1(n655), .A2(n662), .ZN(G66) );
  NAND2_X1 U724 ( .A1(n656), .A2(G469), .ZN(n661) );
  XNOR2_X1 U725 ( .A(KEYINPUT123), .B(KEYINPUT57), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT58), .ZN(n659) );
  XNOR2_X1 U727 ( .A(n657), .B(n659), .ZN(n660) );
  XNOR2_X1 U728 ( .A(n661), .B(n660), .ZN(n663) );
  NOR2_X1 U729 ( .A1(n663), .A2(n662), .ZN(G54) );
  XNOR2_X1 U730 ( .A(n664), .B(G101), .ZN(n665) );
  XNOR2_X1 U731 ( .A(KEYINPUT114), .B(n665), .ZN(G3) );
  NOR2_X1 U732 ( .A1(n666), .A2(n669), .ZN(n668) );
  XNOR2_X1 U733 ( .A(G104), .B(KEYINPUT115), .ZN(n667) );
  XNOR2_X1 U734 ( .A(n668), .B(n667), .ZN(G6) );
  NOR2_X1 U735 ( .A1(n675), .A2(n669), .ZN(n674) );
  XOR2_X1 U736 ( .A(KEYINPUT27), .B(KEYINPUT117), .Z(n671) );
  XNOR2_X1 U737 ( .A(G107), .B(KEYINPUT26), .ZN(n670) );
  XNOR2_X1 U738 ( .A(n671), .B(n670), .ZN(n672) );
  XNOR2_X1 U739 ( .A(KEYINPUT116), .B(n672), .ZN(n673) );
  XNOR2_X1 U740 ( .A(n674), .B(n673), .ZN(G9) );
  XOR2_X1 U741 ( .A(G128), .B(KEYINPUT29), .Z(n678) );
  INV_X1 U742 ( .A(n675), .ZN(n676) );
  NAND2_X1 U743 ( .A1(n680), .A2(n676), .ZN(n677) );
  XNOR2_X1 U744 ( .A(n678), .B(n677), .ZN(G30) );
  NAND2_X1 U745 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U746 ( .A(n681), .B(KEYINPUT118), .ZN(n682) );
  XNOR2_X1 U747 ( .A(G146), .B(n682), .ZN(G48) );
  XNOR2_X1 U748 ( .A(n683), .B(G125), .ZN(n684) );
  XNOR2_X1 U749 ( .A(n684), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U750 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n726) );
  NOR2_X1 U751 ( .A1(n685), .A2(G953), .ZN(n724) );
  NAND2_X1 U752 ( .A1(n687), .A2(n686), .ZN(n688) );
  XOR2_X1 U753 ( .A(KEYINPUT49), .B(n688), .Z(n695) );
  NOR2_X1 U754 ( .A1(n689), .A2(n529), .ZN(n691) );
  XNOR2_X1 U755 ( .A(KEYINPUT50), .B(KEYINPUT120), .ZN(n690) );
  XNOR2_X1 U756 ( .A(n691), .B(n690), .ZN(n693) );
  NOR2_X1 U757 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U758 ( .A1(n695), .A2(n694), .ZN(n697) );
  NAND2_X1 U759 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U760 ( .A(n698), .B(KEYINPUT51), .ZN(n700) );
  INV_X1 U761 ( .A(n699), .ZN(n719) );
  NOR2_X1 U762 ( .A1(n700), .A2(n719), .ZN(n715) );
  NOR2_X1 U763 ( .A1(KEYINPUT121), .A2(n709), .ZN(n703) );
  AND2_X1 U764 ( .A1(n701), .A2(n705), .ZN(n702) );
  NOR2_X1 U765 ( .A1(n703), .A2(n702), .ZN(n704) );
  NOR2_X1 U766 ( .A1(n381), .A2(n704), .ZN(n711) );
  XOR2_X1 U767 ( .A(KEYINPUT121), .B(n705), .Z(n707) );
  NAND2_X1 U768 ( .A1(n707), .A2(n381), .ZN(n708) );
  NOR2_X1 U769 ( .A1(n709), .A2(n708), .ZN(n710) );
  NOR2_X1 U770 ( .A1(n711), .A2(n710), .ZN(n713) );
  BUF_X1 U771 ( .A(n712), .Z(n720) );
  NOR2_X1 U772 ( .A1(n713), .A2(n720), .ZN(n714) );
  NOR2_X1 U773 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U774 ( .A(n716), .B(KEYINPUT52), .ZN(n717) );
  NOR2_X1 U775 ( .A1(n718), .A2(n717), .ZN(n722) );
  NOR2_X1 U776 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U777 ( .A1(n722), .A2(n721), .ZN(n723) );
  NAND2_X1 U778 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U779 ( .A(n726), .B(n725), .ZN(G75) );
  NAND2_X1 U780 ( .A1(n616), .A2(n744), .ZN(n731) );
  NAND2_X1 U781 ( .A1(G953), .A2(G224), .ZN(n728) );
  XNOR2_X1 U782 ( .A(KEYINPUT61), .B(n728), .ZN(n729) );
  NAND2_X1 U783 ( .A1(n729), .A2(G898), .ZN(n730) );
  NAND2_X1 U784 ( .A1(n731), .A2(n730), .ZN(n737) );
  XNOR2_X1 U785 ( .A(n732), .B(G110), .ZN(n733) );
  XNOR2_X1 U786 ( .A(n733), .B(KEYINPUT125), .ZN(n735) );
  NAND2_X1 U787 ( .A1(n735), .A2(n734), .ZN(n736) );
  XOR2_X1 U788 ( .A(n737), .B(n736), .Z(G69) );
  XOR2_X1 U789 ( .A(n739), .B(n738), .Z(n742) );
  XNOR2_X1 U790 ( .A(n740), .B(n742), .ZN(n741) );
  NOR2_X1 U791 ( .A1(n741), .A2(G953), .ZN(n747) );
  XNOR2_X1 U792 ( .A(n742), .B(G227), .ZN(n743) );
  NAND2_X1 U793 ( .A1(n743), .A2(G900), .ZN(n745) );
  NOR2_X1 U794 ( .A1(n745), .A2(n744), .ZN(n746) );
  NOR2_X1 U795 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U796 ( .A(KEYINPUT126), .B(n748), .ZN(G72) );
  XNOR2_X1 U797 ( .A(G110), .B(n749), .ZN(G12) );
  XOR2_X1 U798 ( .A(G137), .B(n750), .Z(G39) );
endmodule

