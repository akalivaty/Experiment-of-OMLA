

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XNOR2_X1 U558 ( .A(n552), .B(n551), .ZN(n554) );
  XNOR2_X1 U559 ( .A(n550), .B(KEYINPUT64), .ZN(n551) );
  AND2_X1 U560 ( .A1(n557), .A2(n556), .ZN(G160) );
  AND2_X1 U561 ( .A1(n811), .A2(n801), .ZN(n524) );
  INV_X1 U562 ( .A(KEYINPUT101), .ZN(n721) );
  INV_X1 U563 ( .A(n732), .ZN(n694) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n716) );
  INV_X1 U565 ( .A(KEYINPUT31), .ZN(n728) );
  XNOR2_X1 U566 ( .A(n717), .B(n716), .ZN(n718) );
  INV_X1 U567 ( .A(n982), .ZN(n752) );
  AND2_X1 U568 ( .A1(n754), .A2(n753), .ZN(n755) );
  OR2_X1 U569 ( .A1(n769), .A2(n686), .ZN(n732) );
  INV_X1 U570 ( .A(KEYINPUT23), .ZN(n550) );
  NOR2_X1 U571 ( .A1(G2104), .A2(n542), .ZN(n878) );
  NAND2_X1 U572 ( .A1(n524), .A2(n802), .ZN(n803) );
  AND2_X1 U573 ( .A1(n542), .A2(G2104), .ZN(n874) );
  OR2_X1 U574 ( .A1(n804), .A2(n803), .ZN(n819) );
  NOR2_X1 U575 ( .A1(G651), .A2(n633), .ZN(n648) );
  NOR2_X1 U576 ( .A1(G651), .A2(G543), .ZN(n652) );
  NAND2_X1 U577 ( .A1(G89), .A2(n652), .ZN(n525) );
  XNOR2_X1 U578 ( .A(n525), .B(KEYINPUT76), .ZN(n526) );
  XNOR2_X1 U579 ( .A(n526), .B(KEYINPUT4), .ZN(n528) );
  XOR2_X1 U580 ( .A(KEYINPUT0), .B(G543), .Z(n633) );
  INV_X1 U581 ( .A(G651), .ZN(n530) );
  NOR2_X1 U582 ( .A1(n633), .A2(n530), .ZN(n651) );
  NAND2_X1 U583 ( .A1(G76), .A2(n651), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U585 ( .A(n529), .B(KEYINPUT5), .ZN(n536) );
  NOR2_X1 U586 ( .A1(G543), .A2(n530), .ZN(n531) );
  XOR2_X1 U587 ( .A(KEYINPUT1), .B(n531), .Z(n647) );
  NAND2_X1 U588 ( .A1(G63), .A2(n647), .ZN(n533) );
  NAND2_X1 U589 ( .A1(G51), .A2(n648), .ZN(n532) );
  NAND2_X1 U590 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U591 ( .A(KEYINPUT6), .B(n534), .Z(n535) );
  NAND2_X1 U592 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U593 ( .A(n537), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U594 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U595 ( .A(G2105), .ZN(n542) );
  NAND2_X1 U596 ( .A1(n878), .A2(G126), .ZN(n538) );
  XNOR2_X1 U597 ( .A(n538), .B(KEYINPUT90), .ZN(n541) );
  NOR2_X1 U598 ( .A1(G2105), .A2(G2104), .ZN(n539) );
  XOR2_X1 U599 ( .A(KEYINPUT17), .B(n539), .Z(n873) );
  NAND2_X1 U600 ( .A1(G138), .A2(n873), .ZN(n540) );
  NAND2_X1 U601 ( .A1(n541), .A2(n540), .ZN(n547) );
  NAND2_X1 U602 ( .A1(G102), .A2(n874), .ZN(n545) );
  NAND2_X1 U603 ( .A1(G2104), .A2(G2105), .ZN(n543) );
  XOR2_X1 U604 ( .A(KEYINPUT66), .B(n543), .Z(n877) );
  NAND2_X1 U605 ( .A1(G114), .A2(n877), .ZN(n544) );
  NAND2_X1 U606 ( .A1(n545), .A2(n544), .ZN(n546) );
  NOR2_X1 U607 ( .A1(n547), .A2(n546), .ZN(G164) );
  NAND2_X1 U608 ( .A1(G137), .A2(n873), .ZN(n549) );
  NAND2_X1 U609 ( .A1(G113), .A2(n877), .ZN(n548) );
  AND2_X1 U610 ( .A1(n549), .A2(n548), .ZN(n557) );
  NAND2_X1 U611 ( .A1(G101), .A2(n874), .ZN(n552) );
  NAND2_X1 U612 ( .A1(G125), .A2(n878), .ZN(n553) );
  NAND2_X1 U613 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U614 ( .A(KEYINPUT65), .B(n555), .ZN(n556) );
  AND2_X1 U615 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U616 ( .A(G132), .ZN(G219) );
  INV_X1 U617 ( .A(G82), .ZN(G220) );
  INV_X1 U618 ( .A(G108), .ZN(G238) );
  XOR2_X1 U619 ( .A(KEYINPUT73), .B(KEYINPUT11), .Z(n561) );
  XOR2_X1 U620 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n559) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n558) );
  XOR2_X1 U622 ( .A(n559), .B(n558), .Z(n922) );
  NAND2_X1 U623 ( .A1(G567), .A2(n922), .ZN(n560) );
  XNOR2_X1 U624 ( .A(n561), .B(n560), .ZN(n562) );
  XOR2_X1 U625 ( .A(KEYINPUT72), .B(n562), .Z(G234) );
  XOR2_X1 U626 ( .A(KEYINPUT14), .B(KEYINPUT74), .Z(n564) );
  NAND2_X1 U627 ( .A1(G56), .A2(n647), .ZN(n563) );
  XNOR2_X1 U628 ( .A(n564), .B(n563), .ZN(n572) );
  NAND2_X1 U629 ( .A1(n652), .A2(G81), .ZN(n565) );
  XNOR2_X1 U630 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U631 ( .A1(G68), .A2(n651), .ZN(n566) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U634 ( .A1(G43), .A2(n648), .ZN(n569) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n571) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n904) );
  NAND2_X1 U637 ( .A1(n904), .A2(G860), .ZN(G153) );
  NAND2_X1 U638 ( .A1(G64), .A2(n647), .ZN(n574) );
  NAND2_X1 U639 ( .A1(G52), .A2(n648), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n579) );
  NAND2_X1 U641 ( .A1(G77), .A2(n651), .ZN(n576) );
  NAND2_X1 U642 ( .A1(G90), .A2(n652), .ZN(n575) );
  NAND2_X1 U643 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U644 ( .A(KEYINPUT9), .B(n577), .Z(n578) );
  NOR2_X1 U645 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U646 ( .A(KEYINPUT69), .B(n580), .ZN(G301) );
  NAND2_X1 U647 ( .A1(G868), .A2(G301), .ZN(n590) );
  NAND2_X1 U648 ( .A1(G66), .A2(n647), .ZN(n582) );
  NAND2_X1 U649 ( .A1(G92), .A2(n652), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(n587) );
  NAND2_X1 U651 ( .A1(G79), .A2(n651), .ZN(n584) );
  NAND2_X1 U652 ( .A1(G54), .A2(n648), .ZN(n583) );
  NAND2_X1 U653 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U654 ( .A(KEYINPUT75), .B(n585), .Z(n586) );
  NOR2_X1 U655 ( .A1(n587), .A2(n586), .ZN(n588) );
  XOR2_X1 U656 ( .A(KEYINPUT15), .B(n588), .Z(n973) );
  INV_X1 U657 ( .A(n973), .ZN(n703) );
  INV_X1 U658 ( .A(G868), .ZN(n667) );
  NAND2_X1 U659 ( .A1(n703), .A2(n667), .ZN(n589) );
  NAND2_X1 U660 ( .A1(n590), .A2(n589), .ZN(G284) );
  NAND2_X1 U661 ( .A1(G65), .A2(n647), .ZN(n592) );
  NAND2_X1 U662 ( .A1(G91), .A2(n652), .ZN(n591) );
  NAND2_X1 U663 ( .A1(n592), .A2(n591), .ZN(n595) );
  NAND2_X1 U664 ( .A1(n651), .A2(G78), .ZN(n593) );
  XOR2_X1 U665 ( .A(KEYINPUT70), .B(n593), .Z(n594) );
  NOR2_X1 U666 ( .A1(n595), .A2(n594), .ZN(n597) );
  NAND2_X1 U667 ( .A1(n648), .A2(G53), .ZN(n596) );
  NAND2_X1 U668 ( .A1(n597), .A2(n596), .ZN(G299) );
  NOR2_X1 U669 ( .A1(G286), .A2(n667), .ZN(n599) );
  NOR2_X1 U670 ( .A1(G868), .A2(G299), .ZN(n598) );
  NOR2_X1 U671 ( .A1(n599), .A2(n598), .ZN(G297) );
  INV_X1 U672 ( .A(G860), .ZN(n600) );
  NAND2_X1 U673 ( .A1(n600), .A2(G559), .ZN(n601) );
  NAND2_X1 U674 ( .A1(n601), .A2(n973), .ZN(n602) );
  XNOR2_X1 U675 ( .A(n602), .B(KEYINPUT77), .ZN(n603) );
  XOR2_X1 U676 ( .A(KEYINPUT16), .B(n603), .Z(G148) );
  INV_X1 U677 ( .A(n904), .ZN(n980) );
  NOR2_X1 U678 ( .A1(G868), .A2(n980), .ZN(n606) );
  NAND2_X1 U679 ( .A1(n973), .A2(G868), .ZN(n604) );
  NOR2_X1 U680 ( .A1(G559), .A2(n604), .ZN(n605) );
  NOR2_X1 U681 ( .A1(n606), .A2(n605), .ZN(G282) );
  XOR2_X1 U682 ( .A(KEYINPUT18), .B(KEYINPUT79), .Z(n608) );
  NAND2_X1 U683 ( .A1(G123), .A2(n878), .ZN(n607) );
  XNOR2_X1 U684 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U685 ( .A(n609), .B(KEYINPUT78), .ZN(n611) );
  NAND2_X1 U686 ( .A1(n874), .A2(G99), .ZN(n610) );
  NAND2_X1 U687 ( .A1(n611), .A2(n610), .ZN(n615) );
  NAND2_X1 U688 ( .A1(G135), .A2(n873), .ZN(n613) );
  NAND2_X1 U689 ( .A1(G111), .A2(n877), .ZN(n612) );
  NAND2_X1 U690 ( .A1(n613), .A2(n612), .ZN(n614) );
  NOR2_X1 U691 ( .A1(n615), .A2(n614), .ZN(n939) );
  XNOR2_X1 U692 ( .A(n939), .B(G2096), .ZN(n616) );
  INV_X1 U693 ( .A(G2100), .ZN(n836) );
  NAND2_X1 U694 ( .A1(n616), .A2(n836), .ZN(G156) );
  NAND2_X1 U695 ( .A1(n652), .A2(G85), .ZN(n623) );
  NAND2_X1 U696 ( .A1(G60), .A2(n647), .ZN(n618) );
  NAND2_X1 U697 ( .A1(G47), .A2(n648), .ZN(n617) );
  NAND2_X1 U698 ( .A1(n618), .A2(n617), .ZN(n621) );
  NAND2_X1 U699 ( .A1(G72), .A2(n651), .ZN(n619) );
  XNOR2_X1 U700 ( .A(KEYINPUT67), .B(n619), .ZN(n620) );
  NOR2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U702 ( .A1(n623), .A2(n622), .ZN(n624) );
  XNOR2_X1 U703 ( .A(n624), .B(KEYINPUT68), .ZN(G290) );
  NAND2_X1 U704 ( .A1(G73), .A2(n651), .ZN(n625) );
  XOR2_X1 U705 ( .A(KEYINPUT2), .B(n625), .Z(n630) );
  NAND2_X1 U706 ( .A1(G61), .A2(n647), .ZN(n627) );
  NAND2_X1 U707 ( .A1(G86), .A2(n652), .ZN(n626) );
  NAND2_X1 U708 ( .A1(n627), .A2(n626), .ZN(n628) );
  XOR2_X1 U709 ( .A(KEYINPUT83), .B(n628), .Z(n629) );
  NOR2_X1 U710 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U711 ( .A1(n648), .A2(G48), .ZN(n631) );
  NAND2_X1 U712 ( .A1(n632), .A2(n631), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G49), .A2(n648), .ZN(n635) );
  NAND2_X1 U714 ( .A1(G87), .A2(n633), .ZN(n634) );
  NAND2_X1 U715 ( .A1(n635), .A2(n634), .ZN(n636) );
  NOR2_X1 U716 ( .A1(n647), .A2(n636), .ZN(n638) );
  NAND2_X1 U717 ( .A1(G651), .A2(G74), .ZN(n637) );
  NAND2_X1 U718 ( .A1(n638), .A2(n637), .ZN(G288) );
  NAND2_X1 U719 ( .A1(G62), .A2(n647), .ZN(n640) );
  NAND2_X1 U720 ( .A1(G50), .A2(n648), .ZN(n639) );
  NAND2_X1 U721 ( .A1(n640), .A2(n639), .ZN(n641) );
  XOR2_X1 U722 ( .A(KEYINPUT84), .B(n641), .Z(n645) );
  NAND2_X1 U723 ( .A1(n651), .A2(G75), .ZN(n643) );
  NAND2_X1 U724 ( .A1(G88), .A2(n652), .ZN(n642) );
  AND2_X1 U725 ( .A1(n643), .A2(n642), .ZN(n644) );
  NAND2_X1 U726 ( .A1(n645), .A2(n644), .ZN(G303) );
  INV_X1 U727 ( .A(G303), .ZN(G166) );
  NAND2_X1 U728 ( .A1(G559), .A2(n973), .ZN(n646) );
  XOR2_X1 U729 ( .A(n646), .B(n980), .Z(n915) );
  NAND2_X1 U730 ( .A1(G67), .A2(n647), .ZN(n650) );
  NAND2_X1 U731 ( .A1(G55), .A2(n648), .ZN(n649) );
  NAND2_X1 U732 ( .A1(n650), .A2(n649), .ZN(n657) );
  NAND2_X1 U733 ( .A1(G80), .A2(n651), .ZN(n654) );
  NAND2_X1 U734 ( .A1(G93), .A2(n652), .ZN(n653) );
  NAND2_X1 U735 ( .A1(n654), .A2(n653), .ZN(n655) );
  XOR2_X1 U736 ( .A(KEYINPUT81), .B(n655), .Z(n656) );
  NOR2_X1 U737 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U738 ( .A(KEYINPUT82), .B(n658), .Z(n918) );
  XNOR2_X1 U739 ( .A(G290), .B(n918), .ZN(n664) );
  XOR2_X1 U740 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n659) );
  XNOR2_X1 U741 ( .A(G288), .B(n659), .ZN(n660) );
  XNOR2_X1 U742 ( .A(G305), .B(n660), .ZN(n662) );
  XOR2_X1 U743 ( .A(G299), .B(G166), .Z(n661) );
  XNOR2_X1 U744 ( .A(n662), .B(n661), .ZN(n663) );
  XNOR2_X1 U745 ( .A(n664), .B(n663), .ZN(n903) );
  XNOR2_X1 U746 ( .A(n915), .B(n903), .ZN(n665) );
  XNOR2_X1 U747 ( .A(KEYINPUT86), .B(n665), .ZN(n666) );
  NOR2_X1 U748 ( .A1(n667), .A2(n666), .ZN(n669) );
  NOR2_X1 U749 ( .A1(n918), .A2(G868), .ZN(n668) );
  NOR2_X1 U750 ( .A1(n669), .A2(n668), .ZN(G295) );
  NAND2_X1 U751 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U752 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U753 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U754 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U755 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U756 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U757 ( .A1(G69), .A2(G120), .ZN(n674) );
  XOR2_X1 U758 ( .A(KEYINPUT87), .B(n674), .Z(n675) );
  NOR2_X1 U759 ( .A1(G238), .A2(n675), .ZN(n676) );
  NAND2_X1 U760 ( .A1(G57), .A2(n676), .ZN(n919) );
  NAND2_X1 U761 ( .A1(n919), .A2(G567), .ZN(n681) );
  NOR2_X1 U762 ( .A1(G220), .A2(G219), .ZN(n677) );
  XOR2_X1 U763 ( .A(KEYINPUT22), .B(n677), .Z(n678) );
  NOR2_X1 U764 ( .A1(G218), .A2(n678), .ZN(n679) );
  NAND2_X1 U765 ( .A1(G96), .A2(n679), .ZN(n920) );
  NAND2_X1 U766 ( .A1(n920), .A2(G2106), .ZN(n680) );
  NAND2_X1 U767 ( .A1(n681), .A2(n680), .ZN(n921) );
  NAND2_X1 U768 ( .A1(G661), .A2(G483), .ZN(n682) );
  XNOR2_X1 U769 ( .A(KEYINPUT88), .B(n682), .ZN(n683) );
  NOR2_X1 U770 ( .A1(n921), .A2(n683), .ZN(n825) );
  NAND2_X1 U771 ( .A1(n825), .A2(G36), .ZN(n684) );
  XOR2_X1 U772 ( .A(KEYINPUT89), .B(n684), .Z(G176) );
  INV_X1 U773 ( .A(G301), .ZN(G171) );
  NAND2_X1 U774 ( .A1(G160), .A2(G40), .ZN(n769) );
  NOR2_X1 U775 ( .A1(G164), .A2(G1384), .ZN(n770) );
  INV_X1 U776 ( .A(n770), .ZN(n686) );
  NAND2_X1 U777 ( .A1(G8), .A2(n732), .ZN(n763) );
  NOR2_X1 U778 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U779 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  NOR2_X1 U780 ( .A1(n763), .A2(n688), .ZN(n768) );
  XNOR2_X1 U781 ( .A(G2078), .B(KEYINPUT25), .ZN(n958) );
  NOR2_X1 U782 ( .A1(n732), .A2(n958), .ZN(n690) );
  INV_X1 U783 ( .A(G1961), .ZN(n1010) );
  NOR2_X1 U784 ( .A1(n694), .A2(n1010), .ZN(n689) );
  NOR2_X1 U785 ( .A1(n690), .A2(n689), .ZN(n720) );
  NAND2_X1 U786 ( .A1(G171), .A2(n720), .ZN(n719) );
  INV_X1 U787 ( .A(G299), .ZN(n984) );
  NAND2_X1 U788 ( .A1(n694), .A2(G2072), .ZN(n691) );
  XNOR2_X1 U789 ( .A(n691), .B(KEYINPUT27), .ZN(n693) );
  XOR2_X1 U790 ( .A(G1956), .B(KEYINPUT98), .Z(n1000) );
  NOR2_X1 U791 ( .A1(n694), .A2(n1000), .ZN(n692) );
  NOR2_X1 U792 ( .A1(n693), .A2(n692), .ZN(n712) );
  NAND2_X1 U793 ( .A1(n984), .A2(n712), .ZN(n711) );
  NAND2_X1 U794 ( .A1(G1996), .A2(n694), .ZN(n695) );
  XNOR2_X1 U795 ( .A(n695), .B(KEYINPUT26), .ZN(n697) );
  NAND2_X1 U796 ( .A1(G1341), .A2(n732), .ZN(n696) );
  NAND2_X1 U797 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U798 ( .A(KEYINPUT99), .B(n698), .ZN(n704) );
  NAND2_X1 U799 ( .A1(n904), .A2(n704), .ZN(n699) );
  NAND2_X1 U800 ( .A1(n699), .A2(n703), .ZN(n709) );
  INV_X1 U801 ( .A(G2067), .ZN(n840) );
  NOR2_X1 U802 ( .A1(n732), .A2(n840), .ZN(n700) );
  XOR2_X1 U803 ( .A(n700), .B(KEYINPUT100), .Z(n702) );
  NAND2_X1 U804 ( .A1(n732), .A2(G1348), .ZN(n701) );
  NAND2_X1 U805 ( .A1(n702), .A2(n701), .ZN(n707) );
  NOR2_X1 U806 ( .A1(n703), .A2(n980), .ZN(n705) );
  NAND2_X1 U807 ( .A1(n705), .A2(n704), .ZN(n706) );
  NAND2_X1 U808 ( .A1(n707), .A2(n706), .ZN(n708) );
  NAND2_X1 U809 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U810 ( .A1(n711), .A2(n710), .ZN(n715) );
  NOR2_X1 U811 ( .A1(n984), .A2(n712), .ZN(n713) );
  XOR2_X1 U812 ( .A(n713), .B(KEYINPUT28), .Z(n714) );
  NAND2_X1 U813 ( .A1(n715), .A2(n714), .ZN(n717) );
  NAND2_X1 U814 ( .A1(n719), .A2(n718), .ZN(n731) );
  NOR2_X1 U815 ( .A1(G171), .A2(n720), .ZN(n727) );
  NOR2_X1 U816 ( .A1(G1966), .A2(n763), .ZN(n744) );
  NOR2_X1 U817 ( .A1(G2084), .A2(n732), .ZN(n740) );
  NOR2_X1 U818 ( .A1(n744), .A2(n740), .ZN(n722) );
  XNOR2_X1 U819 ( .A(n722), .B(n721), .ZN(n723) );
  NAND2_X1 U820 ( .A1(n723), .A2(G8), .ZN(n724) );
  XNOR2_X1 U821 ( .A(KEYINPUT30), .B(n724), .ZN(n725) );
  NOR2_X1 U822 ( .A1(G168), .A2(n725), .ZN(n726) );
  NOR2_X1 U823 ( .A1(n727), .A2(n726), .ZN(n729) );
  XNOR2_X1 U824 ( .A(n729), .B(n728), .ZN(n730) );
  NAND2_X1 U825 ( .A1(n731), .A2(n730), .ZN(n742) );
  NAND2_X1 U826 ( .A1(n742), .A2(G286), .ZN(n737) );
  NOR2_X1 U827 ( .A1(G1971), .A2(n763), .ZN(n734) );
  NOR2_X1 U828 ( .A1(G2090), .A2(n732), .ZN(n733) );
  NOR2_X1 U829 ( .A1(n734), .A2(n733), .ZN(n735) );
  NAND2_X1 U830 ( .A1(n735), .A2(G303), .ZN(n736) );
  NAND2_X1 U831 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U832 ( .A1(G8), .A2(n738), .ZN(n739) );
  XNOR2_X1 U833 ( .A(n739), .B(KEYINPUT32), .ZN(n748) );
  NAND2_X1 U834 ( .A1(G8), .A2(n740), .ZN(n741) );
  XOR2_X1 U835 ( .A(KEYINPUT97), .B(n741), .Z(n746) );
  INV_X1 U836 ( .A(n742), .ZN(n743) );
  NOR2_X1 U837 ( .A1(n744), .A2(n743), .ZN(n745) );
  NAND2_X1 U838 ( .A1(n746), .A2(n745), .ZN(n747) );
  NAND2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n762) );
  NOR2_X1 U840 ( .A1(G1976), .A2(G288), .ZN(n981) );
  NOR2_X1 U841 ( .A1(G1971), .A2(G303), .ZN(n749) );
  NOR2_X1 U842 ( .A1(n981), .A2(n749), .ZN(n750) );
  XNOR2_X1 U843 ( .A(n750), .B(KEYINPUT102), .ZN(n751) );
  NAND2_X1 U844 ( .A1(n762), .A2(n751), .ZN(n754) );
  NAND2_X1 U845 ( .A1(G1976), .A2(G288), .ZN(n982) );
  NOR2_X1 U846 ( .A1(n763), .A2(n752), .ZN(n753) );
  NOR2_X1 U847 ( .A1(KEYINPUT33), .A2(n755), .ZN(n758) );
  NAND2_X1 U848 ( .A1(n981), .A2(KEYINPUT33), .ZN(n756) );
  NOR2_X1 U849 ( .A1(n756), .A2(n763), .ZN(n757) );
  NOR2_X1 U850 ( .A1(n758), .A2(n757), .ZN(n759) );
  XOR2_X1 U851 ( .A(G1981), .B(G305), .Z(n976) );
  NAND2_X1 U852 ( .A1(n759), .A2(n976), .ZN(n766) );
  NOR2_X1 U853 ( .A1(G2090), .A2(G303), .ZN(n760) );
  NAND2_X1 U854 ( .A1(G8), .A2(n760), .ZN(n761) );
  NAND2_X1 U855 ( .A1(n762), .A2(n761), .ZN(n764) );
  NAND2_X1 U856 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U857 ( .A1(n766), .A2(n765), .ZN(n767) );
  NOR2_X1 U858 ( .A1(n768), .A2(n767), .ZN(n804) );
  NOR2_X1 U859 ( .A1(n770), .A2(n769), .ZN(n816) );
  NAND2_X1 U860 ( .A1(n873), .A2(G140), .ZN(n771) );
  XOR2_X1 U861 ( .A(KEYINPUT91), .B(n771), .Z(n773) );
  NAND2_X1 U862 ( .A1(n874), .A2(G104), .ZN(n772) );
  NAND2_X1 U863 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U864 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U865 ( .A1(G128), .A2(n878), .ZN(n776) );
  NAND2_X1 U866 ( .A1(G116), .A2(n877), .ZN(n775) );
  NAND2_X1 U867 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U868 ( .A(KEYINPUT35), .B(n777), .Z(n778) );
  NOR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(n780) );
  XNOR2_X1 U870 ( .A(KEYINPUT36), .B(n780), .ZN(n899) );
  XOR2_X1 U871 ( .A(KEYINPUT37), .B(n840), .Z(n813) );
  NOR2_X1 U872 ( .A1(n899), .A2(n813), .ZN(n929) );
  NAND2_X1 U873 ( .A1(n816), .A2(n929), .ZN(n811) );
  NAND2_X1 U874 ( .A1(G105), .A2(n874), .ZN(n781) );
  XOR2_X1 U875 ( .A(KEYINPUT38), .B(n781), .Z(n786) );
  NAND2_X1 U876 ( .A1(G129), .A2(n878), .ZN(n783) );
  NAND2_X1 U877 ( .A1(G117), .A2(n877), .ZN(n782) );
  NAND2_X1 U878 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U879 ( .A(KEYINPUT95), .B(n784), .Z(n785) );
  NOR2_X1 U880 ( .A1(n786), .A2(n785), .ZN(n788) );
  NAND2_X1 U881 ( .A1(n873), .A2(G141), .ZN(n787) );
  NAND2_X1 U882 ( .A1(n788), .A2(n787), .ZN(n890) );
  AND2_X1 U883 ( .A1(n890), .A2(G1996), .ZN(n799) );
  NAND2_X1 U884 ( .A1(n874), .A2(G95), .ZN(n789) );
  XOR2_X1 U885 ( .A(KEYINPUT93), .B(n789), .Z(n791) );
  NAND2_X1 U886 ( .A1(n873), .A2(G131), .ZN(n790) );
  NAND2_X1 U887 ( .A1(n791), .A2(n790), .ZN(n792) );
  XNOR2_X1 U888 ( .A(KEYINPUT94), .B(n792), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n878), .A2(G119), .ZN(n793) );
  XNOR2_X1 U890 ( .A(n793), .B(KEYINPUT92), .ZN(n795) );
  NAND2_X1 U891 ( .A1(G107), .A2(n877), .ZN(n794) );
  NAND2_X1 U892 ( .A1(n795), .A2(n794), .ZN(n796) );
  NOR2_X1 U893 ( .A1(n797), .A2(n796), .ZN(n887) );
  INV_X1 U894 ( .A(G1991), .ZN(n949) );
  NOR2_X1 U895 ( .A1(n887), .A2(n949), .ZN(n798) );
  NOR2_X1 U896 ( .A1(n799), .A2(n798), .ZN(n931) );
  XOR2_X1 U897 ( .A(n816), .B(KEYINPUT96), .Z(n800) );
  NOR2_X1 U898 ( .A1(n931), .A2(n800), .ZN(n808) );
  INV_X1 U899 ( .A(n808), .ZN(n801) );
  XNOR2_X1 U900 ( .A(G1986), .B(G290), .ZN(n990) );
  NAND2_X1 U901 ( .A1(n990), .A2(n816), .ZN(n802) );
  NOR2_X1 U902 ( .A1(G1996), .A2(n890), .ZN(n937) );
  NOR2_X1 U903 ( .A1(G1986), .A2(G290), .ZN(n806) );
  AND2_X1 U904 ( .A1(n949), .A2(n887), .ZN(n805) );
  XOR2_X1 U905 ( .A(KEYINPUT103), .B(n805), .Z(n940) );
  NOR2_X1 U906 ( .A1(n806), .A2(n940), .ZN(n807) );
  NOR2_X1 U907 ( .A1(n808), .A2(n807), .ZN(n809) );
  NOR2_X1 U908 ( .A1(n937), .A2(n809), .ZN(n810) );
  XNOR2_X1 U909 ( .A(n810), .B(KEYINPUT39), .ZN(n812) );
  NAND2_X1 U910 ( .A1(n812), .A2(n811), .ZN(n814) );
  NAND2_X1 U911 ( .A1(n899), .A2(n813), .ZN(n930) );
  NAND2_X1 U912 ( .A1(n814), .A2(n930), .ZN(n815) );
  XNOR2_X1 U913 ( .A(KEYINPUT104), .B(n815), .ZN(n817) );
  NAND2_X1 U914 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U915 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U916 ( .A(KEYINPUT40), .B(n820), .ZN(G329) );
  NAND2_X1 U917 ( .A1(G2106), .A2(n922), .ZN(G217) );
  INV_X1 U918 ( .A(G661), .ZN(n822) );
  NAND2_X1 U919 ( .A1(G2), .A2(G15), .ZN(n821) );
  NOR2_X1 U920 ( .A1(n822), .A2(n821), .ZN(n823) );
  XOR2_X1 U921 ( .A(KEYINPUT106), .B(n823), .Z(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n824) );
  NAND2_X1 U923 ( .A1(n825), .A2(n824), .ZN(G188) );
  XNOR2_X1 U924 ( .A(G120), .B(KEYINPUT107), .ZN(G236) );
  XNOR2_X1 U925 ( .A(G1341), .B(G2454), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n826), .B(G2430), .ZN(n827) );
  XNOR2_X1 U927 ( .A(n827), .B(G1348), .ZN(n833) );
  XOR2_X1 U928 ( .A(G2443), .B(G2427), .Z(n829) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n828) );
  XNOR2_X1 U930 ( .A(n829), .B(n828), .ZN(n831) );
  XOR2_X1 U931 ( .A(G2451), .B(G2435), .Z(n830) );
  XNOR2_X1 U932 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U933 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U934 ( .A1(n834), .A2(G14), .ZN(n835) );
  XNOR2_X1 U935 ( .A(KEYINPUT105), .B(n835), .ZN(G401) );
  XNOR2_X1 U936 ( .A(n836), .B(G2678), .ZN(n838) );
  XNOR2_X1 U937 ( .A(G2090), .B(KEYINPUT43), .ZN(n837) );
  XNOR2_X1 U938 ( .A(n838), .B(n837), .ZN(n839) );
  XOR2_X1 U939 ( .A(n839), .B(KEYINPUT108), .Z(n842) );
  XOR2_X1 U940 ( .A(n840), .B(G2072), .Z(n841) );
  XNOR2_X1 U941 ( .A(n842), .B(n841), .ZN(n846) );
  XOR2_X1 U942 ( .A(KEYINPUT42), .B(G2096), .Z(n844) );
  XNOR2_X1 U943 ( .A(G2078), .B(G2084), .ZN(n843) );
  XNOR2_X1 U944 ( .A(n844), .B(n843), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(G227) );
  XOR2_X1 U946 ( .A(G1971), .B(G1956), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1986), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U949 ( .A(G1976), .B(G1981), .Z(n850) );
  XOR2_X1 U950 ( .A(G1966), .B(n1010), .Z(n849) );
  XNOR2_X1 U951 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U952 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U953 ( .A(G2474), .B(KEYINPUT41), .ZN(n853) );
  XNOR2_X1 U954 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U955 ( .A(KEYINPUT109), .B(n855), .ZN(n856) );
  XOR2_X1 U956 ( .A(n856), .B(G1991), .Z(G229) );
  NAND2_X1 U957 ( .A1(n878), .A2(G124), .ZN(n857) );
  XNOR2_X1 U958 ( .A(n857), .B(KEYINPUT44), .ZN(n859) );
  NAND2_X1 U959 ( .A1(G136), .A2(n873), .ZN(n858) );
  NAND2_X1 U960 ( .A1(n859), .A2(n858), .ZN(n860) );
  XNOR2_X1 U961 ( .A(KEYINPUT110), .B(n860), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G100), .A2(n874), .ZN(n862) );
  NAND2_X1 U963 ( .A1(G112), .A2(n877), .ZN(n861) );
  NAND2_X1 U964 ( .A1(n862), .A2(n861), .ZN(n863) );
  NOR2_X1 U965 ( .A1(n864), .A2(n863), .ZN(G162) );
  NAND2_X1 U966 ( .A1(G142), .A2(n873), .ZN(n866) );
  NAND2_X1 U967 ( .A1(G106), .A2(n874), .ZN(n865) );
  NAND2_X1 U968 ( .A1(n866), .A2(n865), .ZN(n867) );
  XNOR2_X1 U969 ( .A(n867), .B(KEYINPUT45), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G130), .A2(n878), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n872) );
  NAND2_X1 U972 ( .A1(G118), .A2(n877), .ZN(n870) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n870), .ZN(n871) );
  NOR2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n886) );
  NAND2_X1 U975 ( .A1(G139), .A2(n873), .ZN(n876) );
  NAND2_X1 U976 ( .A1(G103), .A2(n874), .ZN(n875) );
  NAND2_X1 U977 ( .A1(n876), .A2(n875), .ZN(n885) );
  XNOR2_X1 U978 ( .A(KEYINPUT47), .B(KEYINPUT114), .ZN(n883) );
  NAND2_X1 U979 ( .A1(G115), .A2(n877), .ZN(n881) );
  NAND2_X1 U980 ( .A1(n878), .A2(G127), .ZN(n879) );
  XOR2_X1 U981 ( .A(KEYINPUT113), .B(n879), .Z(n880) );
  NAND2_X1 U982 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U983 ( .A(n883), .B(n882), .Z(n884) );
  NOR2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n923) );
  XOR2_X1 U985 ( .A(n886), .B(n923), .Z(n889) );
  XNOR2_X1 U986 ( .A(n887), .B(G162), .ZN(n888) );
  XNOR2_X1 U987 ( .A(n889), .B(n888), .ZN(n901) );
  XOR2_X1 U988 ( .A(G160), .B(n890), .Z(n897) );
  XOR2_X1 U989 ( .A(KEYINPUT112), .B(KEYINPUT48), .Z(n892) );
  XNOR2_X1 U990 ( .A(KEYINPUT116), .B(KEYINPUT115), .ZN(n891) );
  XNOR2_X1 U991 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U992 ( .A(n893), .B(KEYINPUT46), .Z(n895) );
  XNOR2_X1 U993 ( .A(G164), .B(n939), .ZN(n894) );
  XNOR2_X1 U994 ( .A(n895), .B(n894), .ZN(n896) );
  XNOR2_X1 U995 ( .A(n897), .B(n896), .ZN(n898) );
  XNOR2_X1 U996 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U998 ( .A1(G37), .A2(n902), .ZN(G395) );
  XNOR2_X1 U999 ( .A(G286), .B(n903), .ZN(n906) );
  XOR2_X1 U1000 ( .A(n973), .B(n904), .Z(n905) );
  XNOR2_X1 U1001 ( .A(n906), .B(n905), .ZN(n908) );
  XNOR2_X1 U1002 ( .A(G301), .B(KEYINPUT117), .ZN(n907) );
  XNOR2_X1 U1003 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1004 ( .A1(G37), .A2(n909), .ZN(G397) );
  OR2_X1 U1005 ( .A1(n921), .A2(G401), .ZN(n912) );
  NOR2_X1 U1006 ( .A1(G227), .A2(G229), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(KEYINPUT49), .B(n910), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(n912), .A2(n911), .ZN(n914) );
  NOR2_X1 U1009 ( .A1(G395), .A2(G397), .ZN(n913) );
  NAND2_X1 U1010 ( .A1(n914), .A2(n913), .ZN(G225) );
  XOR2_X1 U1011 ( .A(KEYINPUT118), .B(G225), .Z(G308) );
  XOR2_X1 U1013 ( .A(n915), .B(KEYINPUT80), .Z(n916) );
  NOR2_X1 U1014 ( .A1(G860), .A2(n916), .ZN(n917) );
  XOR2_X1 U1015 ( .A(n918), .B(n917), .Z(G145) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  INV_X1 U1017 ( .A(G69), .ZN(G235) );
  NOR2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G325) );
  INV_X1 U1019 ( .A(G325), .ZN(G261) );
  INV_X1 U1020 ( .A(n921), .ZN(G319) );
  INV_X1 U1021 ( .A(G57), .ZN(G237) );
  INV_X1 U1022 ( .A(n922), .ZN(G223) );
  XOR2_X1 U1023 ( .A(G2072), .B(n923), .Z(n925) );
  XOR2_X1 U1024 ( .A(G164), .B(G2078), .Z(n924) );
  NOR2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  XOR2_X1 U1026 ( .A(n926), .B(KEYINPUT120), .Z(n927) );
  XNOR2_X1 U1027 ( .A(KEYINPUT50), .B(n927), .ZN(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n935) );
  NAND2_X1 U1029 ( .A1(n931), .A2(n930), .ZN(n933) );
  XOR2_X1 U1030 ( .A(G160), .B(G2084), .Z(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n945) );
  XOR2_X1 U1033 ( .A(G2090), .B(G162), .Z(n936) );
  NOR2_X1 U1034 ( .A1(n937), .A2(n936), .ZN(n938) );
  XOR2_X1 U1035 ( .A(KEYINPUT51), .B(n938), .Z(n943) );
  NOR2_X1 U1036 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1037 ( .A(KEYINPUT119), .B(n941), .Z(n942) );
  NAND2_X1 U1038 ( .A1(n943), .A2(n942), .ZN(n944) );
  NOR2_X1 U1039 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT52), .B(n946), .ZN(n947) );
  INV_X1 U1041 ( .A(KEYINPUT55), .ZN(n969) );
  NAND2_X1 U1042 ( .A1(n947), .A2(n969), .ZN(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(G29), .ZN(n1031) );
  XNOR2_X1 U1044 ( .A(G29), .B(KEYINPUT123), .ZN(n971) );
  XOR2_X1 U1045 ( .A(n949), .B(G25), .Z(n951) );
  XNOR2_X1 U1046 ( .A(G33), .B(G2072), .ZN(n950) );
  NOR2_X1 U1047 ( .A1(n951), .A2(n950), .ZN(n957) );
  XOR2_X1 U1048 ( .A(G32), .B(G1996), .Z(n952) );
  NAND2_X1 U1049 ( .A1(n952), .A2(G28), .ZN(n955) );
  XNOR2_X1 U1050 ( .A(G26), .B(G2067), .ZN(n953) );
  XNOR2_X1 U1051 ( .A(KEYINPUT122), .B(n953), .ZN(n954) );
  NOR2_X1 U1052 ( .A1(n955), .A2(n954), .ZN(n956) );
  NAND2_X1 U1053 ( .A1(n957), .A2(n956), .ZN(n960) );
  XOR2_X1 U1054 ( .A(G27), .B(n958), .Z(n959) );
  NOR2_X1 U1055 ( .A1(n960), .A2(n959), .ZN(n961) );
  XOR2_X1 U1056 ( .A(KEYINPUT53), .B(n961), .Z(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT54), .B(G34), .Z(n962) );
  XNOR2_X1 U1058 ( .A(G2084), .B(n962), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n967) );
  XOR2_X1 U1060 ( .A(KEYINPUT121), .B(G2090), .Z(n965) );
  XNOR2_X1 U1061 ( .A(G35), .B(n965), .ZN(n966) );
  NOR2_X1 U1062 ( .A1(n967), .A2(n966), .ZN(n968) );
  XOR2_X1 U1063 ( .A(n969), .B(n968), .Z(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  NAND2_X1 U1065 ( .A1(G11), .A2(n972), .ZN(n1029) );
  INV_X1 U1066 ( .A(G16), .ZN(n1025) );
  XOR2_X1 U1067 ( .A(n1025), .B(KEYINPUT56), .Z(n999) );
  XOR2_X1 U1068 ( .A(G1348), .B(n973), .Z(n975) );
  XOR2_X1 U1069 ( .A(G301), .B(n1010), .Z(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n997) );
  XNOR2_X1 U1071 ( .A(G1966), .B(G168), .ZN(n977) );
  NAND2_X1 U1072 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1073 ( .A(n978), .B(KEYINPUT57), .ZN(n979) );
  XNOR2_X1 U1074 ( .A(KEYINPUT124), .B(n979), .ZN(n992) );
  XOR2_X1 U1075 ( .A(n980), .B(G1341), .Z(n988) );
  INV_X1 U1076 ( .A(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n986) );
  XOR2_X1 U1078 ( .A(G1956), .B(n984), .Z(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  NAND2_X1 U1080 ( .A1(n988), .A2(n987), .ZN(n989) );
  NOR2_X1 U1081 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1082 ( .A1(n992), .A2(n991), .ZN(n995) );
  XNOR2_X1 U1083 ( .A(G1971), .B(G166), .ZN(n993) );
  XNOR2_X1 U1084 ( .A(KEYINPUT125), .B(n993), .ZN(n994) );
  NOR2_X1 U1085 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1086 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1087 ( .A1(n999), .A2(n998), .ZN(n1027) );
  XNOR2_X1 U1088 ( .A(n1000), .B(G20), .ZN(n1004) );
  XNOR2_X1 U1089 ( .A(G1341), .B(G19), .ZN(n1002) );
  XNOR2_X1 U1090 ( .A(G1981), .B(G6), .ZN(n1001) );
  NOR2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1092 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XOR2_X1 U1093 ( .A(KEYINPUT59), .B(G1348), .Z(n1005) );
  XNOR2_X1 U1094 ( .A(G4), .B(n1005), .ZN(n1006) );
  NOR2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1009) );
  XOR2_X1 U1096 ( .A(KEYINPUT127), .B(KEYINPUT60), .Z(n1008) );
  XNOR2_X1 U1097 ( .A(n1009), .B(n1008), .ZN(n1020) );
  XOR2_X1 U1098 ( .A(n1010), .B(KEYINPUT126), .Z(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(G5), .ZN(n1018) );
  XNOR2_X1 U1100 ( .A(G1971), .B(G22), .ZN(n1013) );
  XNOR2_X1 U1101 ( .A(G23), .B(G1976), .ZN(n1012) );
  NOR2_X1 U1102 ( .A1(n1013), .A2(n1012), .ZN(n1015) );
  XOR2_X1 U1103 ( .A(G1986), .B(G24), .Z(n1014) );
  NAND2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT58), .B(n1016), .ZN(n1017) );
  NOR2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1022) );
  XNOR2_X1 U1108 ( .A(G21), .B(G1966), .ZN(n1021) );
  NOR2_X1 U1109 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1110 ( .A(KEYINPUT61), .B(n1023), .ZN(n1024) );
  NAND2_X1 U1111 ( .A1(n1025), .A2(n1024), .ZN(n1026) );
  NAND2_X1 U1112 ( .A1(n1027), .A2(n1026), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  NAND2_X1 U1114 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XNOR2_X1 U1115 ( .A(KEYINPUT62), .B(n1032), .ZN(G150) );
  INV_X1 U1116 ( .A(G150), .ZN(G311) );
endmodule

