

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897,
         n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908,
         n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919,
         n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, n930,
         n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
         n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n601) );
  BUF_X1 U557 ( .A(n696), .Z(n697) );
  NAND2_X1 U558 ( .A1(G2105), .A2(G2104), .ZN(n521) );
  AND2_X2 U559 ( .A1(n532), .A2(n531), .ZN(G164) );
  INV_X1 U560 ( .A(KEYINPUT105), .ZN(n636) );
  XOR2_X1 U561 ( .A(KEYINPUT68), .B(n521), .Z(n696) );
  XOR2_X1 U562 ( .A(KEYINPUT93), .B(n526), .Z(n520) );
  INV_X1 U563 ( .A(KEYINPUT26), .ZN(n617) );
  NOR2_X1 U564 ( .A1(n973), .A2(n621), .ZN(n638) );
  XNOR2_X1 U565 ( .A(n637), .B(n636), .ZN(n640) );
  INV_X1 U566 ( .A(KEYINPUT64), .ZN(n686) );
  INV_X1 U567 ( .A(KEYINPUT33), .ZN(n688) );
  XOR2_X1 U568 ( .A(KEYINPUT65), .B(n601), .Z(n695) );
  INV_X1 U569 ( .A(KEYINPUT17), .ZN(n528) );
  NAND2_X1 U570 ( .A1(n885), .A2(G138), .ZN(n530) );
  AND2_X1 U571 ( .A1(n527), .A2(n520), .ZN(n532) );
  INV_X1 U572 ( .A(G2104), .ZN(n525) );
  AND2_X1 U573 ( .A1(n525), .A2(G2105), .ZN(n889) );
  NAND2_X1 U574 ( .A1(G126), .A2(n889), .ZN(n523) );
  NAND2_X1 U575 ( .A1(G114), .A2(n696), .ZN(n522) );
  NAND2_X1 U576 ( .A1(n523), .A2(n522), .ZN(n524) );
  XOR2_X1 U577 ( .A(KEYINPUT92), .B(n524), .Z(n527) );
  NOR2_X1 U578 ( .A1(G2105), .A2(n525), .ZN(n702) );
  NAND2_X1 U579 ( .A1(G102), .A2(n702), .ZN(n526) );
  NOR2_X1 U580 ( .A1(G2105), .A2(G2104), .ZN(n529) );
  XNOR2_X2 U581 ( .A(n529), .B(n528), .ZN(n885) );
  XNOR2_X1 U582 ( .A(n530), .B(KEYINPUT94), .ZN(n531) );
  NAND2_X1 U583 ( .A1(G101), .A2(n702), .ZN(n533) );
  XNOR2_X1 U584 ( .A(n533), .B(KEYINPUT67), .ZN(n534) );
  XNOR2_X1 U585 ( .A(KEYINPUT23), .B(n534), .ZN(n537) );
  NAND2_X1 U586 ( .A1(n696), .A2(G113), .ZN(n535) );
  XOR2_X1 U587 ( .A(KEYINPUT69), .B(n535), .Z(n536) );
  AND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n541) );
  NAND2_X1 U589 ( .A1(G125), .A2(n889), .ZN(n539) );
  NAND2_X1 U590 ( .A1(G137), .A2(n885), .ZN(n538) );
  AND2_X1 U591 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U592 ( .A1(n541), .A2(n540), .ZN(G160) );
  INV_X1 U593 ( .A(G651), .ZN(n546) );
  NOR2_X1 U594 ( .A1(G543), .A2(n546), .ZN(n542) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n542), .Z(n794) );
  NAND2_X1 U596 ( .A1(G64), .A2(n794), .ZN(n545) );
  XOR2_X1 U597 ( .A(KEYINPUT0), .B(G543), .Z(n579) );
  NOR2_X1 U598 ( .A1(G651), .A2(n579), .ZN(n543) );
  XNOR2_X1 U599 ( .A(KEYINPUT66), .B(n543), .ZN(n801) );
  NAND2_X1 U600 ( .A1(G52), .A2(n801), .ZN(n544) );
  NAND2_X1 U601 ( .A1(n545), .A2(n544), .ZN(n552) );
  NOR2_X1 U602 ( .A1(G651), .A2(G543), .ZN(n793) );
  NAND2_X1 U603 ( .A1(G90), .A2(n793), .ZN(n548) );
  NOR2_X1 U604 ( .A1(n579), .A2(n546), .ZN(n797) );
  NAND2_X1 U605 ( .A1(G77), .A2(n797), .ZN(n547) );
  NAND2_X1 U606 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U607 ( .A(KEYINPUT72), .B(n549), .Z(n550) );
  XNOR2_X1 U608 ( .A(KEYINPUT9), .B(n550), .ZN(n551) );
  NOR2_X1 U609 ( .A1(n552), .A2(n551), .ZN(G171) );
  NAND2_X1 U610 ( .A1(G78), .A2(n797), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G53), .A2(n801), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n558) );
  NAND2_X1 U613 ( .A1(G91), .A2(n793), .ZN(n556) );
  NAND2_X1 U614 ( .A1(G65), .A2(n794), .ZN(n555) );
  NAND2_X1 U615 ( .A1(n556), .A2(n555), .ZN(n557) );
  NOR2_X1 U616 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U617 ( .A(n559), .B(KEYINPUT73), .ZN(G299) );
  NAND2_X1 U618 ( .A1(G89), .A2(n793), .ZN(n560) );
  XNOR2_X1 U619 ( .A(n560), .B(KEYINPUT4), .ZN(n561) );
  XNOR2_X1 U620 ( .A(KEYINPUT78), .B(n561), .ZN(n564) );
  NAND2_X1 U621 ( .A1(n797), .A2(G76), .ZN(n562) );
  XOR2_X1 U622 ( .A(KEYINPUT79), .B(n562), .Z(n563) );
  NAND2_X1 U623 ( .A1(n564), .A2(n563), .ZN(n565) );
  XNOR2_X1 U624 ( .A(n565), .B(KEYINPUT5), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G63), .A2(n794), .ZN(n567) );
  NAND2_X1 U626 ( .A1(G51), .A2(n801), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT6), .B(n568), .Z(n569) );
  NAND2_X1 U629 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U630 ( .A(n571), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U631 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U632 ( .A1(G88), .A2(n793), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G75), .A2(n797), .ZN(n572) );
  NAND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n577) );
  NAND2_X1 U635 ( .A1(G62), .A2(n794), .ZN(n575) );
  NAND2_X1 U636 ( .A1(G50), .A2(n801), .ZN(n574) );
  NAND2_X1 U637 ( .A1(n575), .A2(n574), .ZN(n576) );
  NOR2_X1 U638 ( .A1(n577), .A2(n576), .ZN(G166) );
  NAND2_X1 U639 ( .A1(n801), .A2(G49), .ZN(n578) );
  XNOR2_X1 U640 ( .A(n578), .B(KEYINPUT86), .ZN(n584) );
  NAND2_X1 U641 ( .A1(G87), .A2(n579), .ZN(n581) );
  NAND2_X1 U642 ( .A1(G74), .A2(G651), .ZN(n580) );
  NAND2_X1 U643 ( .A1(n581), .A2(n580), .ZN(n582) );
  NOR2_X1 U644 ( .A1(n794), .A2(n582), .ZN(n583) );
  NAND2_X1 U645 ( .A1(n584), .A2(n583), .ZN(G288) );
  INV_X1 U646 ( .A(G166), .ZN(G303) );
  NAND2_X1 U647 ( .A1(G73), .A2(n797), .ZN(n585) );
  XNOR2_X1 U648 ( .A(n585), .B(KEYINPUT2), .ZN(n592) );
  NAND2_X1 U649 ( .A1(G61), .A2(n794), .ZN(n587) );
  NAND2_X1 U650 ( .A1(G48), .A2(n801), .ZN(n586) );
  NAND2_X1 U651 ( .A1(n587), .A2(n586), .ZN(n590) );
  NAND2_X1 U652 ( .A1(G86), .A2(n793), .ZN(n588) );
  XNOR2_X1 U653 ( .A(KEYINPUT87), .B(n588), .ZN(n589) );
  NOR2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  NAND2_X1 U655 ( .A1(n592), .A2(n591), .ZN(G305) );
  NAND2_X1 U656 ( .A1(n793), .A2(G85), .ZN(n593) );
  XNOR2_X1 U657 ( .A(n593), .B(KEYINPUT70), .ZN(n595) );
  NAND2_X1 U658 ( .A1(G72), .A2(n797), .ZN(n594) );
  NAND2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n596), .ZN(n600) );
  NAND2_X1 U661 ( .A1(n801), .A2(G47), .ZN(n598) );
  NAND2_X1 U662 ( .A1(G60), .A2(n794), .ZN(n597) );
  AND2_X1 U663 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n600), .A2(n599), .ZN(G290) );
  INV_X1 U665 ( .A(KEYINPUT95), .ZN(n603) );
  NAND2_X1 U666 ( .A1(G40), .A2(G160), .ZN(n602) );
  XNOR2_X1 U667 ( .A(n603), .B(n602), .ZN(n694) );
  INV_X1 U668 ( .A(n694), .ZN(n604) );
  NAND2_X2 U669 ( .A1(n695), .A2(n604), .ZN(n664) );
  NAND2_X1 U670 ( .A1(G8), .A2(n664), .ZN(n741) );
  XNOR2_X1 U671 ( .A(G2078), .B(KEYINPUT25), .ZN(n926) );
  INV_X1 U672 ( .A(KEYINPUT102), .ZN(n605) );
  XNOR2_X1 U673 ( .A(n664), .B(n605), .ZN(n641) );
  NAND2_X1 U674 ( .A1(n926), .A2(n641), .ZN(n607) );
  INV_X1 U675 ( .A(G1961), .ZN(n1002) );
  NAND2_X1 U676 ( .A1(n664), .A2(n1002), .ZN(n606) );
  NAND2_X1 U677 ( .A1(n607), .A2(n606), .ZN(n658) );
  NAND2_X1 U678 ( .A1(n658), .A2(G171), .ZN(n654) );
  NAND2_X1 U679 ( .A1(G56), .A2(n794), .ZN(n608) );
  XOR2_X1 U680 ( .A(KEYINPUT14), .B(n608), .Z(n614) );
  NAND2_X1 U681 ( .A1(n793), .A2(G81), .ZN(n609) );
  XNOR2_X1 U682 ( .A(n609), .B(KEYINPUT12), .ZN(n611) );
  NAND2_X1 U683 ( .A1(G68), .A2(n797), .ZN(n610) );
  NAND2_X1 U684 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U685 ( .A(KEYINPUT13), .B(n612), .Z(n613) );
  NOR2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n616) );
  NAND2_X1 U687 ( .A1(G43), .A2(n801), .ZN(n615) );
  NAND2_X1 U688 ( .A1(n616), .A2(n615), .ZN(n973) );
  INV_X1 U689 ( .A(G1996), .ZN(n923) );
  NOR2_X1 U690 ( .A1(n664), .A2(n923), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n618), .B(n617), .ZN(n620) );
  NAND2_X1 U692 ( .A1(n664), .A2(G1341), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G92), .A2(n793), .ZN(n623) );
  NAND2_X1 U695 ( .A1(G66), .A2(n794), .ZN(n622) );
  NAND2_X1 U696 ( .A1(n623), .A2(n622), .ZN(n627) );
  NAND2_X1 U697 ( .A1(G79), .A2(n797), .ZN(n625) );
  NAND2_X1 U698 ( .A1(G54), .A2(n801), .ZN(n624) );
  NAND2_X1 U699 ( .A1(n625), .A2(n624), .ZN(n626) );
  NOR2_X1 U700 ( .A1(n627), .A2(n626), .ZN(n629) );
  XNOR2_X1 U701 ( .A(KEYINPUT15), .B(KEYINPUT76), .ZN(n628) );
  XNOR2_X1 U702 ( .A(n629), .B(n628), .ZN(n630) );
  XNOR2_X1 U703 ( .A(KEYINPUT77), .B(n630), .ZN(n994) );
  NAND2_X1 U704 ( .A1(n638), .A2(n994), .ZN(n635) );
  NAND2_X1 U705 ( .A1(G2067), .A2(n641), .ZN(n632) );
  NAND2_X1 U706 ( .A1(G1348), .A2(n664), .ZN(n631) );
  NAND2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n633) );
  XNOR2_X1 U708 ( .A(n633), .B(KEYINPUT104), .ZN(n634) );
  NAND2_X1 U709 ( .A1(n635), .A2(n634), .ZN(n637) );
  OR2_X1 U710 ( .A1(n994), .A2(n638), .ZN(n639) );
  NAND2_X1 U711 ( .A1(n640), .A2(n639), .ZN(n646) );
  INV_X1 U712 ( .A(G299), .ZN(n976) );
  NAND2_X1 U713 ( .A1(n641), .A2(G2072), .ZN(n642) );
  XNOR2_X1 U714 ( .A(n642), .B(KEYINPUT27), .ZN(n644) );
  XNOR2_X1 U715 ( .A(G1956), .B(KEYINPUT103), .ZN(n1003) );
  NOR2_X1 U716 ( .A1(n641), .A2(n1003), .ZN(n643) );
  NOR2_X1 U717 ( .A1(n644), .A2(n643), .ZN(n647) );
  NAND2_X1 U718 ( .A1(n976), .A2(n647), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n650) );
  NOR2_X1 U720 ( .A1(n976), .A2(n647), .ZN(n648) );
  XOR2_X1 U721 ( .A(n648), .B(KEYINPUT28), .Z(n649) );
  NAND2_X1 U722 ( .A1(n650), .A2(n649), .ZN(n652) );
  XOR2_X1 U723 ( .A(KEYINPUT29), .B(KEYINPUT106), .Z(n651) );
  XNOR2_X1 U724 ( .A(n652), .B(n651), .ZN(n653) );
  NAND2_X1 U725 ( .A1(n654), .A2(n653), .ZN(n663) );
  NOR2_X1 U726 ( .A1(G1966), .A2(n741), .ZN(n677) );
  NOR2_X1 U727 ( .A1(G2084), .A2(n664), .ZN(n674) );
  NOR2_X1 U728 ( .A1(n677), .A2(n674), .ZN(n655) );
  NAND2_X1 U729 ( .A1(G8), .A2(n655), .ZN(n656) );
  XNOR2_X1 U730 ( .A(KEYINPUT30), .B(n656), .ZN(n657) );
  NOR2_X1 U731 ( .A1(G168), .A2(n657), .ZN(n660) );
  NOR2_X1 U732 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U733 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U734 ( .A(KEYINPUT31), .B(n661), .Z(n662) );
  NAND2_X1 U735 ( .A1(n663), .A2(n662), .ZN(n675) );
  NAND2_X1 U736 ( .A1(n675), .A2(G286), .ZN(n671) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n664), .ZN(n665) );
  XNOR2_X1 U738 ( .A(KEYINPUT107), .B(n665), .ZN(n668) );
  NOR2_X1 U739 ( .A1(G1971), .A2(n741), .ZN(n666) );
  NOR2_X1 U740 ( .A1(G166), .A2(n666), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n668), .A2(n667), .ZN(n669) );
  XNOR2_X1 U742 ( .A(n669), .B(KEYINPUT108), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n671), .A2(n670), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n672), .A2(G8), .ZN(n673) );
  XNOR2_X1 U745 ( .A(n673), .B(KEYINPUT32), .ZN(n681) );
  NAND2_X1 U746 ( .A1(G8), .A2(n674), .ZN(n679) );
  INV_X1 U747 ( .A(n675), .ZN(n676) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U749 ( .A1(n679), .A2(n678), .ZN(n680) );
  NAND2_X1 U750 ( .A1(n681), .A2(n680), .ZN(n739) );
  NOR2_X1 U751 ( .A1(G1976), .A2(G288), .ZN(n978) );
  NOR2_X1 U752 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U753 ( .A1(n978), .A2(n682), .ZN(n683) );
  NAND2_X1 U754 ( .A1(n739), .A2(n683), .ZN(n684) );
  NAND2_X1 U755 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NAND2_X1 U756 ( .A1(n684), .A2(n979), .ZN(n685) );
  NOR2_X1 U757 ( .A1(n741), .A2(n685), .ZN(n687) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(n689) );
  NAND2_X1 U759 ( .A1(n689), .A2(n688), .ZN(n733) );
  NAND2_X1 U760 ( .A1(n978), .A2(KEYINPUT33), .ZN(n690) );
  NOR2_X1 U761 ( .A1(n690), .A2(n741), .ZN(n693) );
  XNOR2_X1 U762 ( .A(G1981), .B(KEYINPUT109), .ZN(n691) );
  XNOR2_X1 U763 ( .A(n691), .B(G305), .ZN(n989) );
  INV_X1 U764 ( .A(n989), .ZN(n692) );
  NOR2_X1 U765 ( .A1(n693), .A2(n692), .ZN(n731) );
  NOR2_X1 U766 ( .A1(n695), .A2(n694), .ZN(n760) );
  XNOR2_X1 U767 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  XNOR2_X1 U768 ( .A(KEYINPUT35), .B(KEYINPUT97), .ZN(n701) );
  NAND2_X1 U769 ( .A1(G128), .A2(n889), .ZN(n699) );
  NAND2_X1 U770 ( .A1(G116), .A2(n697), .ZN(n698) );
  NAND2_X1 U771 ( .A1(n699), .A2(n698), .ZN(n700) );
  XNOR2_X1 U772 ( .A(n701), .B(n700), .ZN(n708) );
  BUF_X1 U773 ( .A(n702), .Z(n886) );
  NAND2_X1 U774 ( .A1(n886), .A2(G104), .ZN(n703) );
  XNOR2_X1 U775 ( .A(n703), .B(KEYINPUT96), .ZN(n705) );
  NAND2_X1 U776 ( .A1(G140), .A2(n885), .ZN(n704) );
  NAND2_X1 U777 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U778 ( .A(KEYINPUT34), .B(n706), .ZN(n707) );
  NOR2_X1 U779 ( .A1(n708), .A2(n707), .ZN(n709) );
  XNOR2_X1 U780 ( .A(KEYINPUT36), .B(n709), .ZN(n882) );
  NOR2_X1 U781 ( .A1(n758), .A2(n882), .ZN(n710) );
  XNOR2_X1 U782 ( .A(KEYINPUT98), .B(n710), .ZN(n962) );
  NAND2_X1 U783 ( .A1(n760), .A2(n962), .ZN(n755) );
  NAND2_X1 U784 ( .A1(G131), .A2(n885), .ZN(n712) );
  NAND2_X1 U785 ( .A1(G95), .A2(n886), .ZN(n711) );
  NAND2_X1 U786 ( .A1(n712), .A2(n711), .ZN(n716) );
  NAND2_X1 U787 ( .A1(G119), .A2(n889), .ZN(n714) );
  NAND2_X1 U788 ( .A1(G107), .A2(n697), .ZN(n713) );
  NAND2_X1 U789 ( .A1(n714), .A2(n713), .ZN(n715) );
  OR2_X1 U790 ( .A1(n716), .A2(n715), .ZN(n881) );
  AND2_X1 U791 ( .A1(n881), .A2(G1991), .ZN(n727) );
  NAND2_X1 U792 ( .A1(G105), .A2(n886), .ZN(n717) );
  XOR2_X1 U793 ( .A(KEYINPUT38), .B(n717), .Z(n718) );
  XNOR2_X1 U794 ( .A(n718), .B(KEYINPUT99), .ZN(n720) );
  NAND2_X1 U795 ( .A1(G129), .A2(n889), .ZN(n719) );
  NAND2_X1 U796 ( .A1(n720), .A2(n719), .ZN(n724) );
  NAND2_X1 U797 ( .A1(n885), .A2(G141), .ZN(n722) );
  NAND2_X1 U798 ( .A1(G117), .A2(n697), .ZN(n721) );
  NAND2_X1 U799 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U800 ( .A1(n724), .A2(n723), .ZN(n725) );
  XNOR2_X1 U801 ( .A(KEYINPUT100), .B(n725), .ZN(n876) );
  NOR2_X1 U802 ( .A1(n923), .A2(n876), .ZN(n726) );
  NOR2_X1 U803 ( .A1(n727), .A2(n726), .ZN(n945) );
  INV_X1 U804 ( .A(n760), .ZN(n728) );
  NOR2_X1 U805 ( .A1(n945), .A2(n728), .ZN(n752) );
  INV_X1 U806 ( .A(n752), .ZN(n729) );
  NAND2_X1 U807 ( .A1(n755), .A2(n729), .ZN(n745) );
  INV_X1 U808 ( .A(n745), .ZN(n730) );
  AND2_X1 U809 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U810 ( .A1(n733), .A2(n732), .ZN(n747) );
  NOR2_X1 U811 ( .A1(G1981), .A2(G305), .ZN(n734) );
  XNOR2_X1 U812 ( .A(n734), .B(KEYINPUT24), .ZN(n735) );
  XNOR2_X1 U813 ( .A(KEYINPUT101), .B(n735), .ZN(n736) );
  OR2_X1 U814 ( .A1(n741), .A2(n736), .ZN(n743) );
  NOR2_X1 U815 ( .A1(G2090), .A2(G303), .ZN(n737) );
  NAND2_X1 U816 ( .A1(G8), .A2(n737), .ZN(n738) );
  NAND2_X1 U817 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U818 ( .A1(n741), .A2(n740), .ZN(n742) );
  AND2_X1 U819 ( .A1(n743), .A2(n742), .ZN(n744) );
  OR2_X1 U820 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n749) );
  XNOR2_X1 U822 ( .A(G1986), .B(G290), .ZN(n982) );
  NAND2_X1 U823 ( .A1(n982), .A2(n760), .ZN(n748) );
  NAND2_X1 U824 ( .A1(n749), .A2(n748), .ZN(n763) );
  AND2_X1 U825 ( .A1(n923), .A2(n876), .ZN(n949) );
  NOR2_X1 U826 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U827 ( .A1(G1991), .A2(n881), .ZN(n942) );
  NOR2_X1 U828 ( .A1(n750), .A2(n942), .ZN(n751) );
  NOR2_X1 U829 ( .A1(n752), .A2(n751), .ZN(n753) );
  NOR2_X1 U830 ( .A1(n949), .A2(n753), .ZN(n754) );
  XNOR2_X1 U831 ( .A(n754), .B(KEYINPUT39), .ZN(n756) );
  NAND2_X1 U832 ( .A1(n756), .A2(n755), .ZN(n757) );
  XNOR2_X1 U833 ( .A(n757), .B(KEYINPUT110), .ZN(n759) );
  NAND2_X1 U834 ( .A1(n758), .A2(n882), .ZN(n951) );
  NAND2_X1 U835 ( .A1(n759), .A2(n951), .ZN(n761) );
  NAND2_X1 U836 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U837 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U838 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U839 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U840 ( .A(G69), .ZN(G235) );
  INV_X1 U841 ( .A(G108), .ZN(G238) );
  INV_X1 U842 ( .A(G132), .ZN(G219) );
  INV_X1 U843 ( .A(G82), .ZN(G220) );
  XOR2_X1 U844 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n766) );
  NAND2_X1 U845 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U846 ( .A(n766), .B(n765), .ZN(G223) );
  INV_X1 U847 ( .A(G223), .ZN(n833) );
  NAND2_X1 U848 ( .A1(n833), .A2(G567), .ZN(n767) );
  XOR2_X1 U849 ( .A(KEYINPUT11), .B(n767), .Z(G234) );
  INV_X1 U850 ( .A(G860), .ZN(n772) );
  OR2_X1 U851 ( .A1(n973), .A2(n772), .ZN(G153) );
  INV_X1 U852 ( .A(G171), .ZN(G301) );
  INV_X1 U853 ( .A(n994), .ZN(n898) );
  NOR2_X1 U854 ( .A1(n898), .A2(G868), .ZN(n769) );
  INV_X1 U855 ( .A(G868), .ZN(n814) );
  NOR2_X1 U856 ( .A1(n814), .A2(G301), .ZN(n768) );
  NOR2_X1 U857 ( .A1(n769), .A2(n768), .ZN(G284) );
  NAND2_X1 U858 ( .A1(G286), .A2(G868), .ZN(n771) );
  NAND2_X1 U859 ( .A1(G299), .A2(n814), .ZN(n770) );
  NAND2_X1 U860 ( .A1(n771), .A2(n770), .ZN(G297) );
  NAND2_X1 U861 ( .A1(n772), .A2(G559), .ZN(n773) );
  NAND2_X1 U862 ( .A1(n773), .A2(n994), .ZN(n774) );
  XNOR2_X1 U863 ( .A(n774), .B(KEYINPUT80), .ZN(n775) );
  XNOR2_X1 U864 ( .A(KEYINPUT16), .B(n775), .ZN(G148) );
  NOR2_X1 U865 ( .A1(G868), .A2(n973), .ZN(n776) );
  XOR2_X1 U866 ( .A(KEYINPUT81), .B(n776), .Z(n779) );
  NAND2_X1 U867 ( .A1(G868), .A2(n994), .ZN(n777) );
  NOR2_X1 U868 ( .A1(G559), .A2(n777), .ZN(n778) );
  NOR2_X1 U869 ( .A1(n779), .A2(n778), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G123), .A2(n889), .ZN(n780) );
  XNOR2_X1 U871 ( .A(n780), .B(KEYINPUT18), .ZN(n781) );
  XNOR2_X1 U872 ( .A(KEYINPUT82), .B(n781), .ZN(n784) );
  NAND2_X1 U873 ( .A1(G99), .A2(n886), .ZN(n782) );
  XOR2_X1 U874 ( .A(KEYINPUT83), .B(n782), .Z(n783) );
  NAND2_X1 U875 ( .A1(n784), .A2(n783), .ZN(n788) );
  NAND2_X1 U876 ( .A1(n885), .A2(G135), .ZN(n786) );
  NAND2_X1 U877 ( .A1(G111), .A2(n697), .ZN(n785) );
  NAND2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  NOR2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n941) );
  XNOR2_X1 U880 ( .A(G2096), .B(n941), .ZN(n790) );
  INV_X1 U881 ( .A(G2100), .ZN(n789) );
  NAND2_X1 U882 ( .A1(n790), .A2(n789), .ZN(G156) );
  XNOR2_X1 U883 ( .A(KEYINPUT84), .B(n973), .ZN(n791) );
  NAND2_X1 U884 ( .A1(G559), .A2(n994), .ZN(n812) );
  XNOR2_X1 U885 ( .A(n791), .B(n812), .ZN(n792) );
  NOR2_X1 U886 ( .A1(G860), .A2(n792), .ZN(n804) );
  NAND2_X1 U887 ( .A1(G93), .A2(n793), .ZN(n796) );
  NAND2_X1 U888 ( .A1(G67), .A2(n794), .ZN(n795) );
  NAND2_X1 U889 ( .A1(n796), .A2(n795), .ZN(n800) );
  NAND2_X1 U890 ( .A1(G80), .A2(n797), .ZN(n798) );
  XNOR2_X1 U891 ( .A(KEYINPUT85), .B(n798), .ZN(n799) );
  NOR2_X1 U892 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U893 ( .A1(G55), .A2(n801), .ZN(n802) );
  NAND2_X1 U894 ( .A1(n803), .A2(n802), .ZN(n815) );
  XOR2_X1 U895 ( .A(n804), .B(n815), .Z(G145) );
  XNOR2_X1 U896 ( .A(G305), .B(n815), .ZN(n811) );
  XNOR2_X1 U897 ( .A(G290), .B(n973), .ZN(n809) );
  XNOR2_X1 U898 ( .A(G166), .B(KEYINPUT19), .ZN(n805) );
  XNOR2_X1 U899 ( .A(n805), .B(KEYINPUT88), .ZN(n806) );
  XNOR2_X1 U900 ( .A(n976), .B(n806), .ZN(n807) );
  XNOR2_X1 U901 ( .A(n807), .B(G288), .ZN(n808) );
  XNOR2_X1 U902 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U903 ( .A(n811), .B(n810), .ZN(n901) );
  XOR2_X1 U904 ( .A(n901), .B(n812), .Z(n813) );
  NOR2_X1 U905 ( .A1(n814), .A2(n813), .ZN(n817) );
  NOR2_X1 U906 ( .A1(G868), .A2(n815), .ZN(n816) );
  NOR2_X1 U907 ( .A1(n817), .A2(n816), .ZN(G295) );
  NAND2_X1 U908 ( .A1(G2084), .A2(G2078), .ZN(n818) );
  XNOR2_X1 U909 ( .A(n818), .B(KEYINPUT20), .ZN(n819) );
  XNOR2_X1 U910 ( .A(KEYINPUT89), .B(n819), .ZN(n820) );
  NAND2_X1 U911 ( .A1(n820), .A2(G2090), .ZN(n821) );
  XNOR2_X1 U912 ( .A(KEYINPUT21), .B(n821), .ZN(n822) );
  NAND2_X1 U913 ( .A1(n822), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U914 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  XOR2_X1 U915 ( .A(KEYINPUT74), .B(G57), .Z(G237) );
  NOR2_X1 U916 ( .A1(G220), .A2(G219), .ZN(n823) );
  XOR2_X1 U917 ( .A(KEYINPUT22), .B(n823), .Z(n824) );
  NOR2_X1 U918 ( .A1(G218), .A2(n824), .ZN(n825) );
  XNOR2_X1 U919 ( .A(KEYINPUT90), .B(n825), .ZN(n826) );
  NAND2_X1 U920 ( .A1(n826), .A2(G96), .ZN(n839) );
  NAND2_X1 U921 ( .A1(n839), .A2(G2106), .ZN(n831) );
  NOR2_X1 U922 ( .A1(G237), .A2(G238), .ZN(n827) );
  NAND2_X1 U923 ( .A1(G120), .A2(n827), .ZN(n828) );
  NOR2_X1 U924 ( .A1(n828), .A2(G235), .ZN(n829) );
  XNOR2_X1 U925 ( .A(n829), .B(KEYINPUT91), .ZN(n838) );
  NAND2_X1 U926 ( .A1(n838), .A2(G567), .ZN(n830) );
  NAND2_X1 U927 ( .A1(n831), .A2(n830), .ZN(n841) );
  NAND2_X1 U928 ( .A1(G661), .A2(G483), .ZN(n832) );
  NOR2_X1 U929 ( .A1(n841), .A2(n832), .ZN(n837) );
  NAND2_X1 U930 ( .A1(n837), .A2(G36), .ZN(G176) );
  NAND2_X1 U931 ( .A1(n833), .A2(G2106), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n834), .B(KEYINPUT112), .ZN(G217) );
  AND2_X1 U933 ( .A1(G15), .A2(G2), .ZN(n835) );
  NAND2_X1 U934 ( .A1(G661), .A2(n835), .ZN(G259) );
  NAND2_X1 U935 ( .A1(G3), .A2(G1), .ZN(n836) );
  NAND2_X1 U936 ( .A1(n837), .A2(n836), .ZN(G188) );
  XNOR2_X1 U937 ( .A(G120), .B(KEYINPUT113), .ZN(G236) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n839), .A2(n838), .ZN(n840) );
  XNOR2_X1 U941 ( .A(n840), .B(KEYINPUT114), .ZN(G325) );
  INV_X1 U942 ( .A(G325), .ZN(G261) );
  INV_X1 U943 ( .A(n841), .ZN(G319) );
  XOR2_X1 U944 ( .A(KEYINPUT115), .B(G2084), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2072), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U947 ( .A(n844), .B(G2096), .Z(n846) );
  XNOR2_X1 U948 ( .A(G2067), .B(G2090), .ZN(n845) );
  XNOR2_X1 U949 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U950 ( .A(KEYINPUT43), .B(G2678), .Z(n848) );
  XNOR2_X1 U951 ( .A(KEYINPUT42), .B(G2100), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U953 ( .A(n850), .B(n849), .Z(G227) );
  XOR2_X1 U954 ( .A(G1971), .B(G1956), .Z(n852) );
  XNOR2_X1 U955 ( .A(G1966), .B(G1961), .ZN(n851) );
  XNOR2_X1 U956 ( .A(n852), .B(n851), .ZN(n853) );
  XOR2_X1 U957 ( .A(n853), .B(G2474), .Z(n855) );
  XNOR2_X1 U958 ( .A(G1986), .B(G1976), .ZN(n854) );
  XNOR2_X1 U959 ( .A(n855), .B(n854), .ZN(n859) );
  XOR2_X1 U960 ( .A(KEYINPUT41), .B(G1981), .Z(n857) );
  XNOR2_X1 U961 ( .A(G1996), .B(G1991), .ZN(n856) );
  XNOR2_X1 U962 ( .A(n857), .B(n856), .ZN(n858) );
  XNOR2_X1 U963 ( .A(n859), .B(n858), .ZN(G229) );
  NAND2_X1 U964 ( .A1(n889), .A2(G124), .ZN(n860) );
  XNOR2_X1 U965 ( .A(n860), .B(KEYINPUT44), .ZN(n862) );
  NAND2_X1 U966 ( .A1(G100), .A2(n886), .ZN(n861) );
  NAND2_X1 U967 ( .A1(n862), .A2(n861), .ZN(n866) );
  NAND2_X1 U968 ( .A1(n885), .A2(G136), .ZN(n864) );
  NAND2_X1 U969 ( .A1(G112), .A2(n697), .ZN(n863) );
  NAND2_X1 U970 ( .A1(n864), .A2(n863), .ZN(n865) );
  NOR2_X1 U971 ( .A1(n866), .A2(n865), .ZN(G162) );
  XOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n868) );
  XNOR2_X1 U973 ( .A(G162), .B(n941), .ZN(n867) );
  XNOR2_X1 U974 ( .A(n868), .B(n867), .ZN(n880) );
  NAND2_X1 U975 ( .A1(G130), .A2(n889), .ZN(n870) );
  NAND2_X1 U976 ( .A1(G118), .A2(n697), .ZN(n869) );
  NAND2_X1 U977 ( .A1(n870), .A2(n869), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G142), .A2(n885), .ZN(n872) );
  NAND2_X1 U979 ( .A1(G106), .A2(n886), .ZN(n871) );
  NAND2_X1 U980 ( .A1(n872), .A2(n871), .ZN(n873) );
  XOR2_X1 U981 ( .A(n873), .B(KEYINPUT45), .Z(n874) );
  NOR2_X1 U982 ( .A1(n875), .A2(n874), .ZN(n877) );
  XNOR2_X1 U983 ( .A(n877), .B(n876), .ZN(n878) );
  XOR2_X1 U984 ( .A(G160), .B(n878), .Z(n879) );
  XNOR2_X1 U985 ( .A(n880), .B(n879), .ZN(n884) );
  XOR2_X1 U986 ( .A(n882), .B(n881), .Z(n883) );
  XNOR2_X1 U987 ( .A(n884), .B(n883), .ZN(n896) );
  NAND2_X1 U988 ( .A1(G139), .A2(n885), .ZN(n888) );
  NAND2_X1 U989 ( .A1(G103), .A2(n886), .ZN(n887) );
  NAND2_X1 U990 ( .A1(n888), .A2(n887), .ZN(n894) );
  NAND2_X1 U991 ( .A1(G127), .A2(n889), .ZN(n891) );
  NAND2_X1 U992 ( .A1(G115), .A2(n697), .ZN(n890) );
  NAND2_X1 U993 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U994 ( .A(KEYINPUT47), .B(n892), .Z(n893) );
  NOR2_X1 U995 ( .A1(n894), .A2(n893), .ZN(n953) );
  XNOR2_X1 U996 ( .A(G164), .B(n953), .ZN(n895) );
  XNOR2_X1 U997 ( .A(n896), .B(n895), .ZN(n897) );
  NOR2_X1 U998 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U999 ( .A(KEYINPUT116), .B(G286), .Z(n900) );
  XNOR2_X1 U1000 ( .A(G171), .B(n898), .ZN(n899) );
  XNOR2_X1 U1001 ( .A(n900), .B(n899), .ZN(n902) );
  XNOR2_X1 U1002 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1003 ( .A1(G37), .A2(n903), .ZN(G397) );
  XOR2_X1 U1004 ( .A(G2454), .B(G2435), .Z(n905) );
  XNOR2_X1 U1005 ( .A(G2438), .B(G2427), .ZN(n904) );
  XNOR2_X1 U1006 ( .A(n905), .B(n904), .ZN(n912) );
  XOR2_X1 U1007 ( .A(KEYINPUT111), .B(G2446), .Z(n907) );
  XNOR2_X1 U1008 ( .A(G2443), .B(G2430), .ZN(n906) );
  XNOR2_X1 U1009 ( .A(n907), .B(n906), .ZN(n908) );
  XOR2_X1 U1010 ( .A(n908), .B(G2451), .Z(n910) );
  XNOR2_X1 U1011 ( .A(G1341), .B(G1348), .ZN(n909) );
  XNOR2_X1 U1012 ( .A(n910), .B(n909), .ZN(n911) );
  XNOR2_X1 U1013 ( .A(n912), .B(n911), .ZN(n913) );
  NAND2_X1 U1014 ( .A1(n913), .A2(G14), .ZN(n920) );
  NAND2_X1 U1015 ( .A1(G319), .A2(n920), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(G227), .A2(G229), .ZN(n914) );
  XOR2_X1 U1017 ( .A(KEYINPUT49), .B(n914), .Z(n915) );
  XNOR2_X1 U1018 ( .A(n915), .B(KEYINPUT117), .ZN(n916) );
  NOR2_X1 U1019 ( .A1(n917), .A2(n916), .ZN(n919) );
  NOR2_X1 U1020 ( .A1(G395), .A2(G397), .ZN(n918) );
  NAND2_X1 U1021 ( .A1(n919), .A2(n918), .ZN(G225) );
  INV_X1 U1022 ( .A(G225), .ZN(G308) );
  INV_X1 U1023 ( .A(n920), .ZN(G401) );
  XOR2_X1 U1024 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n1033) );
  XNOR2_X1 U1025 ( .A(G2090), .B(G35), .ZN(n935) );
  XOR2_X1 U1026 ( .A(G25), .B(G1991), .Z(n921) );
  NAND2_X1 U1027 ( .A1(n921), .A2(G28), .ZN(n932) );
  XNOR2_X1 U1028 ( .A(KEYINPUT119), .B(G2072), .ZN(n922) );
  XNOR2_X1 U1029 ( .A(n922), .B(G33), .ZN(n930) );
  XOR2_X1 U1030 ( .A(G2067), .B(G26), .Z(n925) );
  XNOR2_X1 U1031 ( .A(n923), .B(G32), .ZN(n924) );
  NAND2_X1 U1032 ( .A1(n925), .A2(n924), .ZN(n928) );
  XOR2_X1 U1033 ( .A(G27), .B(n926), .Z(n927) );
  NOR2_X1 U1034 ( .A1(n928), .A2(n927), .ZN(n929) );
  NAND2_X1 U1035 ( .A1(n930), .A2(n929), .ZN(n931) );
  NOR2_X1 U1036 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1037 ( .A(KEYINPUT53), .B(n933), .ZN(n934) );
  NOR2_X1 U1038 ( .A1(n935), .A2(n934), .ZN(n938) );
  XOR2_X1 U1039 ( .A(G2084), .B(G34), .Z(n936) );
  XNOR2_X1 U1040 ( .A(KEYINPUT54), .B(n936), .ZN(n937) );
  NAND2_X1 U1041 ( .A1(n938), .A2(n937), .ZN(n966) );
  NOR2_X1 U1042 ( .A1(G29), .A2(KEYINPUT55), .ZN(n939) );
  NAND2_X1 U1043 ( .A1(n966), .A2(n939), .ZN(n940) );
  NAND2_X1 U1044 ( .A1(G11), .A2(n940), .ZN(n971) );
  NOR2_X1 U1045 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1046 ( .A(n943), .B(KEYINPUT118), .ZN(n944) );
  NAND2_X1 U1047 ( .A1(n945), .A2(n944), .ZN(n947) );
  XOR2_X1 U1048 ( .A(G160), .B(G2084), .Z(n946) );
  NOR2_X1 U1049 ( .A1(n947), .A2(n946), .ZN(n960) );
  XOR2_X1 U1050 ( .A(G2090), .B(G162), .Z(n948) );
  NOR2_X1 U1051 ( .A1(n949), .A2(n948), .ZN(n950) );
  XOR2_X1 U1052 ( .A(KEYINPUT51), .B(n950), .Z(n952) );
  NAND2_X1 U1053 ( .A1(n952), .A2(n951), .ZN(n958) );
  XOR2_X1 U1054 ( .A(G2072), .B(n953), .Z(n955) );
  XOR2_X1 U1055 ( .A(G164), .B(G2078), .Z(n954) );
  NOR2_X1 U1056 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1057 ( .A(KEYINPUT50), .B(n956), .Z(n957) );
  NOR2_X1 U1058 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1059 ( .A1(n960), .A2(n959), .ZN(n961) );
  NOR2_X1 U1060 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1061 ( .A(KEYINPUT52), .B(n963), .ZN(n964) );
  INV_X1 U1062 ( .A(KEYINPUT55), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n964), .A2(n967), .ZN(n965) );
  NAND2_X1 U1064 ( .A1(n965), .A2(G29), .ZN(n969) );
  OR2_X1 U1065 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1066 ( .A1(n969), .A2(n968), .ZN(n970) );
  NOR2_X1 U1067 ( .A1(n971), .A2(n970), .ZN(n1031) );
  XNOR2_X1 U1068 ( .A(G16), .B(KEYINPUT56), .ZN(n1001) );
  XNOR2_X1 U1069 ( .A(G171), .B(G1961), .ZN(n972) );
  XNOR2_X1 U1070 ( .A(n972), .B(KEYINPUT121), .ZN(n975) );
  XNOR2_X1 U1071 ( .A(G1341), .B(n973), .ZN(n974) );
  NOR2_X1 U1072 ( .A1(n975), .A2(n974), .ZN(n999) );
  XNOR2_X1 U1073 ( .A(G1956), .B(n976), .ZN(n977) );
  XNOR2_X1 U1074 ( .A(n977), .B(KEYINPUT122), .ZN(n984) );
  INV_X1 U1075 ( .A(n978), .ZN(n980) );
  NAND2_X1 U1076 ( .A1(n980), .A2(n979), .ZN(n981) );
  NOR2_X1 U1077 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1078 ( .A1(n984), .A2(n983), .ZN(n987) );
  XOR2_X1 U1079 ( .A(G1971), .B(G303), .Z(n985) );
  XNOR2_X1 U1080 ( .A(KEYINPUT123), .B(n985), .ZN(n986) );
  NOR2_X1 U1081 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1082 ( .A(KEYINPUT124), .B(n988), .ZN(n993) );
  XNOR2_X1 U1083 ( .A(G1966), .B(G168), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  XNOR2_X1 U1085 ( .A(n991), .B(KEYINPUT57), .ZN(n992) );
  NAND2_X1 U1086 ( .A1(n993), .A2(n992), .ZN(n997) );
  XOR2_X1 U1087 ( .A(G1348), .B(n994), .Z(n995) );
  XNOR2_X1 U1088 ( .A(KEYINPUT120), .B(n995), .ZN(n996) );
  NOR2_X1 U1089 ( .A1(n997), .A2(n996), .ZN(n998) );
  NAND2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1028) );
  INV_X1 U1092 ( .A(G16), .ZN(n1026) );
  XNOR2_X1 U1093 ( .A(G5), .B(n1002), .ZN(n1015) );
  XNOR2_X1 U1094 ( .A(G20), .B(n1003), .ZN(n1007) );
  XNOR2_X1 U1095 ( .A(G1341), .B(G19), .ZN(n1005) );
  XNOR2_X1 U1096 ( .A(G6), .B(G1981), .ZN(n1004) );
  NOR2_X1 U1097 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  NAND2_X1 U1098 ( .A1(n1007), .A2(n1006), .ZN(n1010) );
  XOR2_X1 U1099 ( .A(KEYINPUT59), .B(G1348), .Z(n1008) );
  XNOR2_X1 U1100 ( .A(G4), .B(n1008), .ZN(n1009) );
  NOR2_X1 U1101 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  XOR2_X1 U1102 ( .A(KEYINPUT60), .B(n1011), .Z(n1013) );
  XNOR2_X1 U1103 ( .A(G1966), .B(G21), .ZN(n1012) );
  NOR2_X1 U1104 ( .A1(n1013), .A2(n1012), .ZN(n1014) );
  NAND2_X1 U1105 ( .A1(n1015), .A2(n1014), .ZN(n1023) );
  XNOR2_X1 U1106 ( .A(G1971), .B(G22), .ZN(n1017) );
  XNOR2_X1 U1107 ( .A(G23), .B(G1976), .ZN(n1016) );
  NOR2_X1 U1108 ( .A1(n1017), .A2(n1016), .ZN(n1020) );
  XNOR2_X1 U1109 ( .A(G1986), .B(KEYINPUT125), .ZN(n1018) );
  XNOR2_X1 U1110 ( .A(n1018), .B(G24), .ZN(n1019) );
  NAND2_X1 U1111 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1112 ( .A(KEYINPUT58), .B(n1021), .ZN(n1022) );
  NOR2_X1 U1113 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  XNOR2_X1 U1114 ( .A(KEYINPUT61), .B(n1024), .ZN(n1025) );
  NAND2_X1 U1115 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NAND2_X1 U1116 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  XOR2_X1 U1117 ( .A(KEYINPUT126), .B(n1029), .Z(n1030) );
  NAND2_X1 U1118 ( .A1(n1031), .A2(n1030), .ZN(n1032) );
  XOR2_X1 U1119 ( .A(n1033), .B(n1032), .Z(G311) );
  INV_X1 U1120 ( .A(G311), .ZN(G150) );
endmodule

