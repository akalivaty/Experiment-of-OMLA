

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581;

  XOR2_X1 U322 ( .A(n362), .B(n361), .Z(n518) );
  XOR2_X1 U323 ( .A(KEYINPUT94), .B(n409), .Z(n515) );
  XOR2_X1 U324 ( .A(G120GAT), .B(G57GAT), .Z(n443) );
  INV_X1 U325 ( .A(KEYINPUT92), .ZN(n378) );
  XNOR2_X1 U326 ( .A(n444), .B(n443), .ZN(n445) );
  NOR2_X1 U327 ( .A1(n466), .A2(n465), .ZN(n467) );
  INV_X1 U328 ( .A(KEYINPUT37), .ZN(n414) );
  XNOR2_X1 U329 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U330 ( .A(n446), .B(n445), .ZN(n448) );
  XNOR2_X1 U331 ( .A(n414), .B(KEYINPUT103), .ZN(n415) );
  XNOR2_X1 U332 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U333 ( .A(n416), .B(n415), .ZN(n514) );
  XOR2_X1 U334 ( .A(n570), .B(KEYINPUT41), .Z(n559) );
  INV_X1 U335 ( .A(G43GAT), .ZN(n450) );
  XNOR2_X1 U336 ( .A(KEYINPUT38), .B(n449), .ZN(n498) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n475) );
  XNOR2_X1 U338 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U339 ( .A(n476), .B(n475), .ZN(G1351GAT) );
  XNOR2_X1 U340 ( .A(n453), .B(n452), .ZN(G1330GAT) );
  XOR2_X1 U341 ( .A(KEYINPUT64), .B(KEYINPUT76), .Z(n291) );
  XNOR2_X1 U342 ( .A(KEYINPUT10), .B(KEYINPUT65), .ZN(n290) );
  XNOR2_X1 U343 ( .A(n291), .B(n290), .ZN(n306) );
  XOR2_X1 U344 ( .A(G36GAT), .B(G190GAT), .Z(n355) );
  XOR2_X1 U345 ( .A(KEYINPUT11), .B(n355), .Z(n293) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G85GAT), .ZN(n447) );
  XOR2_X1 U347 ( .A(G218GAT), .B(n447), .Z(n292) );
  XNOR2_X1 U348 ( .A(n293), .B(n292), .ZN(n299) );
  XOR2_X1 U349 ( .A(G29GAT), .B(G134GAT), .Z(n370) );
  XOR2_X1 U350 ( .A(G43GAT), .B(KEYINPUT7), .Z(n295) );
  XNOR2_X1 U351 ( .A(KEYINPUT69), .B(KEYINPUT8), .ZN(n294) );
  XNOR2_X1 U352 ( .A(n295), .B(n294), .ZN(n421) );
  XOR2_X1 U353 ( .A(n370), .B(n421), .Z(n297) );
  NAND2_X1 U354 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U355 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U356 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U357 ( .A(G50GAT), .B(KEYINPUT75), .Z(n387) );
  XOR2_X1 U358 ( .A(KEYINPUT9), .B(G92GAT), .Z(n301) );
  XNOR2_X1 U359 ( .A(G162GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U360 ( .A(n301), .B(n300), .ZN(n302) );
  XNOR2_X1 U361 ( .A(n387), .B(n302), .ZN(n303) );
  XNOR2_X1 U362 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U363 ( .A(n306), .B(n305), .Z(n462) );
  XOR2_X1 U364 ( .A(KEYINPUT36), .B(n462), .Z(n578) );
  XOR2_X1 U365 ( .A(KEYINPUT12), .B(KEYINPUT84), .Z(n308) );
  XNOR2_X1 U366 ( .A(KEYINPUT83), .B(KEYINPUT82), .ZN(n307) );
  XNOR2_X1 U367 ( .A(n308), .B(n307), .ZN(n329) );
  XOR2_X1 U368 ( .A(KEYINPUT81), .B(KEYINPUT77), .Z(n310) );
  XNOR2_X1 U369 ( .A(G8GAT), .B(G64GAT), .ZN(n309) );
  XNOR2_X1 U370 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U371 ( .A(KEYINPUT80), .B(KEYINPUT79), .Z(n312) );
  XNOR2_X1 U372 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n311) );
  XNOR2_X1 U373 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U374 ( .A(n314), .B(n313), .Z(n327) );
  XOR2_X1 U375 ( .A(KEYINPUT70), .B(G1GAT), .Z(n316) );
  XNOR2_X1 U376 ( .A(G22GAT), .B(G15GAT), .ZN(n315) );
  XNOR2_X1 U377 ( .A(n316), .B(n315), .ZN(n418) );
  XOR2_X1 U378 ( .A(n418), .B(KEYINPUT14), .Z(n318) );
  NAND2_X1 U379 ( .A1(G231GAT), .A2(G233GAT), .ZN(n317) );
  XNOR2_X1 U380 ( .A(n318), .B(n317), .ZN(n325) );
  XOR2_X1 U381 ( .A(G57GAT), .B(G211GAT), .Z(n320) );
  XNOR2_X1 U382 ( .A(G127GAT), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U383 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U384 ( .A(G71GAT), .B(KEYINPUT13), .Z(n442) );
  XOR2_X1 U385 ( .A(n321), .B(n442), .Z(n323) );
  XNOR2_X1 U386 ( .A(G183GAT), .B(G78GAT), .ZN(n322) );
  XNOR2_X1 U387 ( .A(n323), .B(n322), .ZN(n324) );
  XNOR2_X1 U388 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U389 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n575) );
  INV_X1 U391 ( .A(n575), .ZN(n479) );
  NAND2_X1 U392 ( .A1(G227GAT), .A2(G233GAT), .ZN(n335) );
  XOR2_X1 U393 ( .A(G120GAT), .B(G190GAT), .Z(n331) );
  XNOR2_X1 U394 ( .A(G15GAT), .B(G99GAT), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n333) );
  XOR2_X1 U396 ( .A(G43GAT), .B(G134GAT), .Z(n332) );
  XNOR2_X1 U397 ( .A(n333), .B(n332), .ZN(n334) );
  XNOR2_X1 U398 ( .A(n335), .B(n334), .ZN(n348) );
  XOR2_X1 U399 ( .A(G176GAT), .B(KEYINPUT86), .Z(n337) );
  XNOR2_X1 U400 ( .A(KEYINPUT88), .B(KEYINPUT20), .ZN(n336) );
  XNOR2_X1 U401 ( .A(n337), .B(n336), .ZN(n346) );
  XOR2_X1 U402 ( .A(G127GAT), .B(KEYINPUT85), .Z(n339) );
  XNOR2_X1 U403 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n338) );
  XNOR2_X1 U404 ( .A(n339), .B(n338), .ZN(n377) );
  XOR2_X1 U405 ( .A(G71GAT), .B(n377), .Z(n344) );
  XOR2_X1 U406 ( .A(KEYINPUT18), .B(KEYINPUT87), .Z(n341) );
  XNOR2_X1 U407 ( .A(KEYINPUT17), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U408 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U409 ( .A(KEYINPUT19), .B(n342), .Z(n352) );
  XNOR2_X1 U410 ( .A(G169GAT), .B(n352), .ZN(n343) );
  XNOR2_X1 U411 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U412 ( .A(n346), .B(n345), .Z(n347) );
  XOR2_X1 U413 ( .A(n348), .B(n347), .Z(n520) );
  INV_X1 U414 ( .A(n520), .ZN(n528) );
  XOR2_X1 U415 ( .A(KEYINPUT89), .B(G218GAT), .Z(n350) );
  XNOR2_X1 U416 ( .A(KEYINPUT21), .B(G211GAT), .ZN(n349) );
  XNOR2_X1 U417 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U418 ( .A(G197GAT), .B(n351), .Z(n396) );
  XNOR2_X1 U419 ( .A(n352), .B(n396), .ZN(n362) );
  XOR2_X1 U420 ( .A(G64GAT), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U421 ( .A(G176GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U422 ( .A(n354), .B(n353), .ZN(n438) );
  XOR2_X1 U423 ( .A(n355), .B(n438), .Z(n357) );
  NAND2_X1 U424 ( .A1(G226GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U425 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U426 ( .A(n358), .B(KEYINPUT95), .Z(n360) );
  XOR2_X1 U427 ( .A(G169GAT), .B(G8GAT), .Z(n417) );
  XNOR2_X1 U428 ( .A(n417), .B(KEYINPUT77), .ZN(n359) );
  XNOR2_X1 U429 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U430 ( .A(n518), .B(KEYINPUT27), .ZN(n363) );
  XNOR2_X1 U431 ( .A(KEYINPUT96), .B(n363), .ZN(n403) );
  XNOR2_X1 U432 ( .A(G155GAT), .B(G162GAT), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n364), .B(KEYINPUT3), .ZN(n365) );
  XOR2_X1 U434 ( .A(n365), .B(KEYINPUT2), .Z(n367) );
  XNOR2_X1 U435 ( .A(G141GAT), .B(G148GAT), .ZN(n366) );
  XNOR2_X1 U436 ( .A(n367), .B(n366), .ZN(n397) );
  XOR2_X1 U437 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n369) );
  XNOR2_X1 U438 ( .A(G1GAT), .B(KEYINPUT6), .ZN(n368) );
  XNOR2_X1 U439 ( .A(n369), .B(n368), .ZN(n374) );
  XOR2_X1 U440 ( .A(KEYINPUT4), .B(G85GAT), .Z(n372) );
  XNOR2_X1 U441 ( .A(n370), .B(n443), .ZN(n371) );
  XNOR2_X1 U442 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U443 ( .A(n374), .B(n373), .Z(n376) );
  NAND2_X1 U444 ( .A1(G225GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U445 ( .A(n376), .B(n375), .ZN(n381) );
  XNOR2_X1 U446 ( .A(n377), .B(KEYINPUT93), .ZN(n379) );
  XOR2_X1 U447 ( .A(n397), .B(n382), .Z(n409) );
  NAND2_X1 U448 ( .A1(n403), .A2(n515), .ZN(n383) );
  XOR2_X1 U449 ( .A(KEYINPUT97), .B(n383), .Z(n525) );
  XOR2_X1 U450 ( .A(KEYINPUT24), .B(KEYINPUT91), .Z(n385) );
  XNOR2_X1 U451 ( .A(G204GAT), .B(KEYINPUT22), .ZN(n384) );
  XNOR2_X1 U452 ( .A(n385), .B(n384), .ZN(n386) );
  XOR2_X1 U453 ( .A(n386), .B(KEYINPUT90), .Z(n389) );
  XNOR2_X1 U454 ( .A(G22GAT), .B(n387), .ZN(n388) );
  XNOR2_X1 U455 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U456 ( .A(G78GAT), .B(KEYINPUT73), .Z(n391) );
  XNOR2_X1 U457 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n390) );
  XNOR2_X1 U458 ( .A(n391), .B(n390), .ZN(n437) );
  XOR2_X1 U459 ( .A(n437), .B(KEYINPUT23), .Z(n393) );
  NAND2_X1 U460 ( .A1(G228GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U461 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U462 ( .A(n395), .B(n394), .Z(n399) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n472) );
  XOR2_X1 U465 ( .A(n472), .B(KEYINPUT66), .Z(n400) );
  XNOR2_X1 U466 ( .A(KEYINPUT28), .B(n400), .ZN(n527) );
  NOR2_X1 U467 ( .A1(n525), .A2(n527), .ZN(n401) );
  NAND2_X1 U468 ( .A1(n528), .A2(n401), .ZN(n412) );
  NOR2_X1 U469 ( .A1(n520), .A2(n472), .ZN(n402) );
  XNOR2_X1 U470 ( .A(n402), .B(KEYINPUT26), .ZN(n565) );
  NAND2_X1 U471 ( .A1(n403), .A2(n565), .ZN(n408) );
  NAND2_X1 U472 ( .A1(n520), .A2(n518), .ZN(n404) );
  NAND2_X1 U473 ( .A1(n404), .A2(n472), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n405), .B(KEYINPUT25), .ZN(n406) );
  XOR2_X1 U475 ( .A(KEYINPUT98), .B(n406), .Z(n407) );
  NAND2_X1 U476 ( .A1(n408), .A2(n407), .ZN(n410) );
  NAND2_X1 U477 ( .A1(n410), .A2(n409), .ZN(n411) );
  NAND2_X1 U478 ( .A1(n412), .A2(n411), .ZN(n481) );
  NAND2_X1 U479 ( .A1(n479), .A2(n481), .ZN(n413) );
  NOR2_X1 U480 ( .A1(n578), .A2(n413), .ZN(n416) );
  XOR2_X1 U481 ( .A(n418), .B(n417), .Z(n420) );
  XNOR2_X1 U482 ( .A(G29GAT), .B(G50GAT), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n425) );
  XOR2_X1 U484 ( .A(n421), .B(KEYINPUT30), .Z(n423) );
  NAND2_X1 U485 ( .A1(G229GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U486 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U487 ( .A(n425), .B(n424), .Z(n433) );
  XOR2_X1 U488 ( .A(G113GAT), .B(G197GAT), .Z(n427) );
  XNOR2_X1 U489 ( .A(G36GAT), .B(G141GAT), .ZN(n426) );
  XNOR2_X1 U490 ( .A(n427), .B(n426), .ZN(n431) );
  XOR2_X1 U491 ( .A(KEYINPUT71), .B(KEYINPUT68), .Z(n429) );
  XNOR2_X1 U492 ( .A(KEYINPUT67), .B(KEYINPUT29), .ZN(n428) );
  XNOR2_X1 U493 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U494 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U495 ( .A(n433), .B(n432), .Z(n500) );
  XOR2_X1 U496 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n435) );
  NAND2_X1 U497 ( .A1(G230GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U498 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U499 ( .A(n436), .B(KEYINPUT32), .Z(n440) );
  XNOR2_X1 U500 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n441), .B(KEYINPUT72), .ZN(n446) );
  XOR2_X1 U503 ( .A(G148GAT), .B(n442), .Z(n444) );
  XNOR2_X1 U504 ( .A(n448), .B(n447), .ZN(n570) );
  OR2_X1 U505 ( .A1(n500), .A2(n570), .ZN(n483) );
  NOR2_X1 U506 ( .A1(n514), .A2(n483), .ZN(n449) );
  NAND2_X1 U507 ( .A1(n498), .A2(n520), .ZN(n453) );
  XOR2_X1 U508 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n451) );
  INV_X1 U509 ( .A(n500), .ZN(n566) );
  NOR2_X1 U510 ( .A1(n578), .A2(n479), .ZN(n454) );
  XOR2_X1 U511 ( .A(KEYINPUT45), .B(n454), .Z(n455) );
  NOR2_X1 U512 ( .A1(n455), .A2(n570), .ZN(n456) );
  XOR2_X1 U513 ( .A(KEYINPUT114), .B(n456), .Z(n457) );
  NOR2_X1 U514 ( .A1(n566), .A2(n457), .ZN(n466) );
  NAND2_X1 U515 ( .A1(n566), .A2(n559), .ZN(n459) );
  XOR2_X1 U516 ( .A(KEYINPUT112), .B(KEYINPUT46), .Z(n458) );
  XNOR2_X1 U517 ( .A(n459), .B(n458), .ZN(n460) );
  NOR2_X1 U518 ( .A1(n460), .A2(n575), .ZN(n461) );
  XNOR2_X1 U519 ( .A(n461), .B(KEYINPUT113), .ZN(n463) );
  BUF_X1 U520 ( .A(n462), .Z(n550) );
  NOR2_X1 U521 ( .A1(n463), .A2(n550), .ZN(n464) );
  XOR2_X1 U522 ( .A(n464), .B(KEYINPUT47), .Z(n465) );
  XNOR2_X1 U523 ( .A(n467), .B(KEYINPUT48), .ZN(n526) );
  XNOR2_X1 U524 ( .A(KEYINPUT123), .B(n518), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n526), .A2(n468), .ZN(n469) );
  XNOR2_X1 U526 ( .A(KEYINPUT54), .B(n469), .ZN(n470) );
  INV_X1 U527 ( .A(n470), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n515), .A2(n471), .ZN(n564) );
  AND2_X1 U529 ( .A1(n564), .A2(n472), .ZN(n473) );
  XNOR2_X1 U530 ( .A(n473), .B(KEYINPUT55), .ZN(n474) );
  NOR2_X2 U531 ( .A1(n528), .A2(n474), .ZN(n562) );
  NAND2_X1 U532 ( .A1(n562), .A2(n550), .ZN(n476) );
  XNOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT100), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n477), .B(KEYINPUT34), .ZN(n478) );
  XOR2_X1 U535 ( .A(KEYINPUT99), .B(n478), .Z(n485) );
  NOR2_X1 U536 ( .A1(n550), .A2(n479), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n480), .B(KEYINPUT16), .ZN(n482) );
  NAND2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n501) );
  NOR2_X1 U539 ( .A1(n483), .A2(n501), .ZN(n491) );
  NAND2_X1 U540 ( .A1(n491), .A2(n515), .ZN(n484) );
  XNOR2_X1 U541 ( .A(n485), .B(n484), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n518), .A2(n491), .ZN(n486) );
  XNOR2_X1 U543 ( .A(n486), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(KEYINPUT35), .B(KEYINPUT102), .Z(n488) );
  NAND2_X1 U545 ( .A1(n491), .A2(n520), .ZN(n487) );
  XNOR2_X1 U546 ( .A(n488), .B(n487), .ZN(n490) );
  XOR2_X1 U547 ( .A(G15GAT), .B(KEYINPUT101), .Z(n489) );
  XNOR2_X1 U548 ( .A(n490), .B(n489), .ZN(G1326GAT) );
  NAND2_X1 U549 ( .A1(n527), .A2(n491), .ZN(n492) );
  XNOR2_X1 U550 ( .A(n492), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U551 ( .A(G29GAT), .B(KEYINPUT104), .Z(n494) );
  NAND2_X1 U552 ( .A1(n515), .A2(n498), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT39), .B(n495), .ZN(G1328GAT) );
  XOR2_X1 U555 ( .A(G36GAT), .B(KEYINPUT105), .Z(n497) );
  NAND2_X1 U556 ( .A1(n498), .A2(n518), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n497), .B(n496), .ZN(G1329GAT) );
  NAND2_X1 U558 ( .A1(n498), .A2(n527), .ZN(n499) );
  XNOR2_X1 U559 ( .A(n499), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U560 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n503) );
  NAND2_X1 U561 ( .A1(n500), .A2(n559), .ZN(n513) );
  NOR2_X1 U562 ( .A1(n513), .A2(n501), .ZN(n509) );
  NAND2_X1 U563 ( .A1(n515), .A2(n509), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1332GAT) );
  XOR2_X1 U565 ( .A(G64GAT), .B(KEYINPUT107), .Z(n505) );
  NAND2_X1 U566 ( .A1(n509), .A2(n518), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n505), .B(n504), .ZN(G1333GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n507) );
  NAND2_X1 U569 ( .A1(n509), .A2(n520), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U571 ( .A(G71GAT), .B(n508), .ZN(G1334GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U573 ( .A1(n509), .A2(n527), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(n512), .ZN(G1335GAT) );
  XOR2_X1 U576 ( .A(G85GAT), .B(KEYINPUT111), .Z(n517) );
  NOR2_X1 U577 ( .A1(n514), .A2(n513), .ZN(n522) );
  NAND2_X1 U578 ( .A1(n522), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U580 ( .A1(n518), .A2(n522), .ZN(n519) );
  XNOR2_X1 U581 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U582 ( .A1(n520), .A2(n522), .ZN(n521) );
  XNOR2_X1 U583 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U584 ( .A1(n527), .A2(n522), .ZN(n523) );
  XNOR2_X1 U585 ( .A(n523), .B(KEYINPUT44), .ZN(n524) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(n524), .ZN(G1339GAT) );
  NOR2_X1 U587 ( .A1(n526), .A2(n525), .ZN(n542) );
  NOR2_X1 U588 ( .A1(n528), .A2(n527), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n542), .A2(n529), .ZN(n530) );
  XNOR2_X1 U590 ( .A(KEYINPUT115), .B(n530), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n539), .A2(n566), .ZN(n531) );
  XNOR2_X1 U592 ( .A(n531), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n533) );
  NAND2_X1 U594 ( .A1(n539), .A2(n559), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(n535) );
  XOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT116), .Z(n534) );
  XNOR2_X1 U597 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  XOR2_X1 U598 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n537) );
  NAND2_X1 U599 ( .A1(n539), .A2(n575), .ZN(n536) );
  XNOR2_X1 U600 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U601 ( .A(G127GAT), .B(n538), .Z(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n541) );
  NAND2_X1 U603 ( .A1(n539), .A2(n550), .ZN(n540) );
  XNOR2_X1 U604 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  AND2_X1 U605 ( .A1(n542), .A2(n565), .ZN(n551) );
  NAND2_X1 U606 ( .A1(n566), .A2(n551), .ZN(n543) );
  XOR2_X1 U607 ( .A(KEYINPUT119), .B(n543), .Z(n544) );
  XNOR2_X1 U608 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XNOR2_X1 U609 ( .A(G148GAT), .B(KEYINPUT120), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U611 ( .A1(n551), .A2(n559), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n575), .A2(n551), .ZN(n549) );
  XNOR2_X1 U615 ( .A(n549), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U616 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n553) );
  NAND2_X1 U617 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n554), .ZN(G1347GAT) );
  NAND2_X1 U620 ( .A1(n562), .A2(n566), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U622 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n557) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(n558) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(n558), .Z(n561) );
  NAND2_X1 U626 ( .A1(n559), .A2(n562), .ZN(n560) );
  XNOR2_X1 U627 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U628 ( .A1(n575), .A2(n562), .ZN(n563) );
  XNOR2_X1 U629 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n568) );
  NAND2_X1 U631 ( .A1(n564), .A2(n565), .ZN(n577) );
  INV_X1 U632 ( .A(n577), .ZN(n574) );
  NAND2_X1 U633 ( .A1(n574), .A2(n566), .ZN(n567) );
  XNOR2_X1 U634 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n572) );
  NAND2_X1 U637 ( .A1(n574), .A2(n570), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n573), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n576), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U642 ( .A1(n578), .A2(n577), .ZN(n580) );
  XNOR2_X1 U643 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G218GAT), .B(n581), .ZN(G1355GAT) );
endmodule

