

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746;

  AND2_X2 U368 ( .A1(n352), .A2(n359), .ZN(n356) );
  INV_X1 U369 ( .A(G953), .ZN(n734) );
  AND2_X2 U370 ( .A1(n390), .A2(n401), .ZN(n353) );
  INV_X2 U371 ( .A(KEYINPUT4), .ZN(n408) );
  XOR2_X2 U372 ( .A(KEYINPUT38), .B(n564), .Z(n674) );
  XNOR2_X2 U373 ( .A(n507), .B(n348), .ZN(n447) );
  XNOR2_X1 U374 ( .A(G119), .B(G113), .ZN(n370) );
  NOR2_X1 U375 ( .A1(n525), .A2(n403), .ZN(n526) );
  OR2_X2 U376 ( .A1(n540), .A2(n657), .ZN(n660) );
  XNOR2_X1 U377 ( .A(n605), .B(n604), .ZN(n606) );
  XNOR2_X1 U378 ( .A(n436), .B(n435), .ZN(n540) );
  NOR2_X1 U379 ( .A1(n611), .A2(G902), .ZN(n418) );
  XNOR2_X1 U380 ( .A(n621), .B(KEYINPUT59), .ZN(n622) );
  XNOR2_X1 U381 ( .A(n421), .B(n420), .ZN(n493) );
  XNOR2_X1 U382 ( .A(n370), .B(n369), .ZN(n460) );
  NAND2_X1 U383 ( .A1(n493), .A2(G221), .ZN(n382) );
  XNOR2_X1 U384 ( .A(n555), .B(n347), .ZN(n439) );
  XNOR2_X1 U385 ( .A(n447), .B(n388), .ZN(n546) );
  INV_X1 U386 ( .A(KEYINPUT90), .ZN(n388) );
  NOR2_X1 U387 ( .A1(n570), .A2(n569), .ZN(n571) );
  INV_X1 U388 ( .A(KEYINPUT46), .ZN(n379) );
  XNOR2_X1 U389 ( .A(G116), .B(G131), .ZN(n410) );
  NAND2_X1 U390 ( .A1(n360), .A2(n401), .ZN(n359) );
  AND2_X1 U391 ( .A1(n402), .A2(KEYINPUT84), .ZN(n363) );
  NOR2_X1 U392 ( .A1(n533), .A2(KEYINPUT44), .ZN(n365) );
  XNOR2_X1 U393 ( .A(G137), .B(G128), .ZN(n422) );
  XNOR2_X1 U394 ( .A(n428), .B(n419), .ZN(n385) );
  XNOR2_X1 U395 ( .A(KEYINPUT94), .B(KEYINPUT24), .ZN(n419) );
  XOR2_X1 U396 ( .A(KEYINPUT8), .B(KEYINPUT70), .Z(n421) );
  NOR2_X1 U397 ( .A1(G953), .A2(G237), .ZN(n479) );
  XOR2_X1 U398 ( .A(G104), .B(G122), .Z(n484) );
  XNOR2_X1 U399 ( .A(n409), .B(G125), .ZN(n450) );
  XNOR2_X1 U400 ( .A(G140), .B(G131), .ZN(n485) );
  NOR2_X1 U401 ( .A1(G902), .A2(n710), .ZN(n436) );
  NOR2_X1 U402 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U403 ( .A(n584), .B(KEYINPUT112), .ZN(n544) );
  INV_X1 U404 ( .A(KEYINPUT79), .ZN(n374) );
  BUF_X1 U405 ( .A(n563), .Z(n564) );
  AND2_X1 U406 ( .A1(n389), .A2(n656), .ZN(n406) );
  INV_X1 U407 ( .A(n439), .ZN(n403) );
  XNOR2_X1 U408 ( .A(n518), .B(n517), .ZN(n528) );
  INV_X1 U409 ( .A(n447), .ZN(n389) );
  NAND2_X1 U410 ( .A1(n389), .A2(n660), .ZN(n661) );
  INV_X1 U411 ( .A(G237), .ZN(n464) );
  XNOR2_X1 U412 ( .A(n354), .B(n377), .ZN(n596) );
  INV_X1 U413 ( .A(KEYINPUT48), .ZN(n377) );
  AND2_X1 U414 ( .A1(n571), .A2(n572), .ZN(n380) );
  NAND2_X1 U415 ( .A1(G234), .A2(G237), .ZN(n469) );
  OR2_X1 U416 ( .A1(n628), .A2(n397), .ZN(n396) );
  NAND2_X1 U417 ( .A1(n398), .A2(n490), .ZN(n397) );
  OR2_X1 U418 ( .A1(n677), .A2(n657), .ZN(n514) );
  XNOR2_X1 U419 ( .A(n375), .B(n440), .ZN(n416) );
  NAND2_X1 U420 ( .A1(n367), .A2(n364), .ZN(n534) );
  NAND2_X1 U421 ( .A1(n366), .A2(n365), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n383), .B(n381), .ZN(n710) );
  XNOR2_X1 U423 ( .A(n382), .B(n424), .ZN(n381) );
  XNOR2_X1 U424 ( .A(n385), .B(n728), .ZN(n383) );
  XOR2_X1 U425 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n481) );
  XNOR2_X1 U426 ( .A(G143), .B(G113), .ZN(n483) );
  XNOR2_X1 U427 ( .A(n450), .B(n384), .ZN(n728) );
  XNOR2_X1 U428 ( .A(KEYINPUT10), .B(KEYINPUT71), .ZN(n384) );
  XNOR2_X1 U429 ( .A(G104), .B(G110), .ZN(n441) );
  NOR2_X1 U430 ( .A1(n677), .A2(n679), .ZN(n579) );
  NOR2_X1 U431 ( .A1(n505), .A2(n389), .ZN(n667) );
  NOR2_X1 U432 ( .A1(n562), .A2(n660), .ZN(n573) );
  NOR2_X1 U433 ( .A1(n580), .A2(n404), .ZN(n552) );
  XNOR2_X1 U434 ( .A(n492), .B(n491), .ZN(n513) );
  NAND2_X1 U435 ( .A1(n585), .A2(n389), .ZN(n587) );
  XNOR2_X1 U436 ( .A(n545), .B(n357), .ZN(n547) );
  INV_X1 U437 ( .A(KEYINPUT36), .ZN(n357) );
  XNOR2_X1 U438 ( .A(n371), .B(n350), .ZN(n743) );
  NAND2_X1 U439 ( .A1(n406), .A2(n548), .ZN(n405) );
  NAND2_X1 U440 ( .A1(n519), .A2(n389), .ZN(n520) );
  NOR2_X1 U441 ( .A1(n656), .A2(n403), .ZN(n519) );
  INV_X1 U442 ( .A(G146), .ZN(n409) );
  AND2_X1 U443 ( .A1(n400), .A2(n399), .ZN(n346) );
  XOR2_X1 U444 ( .A(KEYINPUT101), .B(KEYINPUT6), .Z(n347) );
  XOR2_X1 U445 ( .A(KEYINPUT66), .B(KEYINPUT1), .Z(n348) );
  AND2_X1 U446 ( .A1(n561), .A2(n559), .ZN(n349) );
  XOR2_X1 U447 ( .A(n527), .B(KEYINPUT32), .Z(n350) );
  XNOR2_X1 U448 ( .A(n445), .B(n730), .ZN(n628) );
  INV_X1 U449 ( .A(KEYINPUT84), .ZN(n401) );
  INV_X1 U450 ( .A(n627), .ZN(n709) );
  NAND2_X1 U451 ( .A1(n716), .A2(n351), .ZN(n697) );
  XNOR2_X1 U452 ( .A(n592), .B(n593), .ZN(n351) );
  XNOR2_X2 U453 ( .A(n534), .B(KEYINPUT45), .ZN(n716) );
  NAND2_X1 U454 ( .A1(n378), .A2(n380), .ZN(n354) );
  NAND2_X1 U455 ( .A1(n353), .A2(n392), .ZN(n352) );
  NAND2_X1 U456 ( .A1(n555), .A2(n673), .ZN(n557) );
  XNOR2_X2 U457 ( .A(n418), .B(n417), .ZN(n555) );
  NAND2_X1 U458 ( .A1(n742), .A2(n746), .ZN(n358) );
  XNOR2_X1 U459 ( .A(n578), .B(KEYINPUT109), .ZN(n742) );
  NAND2_X1 U460 ( .A1(n560), .A2(n349), .ZN(n562) );
  NAND2_X1 U461 ( .A1(n363), .A2(n362), .ZN(n361) );
  NAND2_X2 U462 ( .A1(n346), .A2(n396), .ZN(n507) );
  XNOR2_X1 U463 ( .A(n355), .B(n489), .ZN(n621) );
  XNOR2_X1 U464 ( .A(n488), .B(n728), .ZN(n355) );
  NAND2_X1 U465 ( .A1(n743), .A2(n744), .ZN(n531) );
  NOR2_X1 U466 ( .A1(n528), .A2(n405), .ZN(n530) );
  NAND2_X1 U467 ( .A1(n532), .A2(KEYINPUT44), .ZN(n376) );
  XNOR2_X1 U468 ( .A(n386), .B(KEYINPUT35), .ZN(n532) );
  NAND2_X1 U469 ( .A1(n387), .A2(n503), .ZN(n386) );
  XNOR2_X1 U470 ( .A(n478), .B(n477), .ZN(n387) );
  NAND2_X1 U471 ( .A1(n356), .A2(n361), .ZN(n367) );
  NOR2_X1 U472 ( .A1(n706), .A2(G902), .ZN(n502) );
  XNOR2_X1 U473 ( .A(n501), .B(n500), .ZN(n706) );
  NAND2_X1 U474 ( .A1(n542), .A2(n403), .ZN(n584) );
  NAND2_X1 U475 ( .A1(n516), .A2(n672), .ZN(n478) );
  XNOR2_X2 U476 ( .A(n368), .B(n476), .ZN(n516) );
  XNOR2_X1 U477 ( .A(n358), .B(n379), .ZN(n378) );
  NOR2_X1 U478 ( .A1(n439), .A2(n660), .ZN(n448) );
  XNOR2_X1 U479 ( .A(n449), .B(KEYINPUT33), .ZN(n672) );
  INV_X1 U480 ( .A(n402), .ZN(n360) );
  NAND2_X1 U481 ( .A1(n392), .A2(n390), .ZN(n362) );
  INV_X1 U482 ( .A(n531), .ZN(n366) );
  NAND2_X1 U483 ( .A1(n475), .A2(n407), .ZN(n368) );
  XNOR2_X2 U484 ( .A(n543), .B(KEYINPUT19), .ZN(n475) );
  NAND2_X2 U485 ( .A1(n563), .A2(n673), .ZN(n543) );
  XNOR2_X2 U486 ( .A(KEYINPUT74), .B(KEYINPUT3), .ZN(n369) );
  NAND2_X1 U487 ( .A1(n373), .A2(n372), .ZN(n371) );
  INV_X1 U488 ( .A(n528), .ZN(n372) );
  XNOR2_X1 U489 ( .A(n526), .B(n374), .ZN(n373) );
  XNOR2_X1 U490 ( .A(n375), .B(n444), .ZN(n445) );
  XNOR2_X2 U491 ( .A(n453), .B(G146), .ZN(n375) );
  XNOR2_X2 U492 ( .A(n376), .B(KEYINPUT86), .ZN(n395) );
  NAND2_X1 U493 ( .A1(n596), .A2(n591), .ZN(n592) );
  NAND2_X1 U494 ( .A1(n395), .A2(n391), .ZN(n390) );
  NOR2_X1 U495 ( .A1(n522), .A2(KEYINPUT85), .ZN(n391) );
  NAND2_X1 U496 ( .A1(n393), .A2(KEYINPUT85), .ZN(n392) );
  NAND2_X1 U497 ( .A1(n395), .A2(n394), .ZN(n393) );
  INV_X1 U498 ( .A(n522), .ZN(n394) );
  NAND2_X1 U499 ( .A1(n628), .A2(n446), .ZN(n400) );
  INV_X1 U500 ( .A(n446), .ZN(n398) );
  NAND2_X1 U501 ( .A1(n446), .A2(G902), .ZN(n399) );
  NAND2_X1 U502 ( .A1(n531), .A2(KEYINPUT44), .ZN(n402) );
  XNOR2_X2 U503 ( .A(n440), .B(n485), .ZN(n730) );
  XNOR2_X2 U504 ( .A(n499), .B(G137), .ZN(n440) );
  XNOR2_X2 U505 ( .A(n451), .B(G134), .ZN(n499) );
  XNOR2_X2 U506 ( .A(G143), .B(G128), .ZN(n451) );
  INV_X1 U507 ( .A(n475), .ZN(n404) );
  OR2_X1 U508 ( .A1(n538), .A2(n474), .ZN(n407) );
  XNOR2_X1 U509 ( .A(KEYINPUT107), .B(KEYINPUT30), .ZN(n556) );
  INV_X1 U510 ( .A(n427), .ZN(n428) );
  XNOR2_X1 U511 ( .A(n557), .B(n556), .ZN(n560) );
  BUF_X1 U512 ( .A(n602), .Z(n605) );
  INV_X1 U513 ( .A(KEYINPUT78), .ZN(n527) );
  BUF_X1 U514 ( .A(n555), .Z(n663) );
  INV_X1 U515 ( .A(n715), .ZN(n617) );
  INV_X1 U516 ( .A(KEYINPUT104), .ZN(n529) );
  XNOR2_X2 U517 ( .A(n408), .B(KEYINPUT69), .ZN(n732) );
  XNOR2_X2 U518 ( .A(n732), .B(G101), .ZN(n453) );
  XOR2_X1 U519 ( .A(KEYINPUT98), .B(KEYINPUT5), .Z(n411) );
  XNOR2_X1 U520 ( .A(n411), .B(n410), .ZN(n413) );
  NAND2_X1 U521 ( .A1(n479), .A2(G210), .ZN(n412) );
  XNOR2_X1 U522 ( .A(n413), .B(n412), .ZN(n414) );
  XOR2_X1 U523 ( .A(n414), .B(n460), .Z(n415) );
  XNOR2_X1 U524 ( .A(n416), .B(n415), .ZN(n611) );
  XNOR2_X1 U525 ( .A(G472), .B(KEYINPUT75), .ZN(n417) );
  NAND2_X1 U526 ( .A1(G234), .A2(n734), .ZN(n420) );
  XOR2_X1 U527 ( .A(G110), .B(G119), .Z(n423) );
  XNOR2_X1 U528 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U529 ( .A(KEYINPUT23), .B(KEYINPUT76), .Z(n426) );
  XNOR2_X1 U530 ( .A(G140), .B(KEYINPUT95), .ZN(n425) );
  XNOR2_X1 U531 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U532 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n434) );
  INV_X1 U533 ( .A(KEYINPUT15), .ZN(n429) );
  XNOR2_X1 U534 ( .A(n429), .B(G902), .ZN(n594) );
  INV_X1 U535 ( .A(n594), .ZN(n430) );
  NAND2_X1 U536 ( .A1(n430), .A2(G234), .ZN(n432) );
  XNOR2_X1 U537 ( .A(KEYINPUT96), .B(KEYINPUT20), .ZN(n431) );
  XNOR2_X1 U538 ( .A(n432), .B(n431), .ZN(n437) );
  NAND2_X1 U539 ( .A1(G217), .A2(n437), .ZN(n433) );
  XOR2_X1 U540 ( .A(n434), .B(n433), .Z(n435) );
  NAND2_X1 U541 ( .A1(n437), .A2(G221), .ZN(n438) );
  XNOR2_X1 U542 ( .A(n438), .B(KEYINPUT21), .ZN(n657) );
  XNOR2_X1 U543 ( .A(n441), .B(G107), .ZN(n461) );
  NAND2_X1 U544 ( .A1(n734), .A2(G227), .ZN(n442) );
  XNOR2_X1 U545 ( .A(n442), .B(KEYINPUT77), .ZN(n443) );
  XNOR2_X1 U546 ( .A(n461), .B(n443), .ZN(n444) );
  XNOR2_X1 U547 ( .A(KEYINPUT73), .B(G469), .ZN(n446) );
  NAND2_X1 U548 ( .A1(n448), .A2(n447), .ZN(n449) );
  XNOR2_X1 U549 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U550 ( .A(n453), .B(n452), .ZN(n458) );
  XOR2_X1 U551 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n456) );
  NAND2_X1 U552 ( .A1(G224), .A2(n734), .ZN(n454) );
  XNOR2_X1 U553 ( .A(n454), .B(KEYINPUT88), .ZN(n455) );
  XNOR2_X1 U554 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U555 ( .A(n458), .B(n457), .ZN(n463) );
  XNOR2_X2 U556 ( .A(G122), .B(G116), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n497), .B(KEYINPUT16), .ZN(n459) );
  XNOR2_X1 U558 ( .A(n460), .B(n459), .ZN(n462) );
  XNOR2_X1 U559 ( .A(n462), .B(n461), .ZN(n722) );
  XNOR2_X1 U560 ( .A(n463), .B(n722), .ZN(n602) );
  OR2_X2 U561 ( .A1(n602), .A2(n594), .ZN(n467) );
  INV_X1 U562 ( .A(G902), .ZN(n490) );
  NAND2_X1 U563 ( .A1(n490), .A2(n464), .ZN(n468) );
  NAND2_X1 U564 ( .A1(n468), .A2(G210), .ZN(n465) );
  XNOR2_X1 U565 ( .A(n465), .B(KEYINPUT91), .ZN(n466) );
  XNOR2_X2 U566 ( .A(n467), .B(n466), .ZN(n563) );
  NAND2_X1 U567 ( .A1(n468), .A2(G214), .ZN(n673) );
  XNOR2_X1 U568 ( .A(n469), .B(KEYINPUT92), .ZN(n470) );
  XNOR2_X1 U569 ( .A(KEYINPUT14), .B(n470), .ZN(n472) );
  NAND2_X1 U570 ( .A1(n472), .A2(G952), .ZN(n471) );
  XOR2_X1 U571 ( .A(KEYINPUT93), .B(n471), .Z(n689) );
  NOR2_X1 U572 ( .A1(n689), .A2(G953), .ZN(n538) );
  AND2_X1 U573 ( .A1(n472), .A2(G953), .ZN(n473) );
  NAND2_X1 U574 ( .A1(G902), .A2(n473), .ZN(n535) );
  NOR2_X1 U575 ( .A1(n535), .A2(G898), .ZN(n474) );
  XNOR2_X1 U576 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n476) );
  INV_X1 U577 ( .A(KEYINPUT34), .ZN(n477) );
  NAND2_X1 U578 ( .A1(G214), .A2(n479), .ZN(n480) );
  XNOR2_X1 U579 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U580 ( .A(KEYINPUT11), .B(n482), .ZN(n489) );
  XNOR2_X1 U581 ( .A(n484), .B(n483), .ZN(n487) );
  INV_X1 U582 ( .A(n485), .ZN(n486) );
  XNOR2_X1 U583 ( .A(n487), .B(n486), .ZN(n488) );
  NAND2_X1 U584 ( .A1(n621), .A2(n490), .ZN(n492) );
  XNOR2_X1 U585 ( .A(KEYINPUT13), .B(G475), .ZN(n491) );
  XOR2_X1 U586 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n495) );
  NAND2_X1 U587 ( .A1(G217), .A2(n493), .ZN(n494) );
  XNOR2_X1 U588 ( .A(n495), .B(n494), .ZN(n501) );
  XOR2_X1 U589 ( .A(KEYINPUT100), .B(G107), .Z(n496) );
  XNOR2_X1 U590 ( .A(n497), .B(n496), .ZN(n498) );
  XNOR2_X1 U591 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U592 ( .A(G478), .B(n502), .ZN(n512) );
  OR2_X1 U593 ( .A1(n513), .A2(n512), .ZN(n566) );
  INV_X1 U594 ( .A(n566), .ZN(n503) );
  INV_X1 U595 ( .A(n660), .ZN(n504) );
  NAND2_X1 U596 ( .A1(n504), .A2(n663), .ZN(n505) );
  NAND2_X1 U597 ( .A1(n667), .A2(n516), .ZN(n506) );
  XOR2_X1 U598 ( .A(KEYINPUT31), .B(n506), .Z(n647) );
  INV_X1 U599 ( .A(n663), .ZN(n548) );
  INV_X1 U600 ( .A(n507), .ZN(n561) );
  NAND2_X1 U601 ( .A1(n548), .A2(n561), .ZN(n508) );
  NOR2_X1 U602 ( .A1(n660), .A2(n508), .ZN(n509) );
  NAND2_X1 U603 ( .A1(n509), .A2(n516), .ZN(n638) );
  NAND2_X1 U604 ( .A1(n647), .A2(n638), .ZN(n511) );
  INV_X1 U605 ( .A(n512), .ZN(n510) );
  NAND2_X1 U606 ( .A1(n513), .A2(n510), .ZN(n648) );
  OR2_X1 U607 ( .A1(n513), .A2(n510), .ZN(n645) );
  NAND2_X1 U608 ( .A1(n648), .A2(n645), .ZN(n678) );
  NAND2_X1 U609 ( .A1(n511), .A2(n678), .ZN(n521) );
  NAND2_X1 U610 ( .A1(n513), .A2(n512), .ZN(n677) );
  XOR2_X1 U611 ( .A(KEYINPUT102), .B(n514), .Z(n515) );
  NAND2_X1 U612 ( .A1(n516), .A2(n515), .ZN(n518) );
  XOR2_X1 U613 ( .A(KEYINPUT22), .B(KEYINPUT65), .Z(n517) );
  INV_X1 U614 ( .A(n540), .ZN(n523) );
  INV_X1 U615 ( .A(n523), .ZN(n656) );
  OR2_X1 U616 ( .A1(n528), .A2(n520), .ZN(n633) );
  NAND2_X1 U617 ( .A1(n521), .A2(n633), .ZN(n522) );
  NOR2_X1 U618 ( .A1(n546), .A2(n523), .ZN(n524) );
  XNOR2_X1 U619 ( .A(n524), .B(KEYINPUT103), .ZN(n525) );
  XNOR2_X1 U620 ( .A(n530), .B(n529), .ZN(n744) );
  BUF_X1 U621 ( .A(n532), .Z(n533) );
  INV_X1 U622 ( .A(KEYINPUT82), .ZN(n593) );
  NOR2_X1 U623 ( .A1(G900), .A2(n535), .ZN(n536) );
  XOR2_X1 U624 ( .A(KEYINPUT105), .B(n536), .Z(n537) );
  NOR2_X1 U625 ( .A1(n538), .A2(n537), .ZN(n558) );
  NOR2_X1 U626 ( .A1(n558), .A2(n657), .ZN(n539) );
  NAND2_X1 U627 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U628 ( .A(KEYINPUT72), .B(n541), .ZN(n549) );
  NOR2_X1 U629 ( .A1(n549), .A2(n645), .ZN(n542) );
  NOR2_X1 U630 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U631 ( .A1(n547), .A2(n546), .ZN(n652) );
  XNOR2_X1 U632 ( .A(KEYINPUT83), .B(n652), .ZN(n572) );
  XNOR2_X1 U633 ( .A(KEYINPUT28), .B(n550), .ZN(n551) );
  NAND2_X1 U634 ( .A1(n551), .A2(n561), .ZN(n580) );
  INV_X1 U635 ( .A(n645), .ZN(n575) );
  NAND2_X1 U636 ( .A1(n552), .A2(n575), .ZN(n644) );
  INV_X1 U637 ( .A(n648), .ZN(n590) );
  NAND2_X1 U638 ( .A1(n552), .A2(n590), .ZN(n641) );
  NAND2_X1 U639 ( .A1(n644), .A2(n641), .ZN(n553) );
  NAND2_X1 U640 ( .A1(n553), .A2(KEYINPUT68), .ZN(n554) );
  XNOR2_X1 U641 ( .A(n554), .B(KEYINPUT47), .ZN(n570) );
  INV_X1 U642 ( .A(n558), .ZN(n559) );
  INV_X1 U643 ( .A(n564), .ZN(n565) );
  NOR2_X1 U644 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U645 ( .A1(n573), .A2(n567), .ZN(n568) );
  XNOR2_X1 U646 ( .A(KEYINPUT108), .B(n568), .ZN(n745) );
  XNOR2_X1 U647 ( .A(KEYINPUT81), .B(n745), .ZN(n569) );
  NAND2_X1 U648 ( .A1(n573), .A2(n674), .ZN(n574) );
  XNOR2_X1 U649 ( .A(n574), .B(KEYINPUT39), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n589), .A2(n575), .ZN(n577) );
  XOR2_X1 U651 ( .A(KEYINPUT110), .B(KEYINPUT40), .Z(n576) );
  XNOR2_X1 U652 ( .A(n577), .B(n576), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n674), .A2(n673), .ZN(n679) );
  XNOR2_X1 U654 ( .A(n579), .B(KEYINPUT41), .ZN(n691) );
  NOR2_X1 U655 ( .A1(n691), .A2(n580), .ZN(n582) );
  XNOR2_X1 U656 ( .A(KEYINPUT111), .B(KEYINPUT42), .ZN(n581) );
  XNOR2_X1 U657 ( .A(n582), .B(n581), .ZN(n746) );
  INV_X1 U658 ( .A(n673), .ZN(n583) );
  NOR2_X1 U659 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U660 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n586) );
  XNOR2_X1 U661 ( .A(n587), .B(n586), .ZN(n588) );
  OR2_X1 U662 ( .A1(n588), .A2(n564), .ZN(n620) );
  NAND2_X1 U663 ( .A1(n589), .A2(n590), .ZN(n654) );
  AND2_X1 U664 ( .A1(n620), .A2(n654), .ZN(n595) );
  AND2_X1 U665 ( .A1(n595), .A2(KEYINPUT2), .ZN(n591) );
  AND2_X2 U666 ( .A1(n697), .A2(n594), .ZN(n599) );
  AND2_X1 U667 ( .A1(n596), .A2(n595), .ZN(n733) );
  NAND2_X1 U668 ( .A1(n716), .A2(n733), .ZN(n694) );
  INV_X1 U669 ( .A(KEYINPUT2), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n694), .A2(n597), .ZN(n598) );
  NAND2_X2 U671 ( .A1(n599), .A2(n598), .ZN(n601) );
  INV_X1 U672 ( .A(KEYINPUT64), .ZN(n600) );
  XNOR2_X2 U673 ( .A(n601), .B(n600), .ZN(n626) );
  NAND2_X1 U674 ( .A1(n626), .A2(G210), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT87), .B(KEYINPUT55), .Z(n603) );
  XOR2_X1 U676 ( .A(n603), .B(KEYINPUT54), .Z(n604) );
  XNOR2_X1 U677 ( .A(n607), .B(n606), .ZN(n609) );
  INV_X1 U678 ( .A(G952), .ZN(n608) );
  AND2_X1 U679 ( .A1(n608), .A2(G953), .ZN(n715) );
  NOR2_X2 U680 ( .A1(n609), .A2(n715), .ZN(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U682 ( .A1(n626), .A2(G472), .ZN(n615) );
  XNOR2_X1 U683 ( .A(KEYINPUT89), .B(KEYINPUT113), .ZN(n612) );
  XNOR2_X1 U684 ( .A(n612), .B(KEYINPUT62), .ZN(n613) );
  XNOR2_X1 U685 ( .A(n611), .B(n613), .ZN(n614) );
  XNOR2_X1 U686 ( .A(n615), .B(n614), .ZN(n616) );
  INV_X1 U687 ( .A(n616), .ZN(n618) );
  NAND2_X1 U688 ( .A1(n618), .A2(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(n619), .B(KEYINPUT63), .ZN(G57) );
  XNOR2_X1 U690 ( .A(n620), .B(G140), .ZN(G42) );
  XOR2_X1 U691 ( .A(G122), .B(n533), .Z(G24) );
  NAND2_X1 U692 ( .A1(n626), .A2(G475), .ZN(n623) );
  XNOR2_X1 U693 ( .A(n623), .B(n622), .ZN(n624) );
  NOR2_X2 U694 ( .A1(n624), .A2(n715), .ZN(n625) );
  XNOR2_X1 U695 ( .A(n625), .B(KEYINPUT60), .ZN(G60) );
  INV_X1 U696 ( .A(n626), .ZN(n627) );
  NAND2_X1 U697 ( .A1(n709), .A2(G469), .ZN(n631) );
  XOR2_X1 U698 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n629) );
  XNOR2_X1 U699 ( .A(n628), .B(n629), .ZN(n630) );
  XNOR2_X1 U700 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X1 U701 ( .A1(n632), .A2(n715), .ZN(G54) );
  INV_X1 U702 ( .A(n633), .ZN(n634) );
  XOR2_X1 U703 ( .A(G101), .B(n634), .Z(G3) );
  NOR2_X1 U704 ( .A1(n638), .A2(n645), .ZN(n635) );
  XOR2_X1 U705 ( .A(G104), .B(n635), .Z(G6) );
  XOR2_X1 U706 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  XNOR2_X1 U707 ( .A(G107), .B(KEYINPUT114), .ZN(n636) );
  XNOR2_X1 U708 ( .A(n637), .B(n636), .ZN(n640) );
  NOR2_X1 U709 ( .A1(n638), .A2(n648), .ZN(n639) );
  XOR2_X1 U710 ( .A(n640), .B(n639), .Z(G9) );
  XNOR2_X1 U711 ( .A(KEYINPUT29), .B(KEYINPUT115), .ZN(n642) );
  XNOR2_X1 U712 ( .A(n642), .B(n641), .ZN(n643) );
  XNOR2_X1 U713 ( .A(G128), .B(n643), .ZN(G30) );
  XNOR2_X1 U714 ( .A(G146), .B(n644), .ZN(G48) );
  NOR2_X1 U715 ( .A1(n645), .A2(n647), .ZN(n646) );
  XOR2_X1 U716 ( .A(G113), .B(n646), .Z(G15) );
  NOR2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n650) );
  XNOR2_X1 U718 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n649) );
  XNOR2_X1 U719 ( .A(n650), .B(n649), .ZN(n651) );
  XNOR2_X1 U720 ( .A(G116), .B(n651), .ZN(G18) );
  XNOR2_X1 U721 ( .A(G125), .B(n652), .ZN(n653) );
  XNOR2_X1 U722 ( .A(n653), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U723 ( .A(G134), .B(KEYINPUT118), .ZN(n655) );
  XNOR2_X1 U724 ( .A(n655), .B(n654), .ZN(G36) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U726 ( .A(n658), .B(KEYINPUT49), .ZN(n659) );
  XNOR2_X1 U727 ( .A(KEYINPUT119), .B(n659), .ZN(n666) );
  XNOR2_X1 U728 ( .A(KEYINPUT120), .B(KEYINPUT50), .ZN(n662) );
  XOR2_X1 U729 ( .A(n662), .B(n661), .Z(n664) );
  NOR2_X1 U730 ( .A1(n664), .A2(n663), .ZN(n665) );
  NAND2_X1 U731 ( .A1(n666), .A2(n665), .ZN(n669) );
  INV_X1 U732 ( .A(n667), .ZN(n668) );
  NAND2_X1 U733 ( .A1(n669), .A2(n668), .ZN(n670) );
  XNOR2_X1 U734 ( .A(KEYINPUT51), .B(n670), .ZN(n671) );
  NOR2_X1 U735 ( .A1(n671), .A2(n691), .ZN(n686) );
  INV_X1 U736 ( .A(n672), .ZN(n690) );
  NOR2_X1 U737 ( .A1(n674), .A2(n673), .ZN(n675) );
  XOR2_X1 U738 ( .A(KEYINPUT121), .B(n675), .Z(n676) );
  NOR2_X1 U739 ( .A1(n677), .A2(n676), .ZN(n683) );
  INV_X1 U740 ( .A(n678), .ZN(n680) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U742 ( .A(n681), .B(KEYINPUT122), .ZN(n682) );
  NOR2_X1 U743 ( .A1(n683), .A2(n682), .ZN(n684) );
  NOR2_X1 U744 ( .A1(n690), .A2(n684), .ZN(n685) );
  NOR2_X1 U745 ( .A1(n686), .A2(n685), .ZN(n687) );
  XNOR2_X1 U746 ( .A(n687), .B(KEYINPUT52), .ZN(n688) );
  NOR2_X1 U747 ( .A1(n689), .A2(n688), .ZN(n693) );
  NOR2_X1 U748 ( .A1(n691), .A2(n690), .ZN(n692) );
  OR2_X1 U749 ( .A1(n693), .A2(n692), .ZN(n702) );
  INV_X1 U750 ( .A(n694), .ZN(n696) );
  XNOR2_X1 U751 ( .A(KEYINPUT80), .B(KEYINPUT2), .ZN(n695) );
  NOR2_X1 U752 ( .A1(n696), .A2(n695), .ZN(n700) );
  BUF_X1 U753 ( .A(n697), .Z(n698) );
  INV_X1 U754 ( .A(n698), .ZN(n699) );
  NOR2_X1 U755 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U756 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U757 ( .A(n703), .B(KEYINPUT123), .ZN(n704) );
  NOR2_X1 U758 ( .A1(G953), .A2(n704), .ZN(n705) );
  XNOR2_X1 U759 ( .A(KEYINPUT53), .B(n705), .ZN(G75) );
  NAND2_X1 U760 ( .A1(n709), .A2(G478), .ZN(n707) );
  XNOR2_X1 U761 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U762 ( .A1(n715), .A2(n708), .ZN(G63) );
  NAND2_X1 U763 ( .A1(n709), .A2(G217), .ZN(n713) );
  BUF_X1 U764 ( .A(n710), .Z(n711) );
  XNOR2_X1 U765 ( .A(n711), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U766 ( .A(n713), .B(n712), .ZN(n714) );
  NOR2_X1 U767 ( .A1(n715), .A2(n714), .ZN(G66) );
  BUF_X1 U768 ( .A(n716), .Z(n717) );
  NAND2_X1 U769 ( .A1(n717), .A2(n734), .ZN(n721) );
  NAND2_X1 U770 ( .A1(G953), .A2(G224), .ZN(n718) );
  XNOR2_X1 U771 ( .A(KEYINPUT61), .B(n718), .ZN(n719) );
  NAND2_X1 U772 ( .A1(n719), .A2(G898), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n727) );
  XNOR2_X1 U774 ( .A(n722), .B(G101), .ZN(n724) );
  NOR2_X1 U775 ( .A1(G898), .A2(n734), .ZN(n723) );
  NOR2_X1 U776 ( .A1(n724), .A2(n723), .ZN(n725) );
  XOR2_X1 U777 ( .A(KEYINPUT125), .B(n725), .Z(n726) );
  XNOR2_X1 U778 ( .A(n727), .B(n726), .ZN(G69) );
  XNOR2_X1 U779 ( .A(n728), .B(KEYINPUT126), .ZN(n729) );
  XOR2_X1 U780 ( .A(n730), .B(n729), .Z(n731) );
  XOR2_X1 U781 ( .A(n732), .B(n731), .Z(n736) );
  XNOR2_X1 U782 ( .A(n733), .B(n736), .ZN(n735) );
  NAND2_X1 U783 ( .A1(n735), .A2(n734), .ZN(n741) );
  XOR2_X1 U784 ( .A(G227), .B(n736), .Z(n737) );
  NAND2_X1 U785 ( .A1(n737), .A2(G900), .ZN(n738) );
  NAND2_X1 U786 ( .A1(G953), .A2(n738), .ZN(n739) );
  XOR2_X1 U787 ( .A(KEYINPUT127), .B(n739), .Z(n740) );
  NAND2_X1 U788 ( .A1(n741), .A2(n740), .ZN(G72) );
  XNOR2_X1 U789 ( .A(G131), .B(n742), .ZN(G33) );
  XNOR2_X1 U790 ( .A(n743), .B(G119), .ZN(G21) );
  XNOR2_X1 U791 ( .A(n744), .B(G110), .ZN(G12) );
  XNOR2_X1 U792 ( .A(G143), .B(n745), .ZN(G45) );
  XNOR2_X1 U793 ( .A(G137), .B(n746), .ZN(G39) );
endmodule

