//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 0 0 0 1 1 1 1 0 1 1 0 1 0 0 1 0 0 0 1 0 1 0 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n623,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n864,
    new_n865, new_n866, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1238, new_n1239, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1249, new_n1250, new_n1251, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XNOR2_X1  g005(.A(KEYINPUT64), .B(G2066), .ZN(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT65), .B(G452), .ZN(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(KEYINPUT3), .ZN(new_n460));
  INV_X1    g035(.A(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2104), .ZN(new_n462));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND4_X1  g038(.A1(new_n460), .A2(new_n462), .A3(G137), .A4(new_n463), .ZN(new_n464));
  NOR2_X1   g039(.A1(new_n459), .A2(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(G101), .ZN(new_n466));
  AND3_X1   g041(.A1(new_n464), .A2(KEYINPUT67), .A3(new_n466), .ZN(new_n467));
  AOI21_X1  g042(.A(KEYINPUT67), .B1(new_n464), .B2(new_n466), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n460), .A2(new_n462), .A3(G125), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  NAND2_X1  g050(.A1(new_n460), .A2(new_n462), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n476), .A2(new_n463), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G124), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n476), .A2(G2105), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G136), .ZN(new_n480));
  OR2_X1    g055(.A1(G100), .A2(G2105), .ZN(new_n481));
  OAI211_X1 g056(.A(new_n481), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n482));
  NAND3_X1  g057(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(new_n483), .ZN(G162));
  NAND4_X1  g059(.A1(new_n460), .A2(new_n462), .A3(G138), .A4(new_n463), .ZN(new_n485));
  NAND2_X1  g060(.A1(new_n485), .A2(KEYINPUT4), .ZN(new_n486));
  XNOR2_X1  g061(.A(KEYINPUT3), .B(G2104), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n487), .A2(new_n488), .A3(G138), .A4(new_n463), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n486), .A2(new_n489), .ZN(new_n490));
  OR2_X1    g065(.A1(G102), .A2(G2105), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n491), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n492));
  NAND4_X1  g067(.A1(new_n460), .A2(new_n462), .A3(G126), .A4(G2105), .ZN(new_n493));
  AND2_X1   g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n490), .A2(KEYINPUT68), .A3(new_n494), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(G164));
  INV_X1    g074(.A(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT6), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  AND2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(G543), .ZN(new_n505));
  INV_X1    g080(.A(G50), .ZN(new_n506));
  INV_X1    g081(.A(G88), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT69), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT5), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n510), .A2(KEYINPUT69), .A3(G543), .ZN(new_n511));
  NAND4_X1  g086(.A1(new_n509), .A2(new_n511), .A3(new_n501), .A4(new_n503), .ZN(new_n512));
  OAI22_X1  g087(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n509), .A2(new_n511), .A3(G62), .ZN(new_n514));
  NAND2_X1  g089(.A1(G75), .A2(G543), .ZN(new_n515));
  AOI21_X1  g090(.A(new_n500), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NOR2_X1   g091(.A1(new_n513), .A2(new_n516), .ZN(G166));
  AND3_X1   g092(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT70), .ZN(new_n518));
  AOI21_X1  g093(.A(KEYINPUT70), .B1(new_n509), .B2(new_n511), .ZN(new_n519));
  NAND2_X1  g094(.A1(G63), .A2(G651), .ZN(new_n520));
  NOR3_X1   g095(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  NAND4_X1  g096(.A1(new_n501), .A2(new_n503), .A3(G51), .A4(G543), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n522), .B(new_n527), .C1(new_n512), .C2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n521), .A2(new_n529), .ZN(G168));
  INV_X1    g105(.A(G64), .ZN(new_n531));
  NOR3_X1   g106(.A1(new_n518), .A2(new_n519), .A3(new_n531), .ZN(new_n532));
  INV_X1    g107(.A(G77), .ZN(new_n533));
  INV_X1    g108(.A(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g110(.A(G651), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n512), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n501), .A2(new_n503), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n538), .A2(new_n534), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n537), .A2(G90), .B1(new_n539), .B2(G52), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n536), .A2(new_n540), .ZN(G301));
  INV_X1    g116(.A(G301), .ZN(G171));
  AOI22_X1  g117(.A1(new_n537), .A2(G81), .B1(new_n539), .B2(G43), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT70), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n510), .B1(KEYINPUT69), .B2(G543), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n508), .A2(KEYINPUT5), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n544), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n509), .A2(new_n511), .A3(KEYINPUT70), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n547), .A2(G56), .A3(new_n548), .ZN(new_n549));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n500), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  OAI21_X1  g127(.A(new_n543), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  AOI211_X1 g128(.A(KEYINPUT71), .B(new_n500), .C1(new_n549), .C2(new_n550), .ZN(new_n554));
  NOR2_X1   g129(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  INV_X1    g136(.A(KEYINPUT72), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n504), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n501), .A2(new_n503), .A3(G53), .A4(G543), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(KEYINPUT72), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(KEYINPUT9), .A3(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT9), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n564), .A2(KEYINPUT72), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n537), .A2(G91), .ZN(new_n569));
  NAND2_X1  g144(.A1(G78), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n509), .A2(new_n511), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n566), .A2(new_n568), .A3(new_n569), .A4(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  INV_X1    g151(.A(G166), .ZN(G303));
  NAND2_X1  g152(.A1(new_n537), .A2(G87), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n501), .A2(new_n503), .A3(G49), .A4(G543), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n579), .A2(KEYINPUT73), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(KEYINPUT73), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  INV_X1    g157(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n547), .A2(new_n548), .ZN(new_n584));
  INV_X1    g159(.A(G74), .ZN(new_n585));
  AOI21_X1  g160(.A(new_n500), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT74), .ZN(new_n588));
  NAND3_X1  g163(.A1(new_n583), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(KEYINPUT74), .B1(new_n582), .B2(new_n586), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(G288));
  NAND2_X1  g166(.A1(new_n537), .A2(G86), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G73), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G61), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n571), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n539), .B2(G48), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n537), .A2(KEYINPUT75), .A3(G86), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(G305));
  NOR2_X1   g175(.A1(new_n518), .A2(new_n519), .ZN(new_n601));
  AOI22_X1  g176(.A1(new_n601), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n602));
  NOR2_X1   g177(.A1(new_n602), .A2(new_n500), .ZN(new_n603));
  INV_X1    g178(.A(G47), .ZN(new_n604));
  INV_X1    g179(.A(G85), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n505), .A2(new_n604), .B1(new_n605), .B2(new_n512), .ZN(new_n606));
  NOR2_X1   g181(.A1(new_n603), .A2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(new_n607), .ZN(G290));
  NAND3_X1  g183(.A1(new_n537), .A2(KEYINPUT10), .A3(G92), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT10), .ZN(new_n610));
  INV_X1    g185(.A(G92), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n610), .B1(new_n512), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n509), .A2(new_n511), .A3(G66), .ZN(new_n614));
  NAND2_X1  g189(.A1(G79), .A2(G543), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n616), .A2(G651), .B1(new_n539), .B2(G54), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G868), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n620), .B1(G171), .B2(new_n619), .ZN(G284));
  XNOR2_X1  g196(.A(G284), .B(KEYINPUT76), .ZN(G321));
  NAND2_X1  g197(.A1(G299), .A2(new_n619), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n619), .B2(G168), .ZN(G297));
  OAI21_X1  g199(.A(new_n623), .B1(new_n619), .B2(G168), .ZN(G280));
  AND2_X1   g200(.A1(new_n613), .A2(new_n617), .ZN(new_n626));
  INV_X1    g201(.A(G559), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n626), .B1(new_n627), .B2(G860), .ZN(G148));
  NAND2_X1  g203(.A1(new_n626), .A2(new_n627), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n629), .A2(G868), .ZN(new_n630));
  OAI21_X1  g205(.A(new_n630), .B1(G868), .B2(new_n555), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT77), .Z(G323));
  XNOR2_X1  g207(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g208(.A1(new_n487), .A2(new_n465), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(KEYINPUT12), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT13), .ZN(new_n636));
  OR2_X1    g211(.A1(new_n636), .A2(G2100), .ZN(new_n637));
  AOI22_X1  g212(.A1(G123), .A2(new_n477), .B1(new_n479), .B2(G135), .ZN(new_n638));
  OAI21_X1  g213(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n639));
  INV_X1    g214(.A(G111), .ZN(new_n640));
  AOI22_X1  g215(.A1(new_n639), .A2(KEYINPUT78), .B1(new_n640), .B2(G2105), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n641), .B1(KEYINPUT78), .B2(new_n639), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(G2096), .Z(new_n644));
  NAND2_X1  g219(.A1(new_n636), .A2(G2100), .ZN(new_n645));
  NAND3_X1  g220(.A1(new_n637), .A2(new_n644), .A3(new_n645), .ZN(G156));
  XOR2_X1   g221(.A(G2427), .B(G2430), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n647), .B(KEYINPUT80), .ZN(new_n648));
  XNOR2_X1  g223(.A(KEYINPUT15), .B(G2435), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2438), .ZN(new_n650));
  NAND2_X1  g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n651), .A2(KEYINPUT14), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(KEYINPUT81), .ZN(new_n653));
  OR2_X1    g228(.A1(new_n648), .A2(new_n650), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(KEYINPUT16), .ZN(new_n656));
  INV_X1    g231(.A(KEYINPUT16), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n653), .A2(new_n657), .A3(new_n654), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G2451), .B(G2454), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  OR2_X1    g237(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(G1341), .B(G1348), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT82), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT79), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n659), .A2(new_n662), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n663), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n668), .A2(G14), .ZN(new_n669));
  AOI21_X1  g244(.A(new_n666), .B1(new_n663), .B2(new_n667), .ZN(new_n670));
  OR2_X1    g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G401));
  XNOR2_X1  g247(.A(G2067), .B(G2678), .ZN(new_n673));
  INV_X1    g248(.A(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G2072), .B(G2078), .Z(new_n675));
  XNOR2_X1  g250(.A(KEYINPUT83), .B(KEYINPUT17), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2084), .B(G2090), .Z(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n678), .B1(new_n674), .B2(new_n675), .ZN(new_n680));
  OAI21_X1  g255(.A(new_n674), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n677), .A2(new_n680), .ZN(new_n682));
  INV_X1    g257(.A(new_n675), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n683), .A2(new_n673), .A3(new_n678), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT18), .Z(new_n685));
  NAND3_X1  g260(.A1(new_n681), .A2(new_n682), .A3(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(G2100), .ZN(new_n687));
  XOR2_X1   g262(.A(KEYINPUT84), .B(G2096), .Z(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(G227));
  XNOR2_X1  g264(.A(G1991), .B(G1996), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT85), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G1971), .B(G1976), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT19), .ZN(new_n694));
  XOR2_X1   g269(.A(G1956), .B(G2474), .Z(new_n695));
  XOR2_X1   g270(.A(G1961), .B(G1966), .Z(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT20), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT20), .ZN(new_n700));
  NOR2_X1   g275(.A1(new_n695), .A2(new_n696), .ZN(new_n701));
  INV_X1    g276(.A(new_n701), .ZN(new_n702));
  OR2_X1    g277(.A1(new_n702), .A2(new_n694), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n702), .A2(new_n694), .A3(new_n697), .ZN(new_n704));
  NAND4_X1  g279(.A1(new_n699), .A2(new_n700), .A3(new_n703), .A4(new_n704), .ZN(new_n705));
  OR2_X1    g280(.A1(new_n705), .A2(KEYINPUT21), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n705), .A2(KEYINPUT21), .ZN(new_n707));
  AOI21_X1  g282(.A(KEYINPUT22), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n706), .A2(KEYINPUT22), .A3(new_n707), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n692), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(G1981), .B(G1986), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n709), .A2(new_n692), .A3(new_n710), .ZN(new_n714));
  AND3_X1   g289(.A1(new_n712), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(new_n713), .B1(new_n712), .B2(new_n714), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(G229));
  INV_X1    g293(.A(KEYINPUT30), .ZN(new_n719));
  AND2_X1   g294(.A1(new_n719), .A2(G28), .ZN(new_n720));
  INV_X1    g295(.A(G29), .ZN(new_n721));
  OAI21_X1  g296(.A(new_n721), .B1(new_n719), .B2(G28), .ZN(new_n722));
  AND2_X1   g297(.A1(KEYINPUT31), .A2(G11), .ZN(new_n723));
  NOR2_X1   g298(.A1(KEYINPUT31), .A2(G11), .ZN(new_n724));
  OAI22_X1  g299(.A1(new_n720), .A2(new_n722), .B1(new_n723), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g300(.A1(new_n643), .A2(new_n721), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT96), .Z(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G168), .B2(new_n728), .ZN(new_n730));
  AOI211_X1 g305(.A(new_n725), .B(new_n727), .C1(G1966), .C2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(G5), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(G171), .B2(new_n728), .ZN(new_n733));
  XNOR2_X1  g308(.A(new_n733), .B(KEYINPUT97), .ZN(new_n734));
  INV_X1    g309(.A(G1961), .ZN(new_n735));
  OAI221_X1 g310(.A(new_n731), .B1(G1966), .B2(new_n730), .C1(new_n734), .C2(new_n735), .ZN(new_n736));
  XOR2_X1   g311(.A(new_n736), .B(KEYINPUT98), .Z(new_n737));
  NAND2_X1  g312(.A1(new_n721), .A2(G26), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n477), .A2(G128), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n479), .A2(G140), .ZN(new_n740));
  OR2_X1    g315(.A1(G104), .A2(G2105), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n741), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n739), .A2(new_n740), .A3(new_n742), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n738), .B1(new_n744), .B2(new_n721), .ZN(new_n745));
  MUX2_X1   g320(.A(new_n738), .B(new_n745), .S(KEYINPUT28), .Z(new_n746));
  XNOR2_X1  g321(.A(KEYINPUT95), .B(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT24), .ZN(new_n749));
  INV_X1    g324(.A(G34), .ZN(new_n750));
  AOI21_X1  g325(.A(G29), .B1(new_n749), .B2(new_n750), .ZN(new_n751));
  OAI21_X1  g326(.A(new_n751), .B1(new_n749), .B2(new_n750), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(G160), .B2(new_n721), .ZN(new_n753));
  OAI21_X1  g328(.A(new_n748), .B1(G2084), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(G27), .A2(G29), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n755), .B1(G164), .B2(G29), .ZN(new_n756));
  XOR2_X1   g331(.A(KEYINPUT99), .B(G2078), .Z(new_n757));
  XNOR2_X1  g332(.A(new_n756), .B(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n728), .A2(G20), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT100), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(KEYINPUT23), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G299), .B2(G16), .ZN(new_n762));
  INV_X1    g337(.A(G1956), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  NOR3_X1   g339(.A1(new_n754), .A2(new_n758), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n721), .A2(G33), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n487), .A2(G127), .ZN(new_n767));
  NAND2_X1  g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  AOI21_X1  g343(.A(new_n463), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n465), .A2(G103), .ZN(new_n770));
  OR2_X1    g345(.A1(new_n770), .A2(KEYINPUT25), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(KEYINPUT25), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g348(.A(new_n769), .B(new_n773), .C1(G139), .C2(new_n479), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n766), .B1(new_n774), .B2(new_n721), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(G2072), .ZN(new_n776));
  NOR2_X1   g351(.A1(G29), .A2(G32), .ZN(new_n777));
  NAND3_X1  g352(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT26), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(G105), .B2(new_n465), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n477), .A2(G129), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n479), .A2(G141), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(new_n783), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n777), .B1(new_n784), .B2(G29), .ZN(new_n785));
  XOR2_X1   g360(.A(KEYINPUT27), .B(G1996), .Z(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(new_n776), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n721), .A2(G35), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G162), .B2(new_n721), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n790), .B(KEYINPUT29), .ZN(new_n791));
  INV_X1    g366(.A(G2090), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n753), .A2(G2084), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n788), .A2(new_n793), .A3(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n555), .A2(new_n728), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(new_n728), .B2(G19), .ZN(new_n797));
  INV_X1    g372(.A(G1341), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n728), .A2(G4), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(new_n626), .B2(new_n728), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT93), .B(G1348), .ZN(new_n802));
  XOR2_X1   g377(.A(new_n802), .B(KEYINPUT94), .Z(new_n803));
  XNOR2_X1  g378(.A(new_n801), .B(new_n803), .ZN(new_n804));
  NOR3_X1   g379(.A1(new_n795), .A2(new_n799), .A3(new_n804), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n734), .A2(new_n735), .B1(new_n797), .B2(new_n798), .ZN(new_n806));
  NAND4_X1  g381(.A1(new_n737), .A2(new_n765), .A3(new_n805), .A4(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n479), .A2(KEYINPUT86), .A3(G131), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT86), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n487), .A2(new_n463), .ZN(new_n810));
  INV_X1    g385(.A(G131), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n477), .A2(G119), .ZN(new_n813));
  OR2_X1    g388(.A1(G95), .A2(G2105), .ZN(new_n814));
  OAI211_X1 g389(.A(new_n814), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n808), .A2(new_n812), .A3(new_n813), .A4(new_n815), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(KEYINPUT87), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G29), .ZN(new_n818));
  OAI21_X1  g393(.A(new_n818), .B1(G25), .B2(G29), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT88), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT35), .B(G1991), .ZN(new_n821));
  INV_X1    g396(.A(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n728), .A2(G24), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(new_n607), .B2(new_n728), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n825), .B(G1986), .Z(new_n826));
  AND2_X1   g401(.A1(new_n823), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(KEYINPUT92), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n728), .A2(G23), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n582), .A2(new_n586), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(new_n728), .ZN(new_n831));
  XNOR2_X1  g406(.A(KEYINPUT33), .B(G1976), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n832), .B(KEYINPUT90), .ZN(new_n833));
  OR2_X1    g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n833), .ZN(new_n835));
  XOR2_X1   g410(.A(KEYINPUT32), .B(G1981), .Z(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT89), .ZN(new_n837));
  AND2_X1   g412(.A1(new_n728), .A2(G6), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n838), .B1(G305), .B2(G16), .ZN(new_n839));
  OAI211_X1 g414(.A(new_n834), .B(new_n835), .C1(new_n837), .C2(new_n839), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n728), .A2(G22), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(G166), .B2(new_n728), .ZN(new_n842));
  INV_X1    g417(.A(G1971), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n842), .B(new_n843), .ZN(new_n844));
  INV_X1    g419(.A(new_n837), .ZN(new_n845));
  INV_X1    g420(.A(new_n839), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n844), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g422(.A(KEYINPUT91), .ZN(new_n848));
  OR3_X1    g423(.A1(new_n840), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  OAI21_X1  g424(.A(new_n848), .B1(new_n840), .B2(new_n847), .ZN(new_n850));
  AOI21_X1  g425(.A(KEYINPUT34), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n820), .A2(new_n822), .ZN(new_n853));
  NAND4_X1  g428(.A1(new_n827), .A2(new_n828), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n823), .A2(new_n853), .A3(new_n826), .ZN(new_n855));
  OAI21_X1  g430(.A(KEYINPUT92), .B1(new_n855), .B2(new_n851), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n849), .A2(KEYINPUT34), .A3(new_n850), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n859), .A2(KEYINPUT36), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT36), .ZN(new_n861));
  NAND3_X1  g436(.A1(new_n857), .A2(new_n861), .A3(new_n858), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n807), .B1(new_n860), .B2(new_n862), .ZN(G311));
  INV_X1    g438(.A(new_n807), .ZN(new_n864));
  INV_X1    g439(.A(new_n862), .ZN(new_n865));
  AOI21_X1  g440(.A(new_n861), .B1(new_n857), .B2(new_n858), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n864), .B1(new_n865), .B2(new_n866), .ZN(G150));
  INV_X1    g442(.A(KEYINPUT101), .ZN(new_n868));
  INV_X1    g443(.A(G67), .ZN(new_n869));
  NOR3_X1   g444(.A1(new_n518), .A2(new_n519), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(G80), .A2(G543), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  OAI21_X1  g447(.A(G651), .B1(new_n870), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G55), .ZN(new_n874));
  INV_X1    g449(.A(G93), .ZN(new_n875));
  OAI22_X1  g450(.A1(new_n505), .A2(new_n874), .B1(new_n875), .B2(new_n512), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n868), .B1(new_n873), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n547), .A2(G67), .A3(new_n548), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n500), .B1(new_n879), .B2(new_n871), .ZN(new_n880));
  NOR3_X1   g455(.A1(new_n880), .A2(KEYINPUT101), .A3(new_n876), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n878), .A2(new_n881), .ZN(new_n882));
  XOR2_X1   g457(.A(KEYINPUT103), .B(G860), .Z(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n884), .B(KEYINPUT37), .Z(new_n885));
  INV_X1    g460(.A(new_n554), .ZN(new_n886));
  INV_X1    g461(.A(new_n543), .ZN(new_n887));
  INV_X1    g462(.A(G56), .ZN(new_n888));
  NOR3_X1   g463(.A1(new_n518), .A2(new_n519), .A3(new_n888), .ZN(new_n889));
  INV_X1    g464(.A(new_n550), .ZN(new_n890));
  OAI21_X1  g465(.A(G651), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n891), .B2(KEYINPUT71), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n873), .A2(new_n868), .A3(new_n877), .ZN(new_n893));
  OAI21_X1  g468(.A(KEYINPUT101), .B1(new_n880), .B2(new_n876), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n886), .A2(new_n892), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n880), .A2(new_n876), .ZN(new_n896));
  NOR3_X1   g471(.A1(new_n553), .A2(new_n896), .A3(new_n554), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  NOR2_X1   g473(.A1(new_n618), .A2(new_n627), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT39), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n898), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n902));
  AND2_X1   g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OR2_X1    g478(.A1(new_n903), .A2(new_n883), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n901), .A2(new_n902), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n885), .B1(new_n904), .B2(new_n905), .ZN(G145));
  NAND2_X1  g481(.A1(new_n477), .A2(G130), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n479), .A2(G142), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n463), .A2(G118), .ZN(new_n909));
  OAI21_X1  g484(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n910));
  OAI211_X1 g485(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n774), .B(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n784), .A2(new_n743), .ZN(new_n914));
  INV_X1    g489(.A(new_n495), .ZN(new_n915));
  NAND2_X1  g490(.A1(new_n744), .A2(new_n783), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n914), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  INV_X1    g492(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(new_n915), .B1(new_n914), .B2(new_n916), .ZN(new_n919));
  NOR3_X1   g494(.A1(new_n918), .A2(new_n919), .A3(new_n635), .ZN(new_n920));
  INV_X1    g495(.A(new_n635), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n914), .A2(new_n916), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(new_n495), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n921), .B1(new_n923), .B2(new_n917), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n913), .B1(new_n920), .B2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n816), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n635), .B1(new_n918), .B2(new_n919), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n923), .A2(new_n921), .A3(new_n917), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n927), .A2(new_n912), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n925), .A2(new_n926), .A3(new_n929), .ZN(new_n930));
  AND2_X1   g505(.A1(new_n930), .A2(KEYINPUT104), .ZN(new_n931));
  INV_X1    g506(.A(new_n929), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n912), .B1(new_n927), .B2(new_n928), .ZN(new_n933));
  OAI21_X1  g508(.A(new_n816), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n931), .A2(new_n934), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n643), .B(new_n483), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(G160), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n935), .A2(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT105), .ZN(new_n940));
  INV_X1    g515(.A(G37), .ZN(new_n941));
  NAND4_X1  g516(.A1(new_n934), .A2(KEYINPUT104), .A3(new_n930), .A4(new_n937), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n939), .A2(new_n940), .A3(new_n941), .A4(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n937), .B1(new_n931), .B2(new_n934), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n942), .A2(new_n941), .ZN(new_n945));
  OAI21_X1  g520(.A(KEYINPUT105), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  XNOR2_X1  g522(.A(new_n947), .B(KEYINPUT40), .ZN(G395));
  XOR2_X1   g523(.A(new_n629), .B(KEYINPUT106), .Z(new_n949));
  XNOR2_X1  g524(.A(new_n949), .B(new_n898), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT41), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n626), .A2(G299), .ZN(new_n952));
  AND3_X1   g527(.A1(new_n574), .A2(new_n568), .A3(new_n569), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT107), .ZN(new_n954));
  NAND4_X1  g529(.A1(new_n618), .A2(new_n953), .A3(new_n954), .A4(new_n566), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  AND4_X1   g531(.A1(new_n566), .A2(new_n568), .A3(new_n569), .A4(new_n574), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n954), .B1(new_n957), .B2(new_n618), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n951), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(KEYINPUT107), .B1(new_n626), .B2(G299), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n960), .A2(KEYINPUT41), .A3(new_n952), .A4(new_n955), .ZN(new_n961));
  AND2_X1   g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n950), .A2(new_n962), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n960), .A2(new_n952), .A3(new_n955), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n950), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(KEYINPUT42), .ZN(new_n967));
  XNOR2_X1  g542(.A(new_n607), .B(G305), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n830), .B(G303), .ZN(new_n969));
  XNOR2_X1  g544(.A(new_n968), .B(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT42), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n963), .A2(new_n971), .A3(new_n965), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n967), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n970), .B1(new_n967), .B2(new_n972), .ZN(new_n974));
  OAI21_X1  g549(.A(G868), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n882), .A2(new_n619), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n975), .A2(new_n976), .ZN(G295));
  NAND2_X1  g552(.A1(new_n975), .A2(new_n976), .ZN(G331));
  OAI21_X1  g553(.A(KEYINPUT108), .B1(new_n521), .B2(new_n529), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n547), .A2(G63), .A3(G651), .A4(new_n548), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n537), .A2(G89), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT108), .ZN(new_n982));
  AND2_X1   g557(.A1(new_n527), .A2(new_n522), .ZN(new_n983));
  NAND4_X1  g558(.A1(new_n980), .A2(new_n981), .A3(new_n982), .A4(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n540), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n547), .A2(G64), .A3(new_n548), .ZN(new_n986));
  INV_X1    g561(.A(new_n535), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n500), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(new_n979), .B(new_n984), .C1(new_n985), .C2(new_n988), .ZN(new_n989));
  NAND4_X1  g564(.A1(new_n536), .A2(G168), .A3(new_n982), .A4(new_n540), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n895), .B2(new_n897), .ZN(new_n993));
  OAI22_X1  g568(.A1(new_n878), .A2(new_n881), .B1(new_n553), .B2(new_n554), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n873), .A2(new_n877), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n892), .A2(new_n886), .A3(new_n995), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n996), .A3(new_n991), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n993), .A2(new_n964), .A3(new_n997), .ZN(new_n998));
  INV_X1    g573(.A(new_n998), .ZN(new_n999));
  AND3_X1   g574(.A1(new_n994), .A2(new_n996), .A3(new_n991), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n991), .B1(new_n994), .B2(new_n996), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT109), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT109), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n993), .A2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n959), .A2(new_n961), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n999), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  AOI21_X1  g582(.A(G37), .B1(new_n1007), .B2(new_n970), .ZN(new_n1008));
  INV_X1    g583(.A(new_n970), .ZN(new_n1009));
  AOI21_X1  g584(.A(new_n962), .B1(new_n1002), .B2(new_n1004), .ZN(new_n1010));
  OAI21_X1  g585(.A(new_n1009), .B1(new_n1010), .B2(new_n999), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1008), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1012), .A2(KEYINPUT43), .ZN(new_n1013));
  OAI21_X1  g588(.A(new_n1006), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1002), .A2(new_n964), .A3(new_n1004), .ZN(new_n1015));
  OAI21_X1  g590(.A(new_n1014), .B1(new_n1015), .B2(KEYINPUT110), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT110), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1003), .B1(new_n993), .B2(new_n997), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1001), .A2(KEYINPUT109), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1018), .A2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1017), .B1(new_n1020), .B2(new_n964), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n1009), .B1(new_n1016), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n1008), .ZN(new_n1023));
  OAI21_X1  g598(.A(new_n1013), .B1(KEYINPUT43), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(KEYINPUT44), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1006), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1027));
  NAND3_X1  g602(.A1(new_n1027), .A2(new_n970), .A3(new_n998), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n941), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1020), .A2(new_n1017), .A3(new_n964), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1015), .A2(KEYINPUT110), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(new_n1031), .A3(new_n1014), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1009), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(KEYINPUT43), .ZN(new_n1034));
  OAI21_X1  g609(.A(KEYINPUT44), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n1011), .A2(new_n1034), .A3(new_n941), .A4(new_n1028), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(KEYINPUT111), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT111), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1008), .A2(new_n1038), .A3(new_n1034), .A4(new_n1011), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT112), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n1035), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(new_n1036), .B(new_n1038), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1025), .B1(new_n1023), .B2(KEYINPUT43), .ZN(new_n1044));
  AOI21_X1  g619(.A(KEYINPUT112), .B1(new_n1043), .B2(new_n1044), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1026), .B1(new_n1042), .B2(new_n1045), .ZN(G397));
  INV_X1    g621(.A(G1384), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n495), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT45), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1050));
  NAND4_X1  g625(.A1(new_n469), .A2(KEYINPUT113), .A3(G40), .A4(new_n473), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n464), .A2(new_n466), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT67), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1052), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g629(.A1(new_n464), .A2(KEYINPUT67), .A3(new_n466), .ZN(new_n1055));
  NAND4_X1  g630(.A1(new_n1054), .A2(new_n473), .A3(new_n1055), .A4(G40), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT113), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1050), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1059));
  XNOR2_X1  g634(.A(new_n743), .B(G2067), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1059), .B1(new_n783), .B2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(G1996), .ZN(new_n1062));
  AND2_X1   g637(.A1(new_n1059), .A2(new_n1062), .ZN(new_n1063));
  OR2_X1    g638(.A1(new_n1063), .A2(KEYINPUT115), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1059), .A2(KEYINPUT115), .A3(new_n1062), .ZN(new_n1065));
  AND3_X1   g640(.A1(new_n1064), .A2(KEYINPUT46), .A3(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(KEYINPUT46), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1061), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  OR2_X1    g643(.A1(new_n1068), .A2(KEYINPUT126), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(KEYINPUT126), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1069), .A2(KEYINPUT47), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(new_n784), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1074));
  OR2_X1    g649(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1074), .A2(KEYINPUT116), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n784), .A2(new_n1062), .ZN(new_n1077));
  AOI22_X1  g652(.A1(new_n1075), .A2(new_n1076), .B1(new_n1059), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n817), .A2(new_n822), .ZN(new_n1079));
  XNOR2_X1  g654(.A(new_n1079), .B(KEYINPUT125), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1073), .A2(new_n1078), .A3(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G2067), .B2(new_n743), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1082), .A2(new_n1059), .ZN(new_n1083));
  XNOR2_X1  g658(.A(new_n816), .B(new_n821), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1059), .A2(new_n1084), .ZN(new_n1085));
  NOR2_X1   g660(.A1(G290), .A2(G1986), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1086), .A2(new_n1059), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1087), .B(KEYINPUT48), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1073), .A2(new_n1078), .A3(new_n1085), .A4(new_n1088), .ZN(new_n1089));
  NAND3_X1  g664(.A1(new_n1071), .A2(new_n1083), .A3(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(KEYINPUT47), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT63), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n497), .A2(new_n1047), .A3(new_n498), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1094), .A2(KEYINPUT50), .ZN(new_n1095));
  AOI211_X1 g670(.A(KEYINPUT50), .B(G1384), .C1(new_n490), .C2(new_n494), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1096), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1095), .A2(new_n1097), .A3(new_n792), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1094), .A2(new_n1049), .ZN(new_n1100));
  AOI211_X1 g675(.A(new_n1049), .B(G1384), .C1(new_n490), .C2(new_n494), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1051), .B2(new_n1058), .ZN(new_n1102));
  AOI21_X1  g677(.A(G1971), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(KEYINPUT118), .B1(new_n1099), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n843), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT118), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1106), .A2(new_n1107), .A3(new_n1098), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1104), .A2(new_n1108), .A3(G8), .ZN(new_n1109));
  NAND2_X1  g684(.A1(G303), .A2(G8), .ZN(new_n1110));
  XNOR2_X1  g685(.A(new_n1110), .B(KEYINPUT55), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1109), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1051), .A2(new_n1058), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1048), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n830), .A2(G1976), .ZN(new_n1116));
  AND3_X1   g691(.A1(new_n1115), .A2(G8), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(G1976), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT52), .B1(G288), .B2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(G8), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1122), .A2(new_n1116), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1123), .A2(KEYINPUT52), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n598), .A2(new_n592), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(G1981), .ZN(new_n1126));
  INV_X1    g701(.A(G1981), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n594), .A2(new_n598), .A3(new_n1127), .A4(new_n599), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT49), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1126), .A2(KEYINPUT49), .A3(new_n1128), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1122), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  NAND3_X1  g708(.A1(new_n1120), .A2(new_n1124), .A3(new_n1133), .ZN(new_n1134));
  NAND4_X1  g709(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n1047), .A4(new_n498), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1113), .A2(new_n1135), .A3(new_n1050), .ZN(new_n1136));
  INV_X1    g711(.A(G1966), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(G2084), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1095), .A2(new_n1097), .A3(new_n1139), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1141), .A2(G8), .A3(G168), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g718(.A(new_n1093), .B1(new_n1112), .B2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT50), .ZN(new_n1145));
  NAND4_X1  g720(.A1(new_n497), .A2(new_n1145), .A3(new_n1047), .A4(new_n498), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1048), .A2(KEYINPUT50), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1113), .A2(new_n1146), .A3(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1148), .A2(G2090), .ZN(new_n1149));
  OAI21_X1  g724(.A(G8), .B1(new_n1149), .B2(new_n1103), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1150), .A2(new_n1111), .ZN(new_n1151));
  AOI211_X1 g726(.A(new_n1121), .B(G286), .C1(new_n1138), .C2(new_n1140), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1151), .A2(new_n1093), .A3(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(new_n1111), .ZN(new_n1154));
  NAND4_X1  g729(.A1(new_n1104), .A2(new_n1108), .A3(G8), .A4(new_n1154), .ZN(new_n1155));
  AOI21_X1  g730(.A(new_n1134), .B1(new_n1153), .B2(new_n1155), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G288), .A2(G1976), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1133), .A2(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1158), .A2(new_n1128), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT120), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(KEYINPUT120), .B1(new_n1158), .B2(new_n1128), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1122), .B(KEYINPUT119), .ZN(new_n1163));
  NOR3_X1   g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NOR3_X1   g739(.A1(new_n1144), .A2(new_n1156), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT121), .ZN(new_n1166));
  OR2_X1    g741(.A1(new_n1166), .A2(KEYINPUT57), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1166), .A2(KEYINPUT57), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n957), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g744(.A1(G299), .A2(new_n1166), .A3(KEYINPUT57), .ZN(new_n1170));
  NAND2_X1  g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n1148), .A2(new_n763), .ZN(new_n1173));
  XNOR2_X1  g748(.A(KEYINPUT56), .B(G2072), .ZN(new_n1174));
  NAND3_X1  g749(.A1(new_n1100), .A2(new_n1102), .A3(new_n1174), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1172), .B1(new_n1173), .B2(new_n1175), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1095), .A2(new_n1097), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1177), .A2(new_n802), .ZN(new_n1178));
  INV_X1    g753(.A(G2067), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1113), .A2(new_n1179), .A3(new_n1114), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n618), .B1(new_n1178), .B2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1173), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1176), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(KEYINPUT61), .ZN(new_n1184));
  AND3_X1   g759(.A1(new_n1173), .A2(new_n1172), .A3(new_n1175), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1184), .B1(new_n1185), .B2(new_n1176), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1173), .A2(new_n1175), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1187), .A2(new_n1171), .ZN(new_n1188));
  NAND3_X1  g763(.A1(new_n1188), .A2(KEYINPUT61), .A3(new_n1182), .ZN(new_n1189));
  NOR2_X1   g764(.A1(new_n1105), .A2(G1996), .ZN(new_n1190));
  XNOR2_X1  g765(.A(KEYINPUT58), .B(G1341), .ZN(new_n1191));
  AOI21_X1  g766(.A(new_n1191), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1192));
  OAI21_X1  g767(.A(new_n555), .B1(new_n1190), .B2(new_n1192), .ZN(new_n1193));
  INV_X1    g768(.A(KEYINPUT59), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(new_n1194), .ZN(new_n1195));
  OAI211_X1 g770(.A(KEYINPUT59), .B(new_n555), .C1(new_n1190), .C2(new_n1192), .ZN(new_n1196));
  NAND4_X1  g771(.A1(new_n1186), .A2(new_n1189), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  NAND2_X1  g772(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1198));
  INV_X1    g773(.A(KEYINPUT60), .ZN(new_n1199));
  OAI21_X1  g774(.A(new_n626), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g775(.A1(new_n1178), .A2(KEYINPUT60), .A3(new_n618), .A4(new_n1180), .ZN(new_n1201));
  AOI22_X1  g776(.A1(new_n1200), .A2(new_n1201), .B1(new_n1199), .B2(new_n1198), .ZN(new_n1202));
  OAI21_X1  g777(.A(new_n1183), .B1(new_n1197), .B2(new_n1202), .ZN(new_n1203));
  INV_X1    g778(.A(G2078), .ZN(new_n1204));
  NAND3_X1  g779(.A1(new_n1100), .A2(new_n1102), .A3(new_n1204), .ZN(new_n1205));
  INV_X1    g780(.A(KEYINPUT53), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g782(.A1(new_n1177), .A2(new_n735), .ZN(new_n1208));
  AOI211_X1 g783(.A(new_n1206), .B(G2078), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1209));
  NAND3_X1  g784(.A1(new_n1209), .A2(new_n1113), .A3(new_n1135), .ZN(new_n1210));
  NAND3_X1  g785(.A1(new_n1207), .A2(new_n1208), .A3(new_n1210), .ZN(new_n1211));
  XNOR2_X1  g786(.A(G301), .B(KEYINPUT54), .ZN(new_n1212));
  AOI22_X1  g787(.A1(new_n1205), .A2(new_n1206), .B1(new_n1177), .B2(new_n735), .ZN(new_n1213));
  INV_X1    g788(.A(new_n472), .ZN(new_n1214));
  AOI21_X1  g789(.A(new_n463), .B1(new_n1214), .B2(KEYINPUT123), .ZN(new_n1215));
  OAI21_X1  g790(.A(new_n1215), .B1(KEYINPUT123), .B2(new_n1214), .ZN(new_n1216));
  NAND3_X1  g791(.A1(new_n1216), .A2(new_n469), .A3(G40), .ZN(new_n1217));
  NOR2_X1   g792(.A1(new_n1217), .A2(new_n1101), .ZN(new_n1218));
  AOI21_X1  g793(.A(new_n1212), .B1(new_n1209), .B2(new_n1218), .ZN(new_n1219));
  AOI22_X1  g794(.A1(new_n1211), .A2(new_n1212), .B1(new_n1213), .B2(new_n1219), .ZN(new_n1220));
  INV_X1    g795(.A(KEYINPUT52), .ZN(new_n1221));
  OAI21_X1  g796(.A(new_n1133), .B1(new_n1117), .B2(new_n1221), .ZN(new_n1222));
  AND3_X1   g797(.A1(new_n1119), .A2(new_n1122), .A3(new_n1116), .ZN(new_n1223));
  NOR2_X1   g798(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  NAND4_X1  g799(.A1(new_n1220), .A2(new_n1155), .A3(new_n1224), .A4(new_n1151), .ZN(new_n1225));
  NAND2_X1  g800(.A1(new_n1141), .A2(G8), .ZN(new_n1226));
  NOR2_X1   g801(.A1(G168), .A2(new_n1121), .ZN(new_n1227));
  INV_X1    g802(.A(new_n1227), .ZN(new_n1228));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n1229));
  OAI21_X1  g804(.A(KEYINPUT51), .B1(new_n1227), .B2(new_n1229), .ZN(new_n1230));
  NAND3_X1  g805(.A1(new_n1226), .A2(new_n1228), .A3(new_n1230), .ZN(new_n1231));
  INV_X1    g806(.A(new_n1230), .ZN(new_n1232));
  OAI211_X1 g807(.A(G8), .B(new_n1232), .C1(new_n1141), .C2(G286), .ZN(new_n1233));
  AOI22_X1  g808(.A1(new_n1231), .A2(new_n1233), .B1(new_n1227), .B2(new_n1141), .ZN(new_n1234));
  NOR2_X1   g809(.A1(new_n1225), .A2(new_n1234), .ZN(new_n1235));
  NAND2_X1  g810(.A1(new_n1203), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n1237));
  AND3_X1   g812(.A1(new_n1165), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  AOI21_X1  g813(.A(new_n1237), .B1(new_n1165), .B2(new_n1236), .ZN(new_n1239));
  AOI21_X1  g814(.A(G301), .B1(new_n1213), .B2(new_n1210), .ZN(new_n1240));
  NAND4_X1  g815(.A1(new_n1155), .A2(new_n1224), .A3(new_n1151), .A4(new_n1240), .ZN(new_n1241));
  OR2_X1    g816(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1242));
  NAND2_X1  g817(.A1(new_n1234), .A2(KEYINPUT62), .ZN(new_n1243));
  AOI21_X1  g818(.A(new_n1241), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1244));
  NOR3_X1   g819(.A1(new_n1238), .A2(new_n1239), .A3(new_n1244), .ZN(new_n1245));
  AND2_X1   g820(.A1(G290), .A2(G1986), .ZN(new_n1246));
  OR3_X1    g821(.A1(new_n1246), .A2(new_n1086), .A3(KEYINPUT114), .ZN(new_n1247));
  NAND3_X1  g822(.A1(G290), .A2(KEYINPUT114), .A3(G1986), .ZN(new_n1248));
  NAND3_X1  g823(.A1(new_n1247), .A2(new_n1059), .A3(new_n1248), .ZN(new_n1249));
  NAND4_X1  g824(.A1(new_n1073), .A2(new_n1078), .A3(new_n1085), .A4(new_n1249), .ZN(new_n1250));
  XNOR2_X1  g825(.A(new_n1250), .B(KEYINPUT117), .ZN(new_n1251));
  OAI21_X1  g826(.A(new_n1092), .B1(new_n1245), .B2(new_n1251), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g827(.A(G319), .ZN(new_n1254));
  NOR2_X1   g828(.A1(G227), .A2(new_n1254), .ZN(new_n1255));
  NAND3_X1  g829(.A1(new_n671), .A2(new_n717), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g830(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1257));
  INV_X1    g831(.A(KEYINPUT127), .ZN(new_n1258));
  NAND4_X1  g832(.A1(new_n671), .A2(new_n717), .A3(new_n1258), .A4(new_n1255), .ZN(new_n1259));
  NAND4_X1  g833(.A1(new_n1257), .A2(new_n947), .A3(new_n1024), .A4(new_n1259), .ZN(G225));
  INV_X1    g834(.A(G225), .ZN(G308));
endmodule


