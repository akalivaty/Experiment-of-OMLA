//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 1 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:01 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1240, new_n1241, new_n1242,
    new_n1243, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1287,
    new_n1288, new_n1289, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  NAND2_X1  g0008(.A1(G1), .A2(G20), .ZN(new_n209));
  XNOR2_X1  g0009(.A(KEYINPUT65), .B(G244), .ZN(new_n210));
  AND2_X1   g0010(.A1(new_n210), .A2(G77), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G58), .A2(G232), .B1(G87), .B2(G250), .ZN(new_n212));
  AOI22_X1  g0012(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n213));
  AOI22_X1  g0013(.A1(G97), .A2(G257), .B1(G116), .B2(G270), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G107), .A2(G264), .ZN(new_n215));
  NAND4_X1  g0015(.A1(new_n212), .A2(new_n213), .A3(new_n214), .A4(new_n215), .ZN(new_n216));
  OAI21_X1  g0016(.A(new_n209), .B1(new_n211), .B2(new_n216), .ZN(new_n217));
  OR2_X1    g0017(.A1(new_n217), .A2(KEYINPUT1), .ZN(new_n218));
  XOR2_X1   g0018(.A(new_n218), .B(KEYINPUT66), .Z(new_n219));
  NOR2_X1   g0019(.A1(new_n209), .A2(G13), .ZN(new_n220));
  INV_X1    g0020(.A(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(G250), .B1(G257), .B2(G264), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(G20), .ZN(new_n225));
  NOR2_X1   g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  INV_X1    g0026(.A(new_n226), .ZN(new_n227));
  INV_X1    g0027(.A(new_n201), .ZN(new_n228));
  NAND2_X1  g0028(.A1(new_n228), .A2(G50), .ZN(new_n229));
  OAI22_X1  g0029(.A1(new_n223), .A2(KEYINPUT0), .B1(new_n227), .B2(new_n229), .ZN(new_n230));
  AOI21_X1  g0030(.A(new_n230), .B1(KEYINPUT0), .B2(new_n223), .ZN(new_n231));
  XOR2_X1   g0031(.A(new_n231), .B(KEYINPUT64), .Z(new_n232));
  AOI211_X1 g0032(.A(new_n219), .B(new_n232), .C1(KEYINPUT1), .C2(new_n217), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT2), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(G226), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G250), .B(G257), .Z(new_n239));
  XNOR2_X1  g0039(.A(G264), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XOR2_X1   g0045(.A(G87), .B(G97), .Z(new_n246));
  XNOR2_X1  g0046(.A(G107), .B(G116), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n245), .B(new_n248), .ZN(G351));
  NOR2_X1   g0049(.A1(G20), .A2(G33), .ZN(new_n250));
  AOI22_X1  g0050(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(KEYINPUT8), .B(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n225), .A2(G33), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n251), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g0054(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n224), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G1), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n258), .A2(G13), .A3(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n260), .A2(new_n256), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n202), .B1(new_n258), .B2(G20), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n261), .A2(new_n262), .B1(new_n202), .B2(new_n260), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n257), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g0064(.A(KEYINPUT3), .B(G33), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(G223), .A3(G1698), .ZN(new_n266));
  INV_X1    g0066(.A(G77), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n265), .A2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G222), .ZN(new_n270));
  OAI221_X1 g0070(.A(new_n266), .B1(new_n267), .B2(new_n265), .C1(new_n269), .C2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n258), .B1(G41), .B2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  NOR2_X1   g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(new_n274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n272), .A2(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n276), .B1(new_n278), .B2(G226), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G179), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G169), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n283), .B1(new_n273), .B2(new_n279), .ZN(new_n284));
  OAI21_X1  g0084(.A(new_n264), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  XOR2_X1   g0085(.A(new_n285), .B(KEYINPUT67), .Z(new_n286));
  XNOR2_X1  g0086(.A(new_n264), .B(KEYINPUT9), .ZN(new_n287));
  XNOR2_X1  g0087(.A(KEYINPUT70), .B(G200), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n280), .A2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G190), .ZN(new_n291));
  OAI211_X1 g0091(.A(new_n287), .B(new_n290), .C1(new_n291), .C2(new_n280), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT10), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n265), .A2(G238), .A3(G1698), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n294), .B1(new_n206), .B2(new_n265), .C1(new_n269), .C2(new_n237), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n272), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n276), .B1(new_n278), .B2(new_n210), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n298), .A2(G190), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n299), .B1(new_n298), .B2(new_n288), .ZN(new_n300));
  INV_X1    g0100(.A(new_n252), .ZN(new_n301));
  AOI22_X1  g0101(.A1(new_n301), .A2(new_n250), .B1(G20), .B2(G77), .ZN(new_n302));
  XNOR2_X1  g0102(.A(KEYINPUT15), .B(G87), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n303), .B(KEYINPUT68), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n302), .B1(new_n304), .B2(new_n253), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n305), .A2(new_n256), .B1(new_n267), .B2(new_n260), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n258), .A2(G20), .ZN(new_n307));
  NAND3_X1  g0107(.A1(new_n261), .A2(G77), .A3(new_n307), .ZN(new_n308));
  XNOR2_X1  g0108(.A(new_n308), .B(KEYINPUT69), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n300), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n298), .A2(G169), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n312), .B1(new_n281), .B2(new_n298), .ZN(new_n313));
  AND2_X1   g0113(.A1(new_n313), .A2(new_n310), .ZN(new_n314));
  NOR2_X1   g0114(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n265), .A2(G232), .A3(G1698), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  INV_X1    g0117(.A(G226), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(new_n269), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n272), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n276), .B1(new_n278), .B2(G238), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(KEYINPUT13), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT13), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(new_n324), .A3(new_n321), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G190), .B2(new_n326), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n261), .A2(G68), .A3(new_n307), .ZN(new_n330));
  INV_X1    g0130(.A(G13), .ZN(new_n331));
  NOR2_X1   g0131(.A1(new_n331), .A2(G1), .ZN(new_n332));
  INV_X1    g0132(.A(G68), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(G20), .A3(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(KEYINPUT71), .A3(KEYINPUT12), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(KEYINPUT12), .B2(new_n334), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT71), .B1(new_n334), .B2(KEYINPUT12), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n330), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT72), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n250), .ZN(new_n341));
  OAI22_X1  g0141(.A1(new_n341), .A2(new_n202), .B1(new_n225), .B2(G68), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n253), .A2(new_n267), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n256), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  XNOR2_X1  g0144(.A(new_n344), .B(KEYINPUT11), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n329), .A2(new_n347), .ZN(new_n348));
  AND4_X1   g0148(.A1(new_n286), .A2(new_n293), .A3(new_n315), .A4(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n252), .B1(new_n258), .B2(G20), .ZN(new_n350));
  AOI22_X1  g0150(.A1(new_n350), .A2(new_n261), .B1(new_n260), .B2(new_n252), .ZN(new_n351));
  INV_X1    g0151(.A(G33), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(KEYINPUT3), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT3), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(G33), .ZN(new_n355));
  NAND4_X1  g0155(.A1(new_n353), .A2(new_n355), .A3(G223), .A4(new_n268), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n353), .A2(new_n355), .A3(G226), .A4(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n359), .A2(new_n272), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n276), .B1(new_n278), .B2(G232), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n360), .A2(new_n361), .A3(new_n291), .ZN(new_n362));
  INV_X1    g0162(.A(G41), .ZN(new_n363));
  OAI211_X1 g0163(.A(G1), .B(G13), .C1(new_n352), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n364), .A2(G232), .A3(new_n274), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n365), .B1(new_n275), .B2(new_n274), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n366), .B1(new_n272), .B2(new_n359), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n362), .B1(new_n367), .B2(G200), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT74), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n369), .B1(new_n352), .B2(KEYINPUT3), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT73), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n354), .B2(G33), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n354), .A2(KEYINPUT74), .A3(G33), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n352), .A2(KEYINPUT73), .A3(KEYINPUT3), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n370), .A2(new_n372), .A3(new_n373), .A4(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT7), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n376), .A2(G20), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n265), .B2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G68), .ZN(new_n381));
  INV_X1    g0181(.A(G58), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n382), .A2(new_n333), .ZN(new_n383));
  OAI21_X1  g0183(.A(G20), .B1(new_n383), .B2(new_n201), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n250), .A2(G159), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n386), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT16), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n353), .A2(new_n355), .ZN(new_n389));
  AOI21_X1  g0189(.A(KEYINPUT7), .B1(new_n389), .B2(new_n225), .ZN(new_n390));
  AOI211_X1 g0190(.A(new_n376), .B(G20), .C1(new_n353), .C2(new_n355), .ZN(new_n391));
  OAI21_X1  g0191(.A(G68), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n392), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(new_n256), .ZN(new_n394));
  OAI211_X1 g0194(.A(new_n351), .B(new_n368), .C1(new_n388), .C2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(KEYINPUT17), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(KEYINPUT75), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT75), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n395), .A2(new_n399), .A3(KEYINPUT17), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n396), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n351), .B1(new_n388), .B2(new_n394), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n367), .A2(new_n281), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n360), .A2(new_n361), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(new_n283), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  INV_X1    g0206(.A(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n402), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n351), .ZN(new_n410));
  INV_X1    g0210(.A(new_n256), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n389), .A2(KEYINPUT7), .A3(new_n225), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n379), .A2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n386), .B1(new_n413), .B2(G68), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n414), .B2(KEYINPUT16), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT16), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n333), .B1(new_n378), .B2(new_n379), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n416), .B1(new_n417), .B2(new_n386), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n410), .B1(new_n415), .B2(new_n418), .ZN(new_n419));
  OAI21_X1  g0219(.A(KEYINPUT18), .B1(new_n419), .B2(new_n406), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n409), .A2(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n401), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n283), .B1(new_n323), .B2(new_n325), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT14), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI22_X1  g0226(.A1(new_n423), .A2(new_n424), .B1(new_n326), .B2(new_n281), .ZN(new_n427));
  OAI21_X1  g0227(.A(new_n346), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  AND3_X1   g0228(.A1(new_n349), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT4), .ZN(new_n430));
  AOI21_X1  g0230(.A(G1698), .B1(new_n430), .B2(KEYINPUT80), .ZN(new_n431));
  NAND4_X1  g0231(.A1(new_n431), .A2(G244), .A3(new_n353), .A4(new_n355), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n430), .A2(KEYINPUT80), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n265), .A2(G244), .A3(new_n431), .A4(new_n433), .ZN(new_n436));
  NAND2_X1  g0236(.A1(G33), .A2(G283), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n265), .A2(G250), .A3(G1698), .ZN(new_n438));
  NAND4_X1  g0238(.A1(new_n435), .A2(new_n436), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(new_n272), .ZN(new_n440));
  OR2_X1    g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  NAND2_X1  g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n258), .A2(G45), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n446), .A2(G257), .A3(new_n364), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n444), .B1(new_n441), .B2(new_n442), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(G274), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n440), .A2(new_n291), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n439), .B2(new_n272), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n452), .B1(G200), .B2(new_n453), .ZN(new_n454));
  AOI21_X1  g0254(.A(new_n206), .B1(new_n378), .B2(new_n379), .ZN(new_n455));
  NAND2_X1  g0255(.A1(G97), .A2(G107), .ZN(new_n456));
  INV_X1    g0256(.A(new_n456), .ZN(new_n457));
  NOR2_X1   g0257(.A1(G97), .A2(G107), .ZN(new_n458));
  OAI21_X1  g0258(.A(KEYINPUT77), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT77), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n207), .A2(new_n460), .A3(new_n456), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT6), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n459), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  AND2_X1   g0263(.A1(KEYINPUT76), .A2(G97), .ZN(new_n464));
  NOR2_X1   g0264(.A1(KEYINPUT76), .A2(G97), .ZN(new_n465));
  OAI211_X1 g0265(.A(KEYINPUT6), .B(new_n206), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  AOI21_X1  g0266(.A(new_n225), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n341), .A2(new_n267), .ZN(new_n468));
  NOR3_X1   g0268(.A1(new_n455), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  OAI21_X1  g0269(.A(KEYINPUT78), .B1(new_n469), .B2(new_n411), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT78), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n390), .B1(new_n375), .B2(new_n377), .ZN(new_n472));
  OAI22_X1  g0272(.A1(new_n472), .A2(new_n206), .B1(new_n267), .B2(new_n341), .ZN(new_n473));
  OAI211_X1 g0273(.A(new_n471), .B(new_n256), .C1(new_n473), .C2(new_n467), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n260), .A2(new_n205), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n258), .A2(G33), .ZN(new_n476));
  NAND4_X1  g0276(.A1(new_n259), .A2(new_n476), .A3(new_n224), .A4(new_n255), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n475), .B1(new_n477), .B2(new_n205), .ZN(new_n478));
  XNOR2_X1  g0278(.A(new_n478), .B(KEYINPUT79), .ZN(new_n479));
  INV_X1    g0279(.A(new_n479), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n454), .A2(new_n470), .A3(new_n474), .A4(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(KEYINPUT81), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n455), .A2(new_n468), .ZN(new_n483));
  INV_X1    g0283(.A(new_n467), .ZN(new_n484));
  AOI21_X1  g0284(.A(new_n411), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n479), .B1(new_n485), .B2(new_n471), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  NAND4_X1  g0287(.A1(new_n486), .A2(new_n487), .A3(new_n470), .A4(new_n454), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n470), .A2(new_n474), .A3(new_n480), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n453), .A2(G169), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n440), .A2(new_n451), .ZN(new_n491));
  OAI21_X1  g0291(.A(KEYINPUT82), .B1(new_n491), .B2(G179), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n453), .A2(new_n493), .A3(new_n281), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  AOI22_X1  g0295(.A1(new_n482), .A2(new_n488), .B1(new_n489), .B2(new_n495), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n353), .A2(new_n355), .A3(G250), .A4(new_n268), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n353), .A2(new_n355), .A3(G257), .A4(G1698), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G294), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n497), .A2(new_n498), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(new_n272), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n446), .A2(G264), .A3(new_n364), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(new_n449), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(new_n327), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n448), .A2(new_n272), .ZN(new_n505));
  AOI22_X1  g0305(.A1(new_n272), .A2(new_n500), .B1(new_n505), .B2(G264), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n506), .A2(new_n291), .A3(new_n449), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n504), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n332), .A2(G20), .A3(new_n206), .ZN(new_n509));
  XNOR2_X1  g0309(.A(new_n509), .B(KEYINPUT25), .ZN(new_n510));
  INV_X1    g0310(.A(new_n477), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n510), .B1(new_n511), .B2(G107), .ZN(new_n512));
  NAND4_X1  g0312(.A1(new_n353), .A2(new_n355), .A3(new_n225), .A4(G87), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT85), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT85), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n265), .A2(new_n515), .A3(new_n225), .A4(G87), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT22), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n514), .A2(new_n516), .A3(KEYINPUT22), .ZN(new_n520));
  OAI21_X1  g0320(.A(KEYINPUT86), .B1(new_n225), .B2(G107), .ZN(new_n521));
  INV_X1    g0321(.A(KEYINPUT23), .ZN(new_n522));
  OR2_X1    g0322(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n522), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n225), .A2(G33), .A3(G116), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n519), .A2(KEYINPUT24), .A3(new_n520), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n256), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n526), .B1(new_n517), .B2(new_n518), .ZN(new_n530));
  AOI21_X1  g0330(.A(KEYINPUT24), .B1(new_n530), .B2(new_n520), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n508), .B(new_n512), .C1(new_n529), .C2(new_n531), .ZN(new_n532));
  INV_X1    g0332(.A(new_n465), .ZN(new_n533));
  INV_X1    g0333(.A(G87), .ZN(new_n534));
  NAND2_X1  g0334(.A1(KEYINPUT76), .A2(G97), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n533), .A2(new_n534), .A3(new_n206), .A4(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT19), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n537), .B1(new_n317), .B2(new_n225), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n464), .A2(new_n465), .ZN(new_n540));
  OAI21_X1  g0340(.A(new_n537), .B1(new_n540), .B2(new_n253), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n265), .A2(new_n225), .A3(G68), .ZN(new_n542));
  NAND3_X1  g0342(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n543), .A2(new_n256), .B1(new_n304), .B2(new_n260), .ZN(new_n544));
  OAI21_X1  g0344(.A(new_n544), .B1(new_n304), .B2(new_n477), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n444), .A2(G250), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n546), .B1(new_n275), .B2(new_n444), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n364), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n353), .A2(new_n355), .A3(G244), .A4(G1698), .ZN(new_n549));
  NAND4_X1  g0349(.A1(new_n353), .A2(new_n355), .A3(G238), .A4(new_n268), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n549), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT83), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n549), .A2(new_n550), .A3(KEYINPUT83), .A4(new_n551), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n272), .ZN(new_n557));
  OAI211_X1 g0357(.A(new_n281), .B(new_n548), .C1(new_n555), .C2(new_n557), .ZN(new_n558));
  AND2_X1   g0358(.A1(new_n556), .A2(new_n272), .ZN(new_n559));
  AOI22_X1  g0359(.A1(new_n559), .A2(new_n554), .B1(new_n364), .B2(new_n547), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n545), .B(new_n558), .C1(G169), .C2(new_n560), .ZN(new_n561));
  OR3_X1    g0361(.A1(new_n477), .A2(KEYINPUT84), .A3(new_n534), .ZN(new_n562));
  OAI21_X1  g0362(.A(KEYINPUT84), .B1(new_n477), .B2(new_n534), .ZN(new_n563));
  AND2_X1   g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n544), .A2(new_n564), .ZN(new_n565));
  OAI21_X1  g0365(.A(new_n548), .B1(new_n555), .B2(new_n557), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(new_n289), .ZN(new_n567));
  OAI211_X1 g0367(.A(G190), .B(new_n548), .C1(new_n555), .C2(new_n557), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n565), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n532), .A2(new_n561), .A3(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n352), .B1(new_n464), .B2(new_n465), .ZN(new_n571));
  AOI21_X1  g0371(.A(G20), .B1(new_n571), .B2(new_n437), .ZN(new_n572));
  INV_X1    g0372(.A(G116), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n225), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n256), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(KEYINPUT20), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(KEYINPUT20), .B(new_n256), .C1(new_n572), .C2(new_n574), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n477), .A2(G116), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n259), .A2(new_n573), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g0383(.A1(new_n505), .A2(G270), .B1(G274), .B2(new_n448), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n353), .A2(new_n355), .A3(G264), .A4(G1698), .ZN(new_n585));
  NAND4_X1  g0385(.A1(new_n353), .A2(new_n355), .A3(G257), .A4(new_n268), .ZN(new_n586));
  INV_X1    g0386(.A(G303), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n585), .B(new_n586), .C1(new_n587), .C2(new_n265), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(new_n272), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n584), .A2(G179), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  AOI211_X1 g0391(.A(new_n591), .B(new_n283), .C1(new_n584), .C2(new_n589), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n583), .B1(new_n590), .B2(new_n592), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n577), .A2(new_n578), .B1(new_n581), .B2(new_n580), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n584), .A2(new_n589), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G169), .ZN(new_n596));
  OAI21_X1  g0396(.A(new_n591), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(G200), .B1(new_n584), .B2(new_n589), .ZN(new_n598));
  AND3_X1   g0398(.A1(new_n584), .A2(new_n291), .A3(new_n589), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n594), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n593), .A2(new_n597), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n519), .A2(new_n520), .A3(new_n527), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND3_X1  g0404(.A1(new_n604), .A2(new_n256), .A3(new_n528), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n506), .A2(G179), .A3(new_n449), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n503), .A2(G169), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n605), .A2(new_n512), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n570), .A2(new_n601), .A3(new_n608), .ZN(new_n609));
  AND3_X1   g0409(.A1(new_n429), .A2(new_n496), .A3(new_n609), .ZN(G372));
  INV_X1    g0410(.A(new_n286), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n421), .B(KEYINPUT90), .ZN(new_n612));
  INV_X1    g0412(.A(new_n428), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n613), .B1(new_n314), .B2(new_n348), .ZN(new_n614));
  OAI21_X1  g0414(.A(new_n612), .B1(new_n614), .B2(new_n401), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n611), .B1(new_n615), .B2(new_n293), .ZN(new_n616));
  INV_X1    g0416(.A(new_n429), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT88), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n565), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n544), .A2(new_n563), .A3(new_n562), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT88), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n566), .A2(KEYINPUT87), .A3(new_n289), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT87), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n567), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n622), .A2(new_n568), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  AND3_X1   g0426(.A1(new_n626), .A2(new_n532), .A3(new_n561), .ZN(new_n627));
  INV_X1    g0427(.A(new_n608), .ZN(new_n628));
  AND2_X1   g0428(.A1(new_n593), .A2(new_n597), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n627), .A2(new_n496), .A3(new_n630), .ZN(new_n631));
  AND2_X1   g0431(.A1(new_n495), .A2(new_n489), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT26), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n632), .A2(new_n626), .A3(new_n633), .A4(new_n561), .ZN(new_n634));
  INV_X1    g0434(.A(new_n561), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n495), .A2(new_n489), .A3(new_n561), .A4(new_n569), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n636), .B2(KEYINPUT26), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT89), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n634), .B2(new_n637), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n631), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n616), .B1(new_n617), .B2(new_n642), .ZN(G369));
  INV_X1    g0443(.A(new_n332), .ZN(new_n644));
  OR3_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .A3(G20), .ZN(new_n645));
  OAI21_X1  g0445(.A(KEYINPUT27), .B1(new_n644), .B2(G20), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(G343), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NOR2_X1   g0450(.A1(new_n594), .A2(new_n650), .ZN(new_n651));
  MUX2_X1   g0451(.A(new_n601), .B(new_n629), .S(new_n651), .Z(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT91), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n653), .A2(G330), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n605), .A2(new_n512), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n649), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n608), .B1(new_n657), .B2(new_n532), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n608), .A2(new_n650), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n655), .A2(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n629), .A2(new_n649), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT92), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n659), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n662), .A2(new_n667), .ZN(G399));
  NOR2_X1   g0468(.A1(new_n221), .A2(G41), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n670), .A2(G1), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n536), .A2(G116), .ZN(new_n672));
  OAI22_X1  g0472(.A1(new_n671), .A2(new_n672), .B1(new_n229), .B2(new_n670), .ZN(new_n673));
  XNOR2_X1  g0473(.A(new_n673), .B(KEYINPUT28), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT29), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n642), .B2(new_n649), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n626), .A2(new_n561), .ZN(new_n677));
  INV_X1    g0477(.A(new_n632), .ZN(new_n678));
  OAI21_X1  g0478(.A(KEYINPUT26), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  OAI211_X1 g0479(.A(new_n679), .B(new_n561), .C1(KEYINPUT26), .C2(new_n636), .ZN(new_n680));
  INV_X1    g0480(.A(new_n631), .ZN(new_n681));
  OAI211_X1 g0481(.A(KEYINPUT29), .B(new_n650), .C1(new_n680), .C2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n676), .A2(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n496), .A2(new_n609), .A3(new_n650), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT95), .ZN(new_n685));
  AOI21_X1  g0485(.A(G179), .B1(new_n584), .B2(new_n589), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n491), .A2(new_n566), .A3(new_n686), .A4(new_n503), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n560), .A2(new_n590), .A3(new_n453), .A4(new_n506), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT30), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n687), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n440), .A2(new_n451), .A3(new_n506), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n584), .A2(G179), .A3(new_n589), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(KEYINPUT30), .B1(new_n693), .B2(new_n560), .ZN(new_n694));
  OAI211_X1 g0494(.A(KEYINPUT31), .B(new_n649), .C1(new_n690), .C2(new_n694), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT93), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT94), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n690), .B2(new_n694), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n693), .A2(KEYINPUT30), .A3(new_n560), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n688), .A2(new_n689), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n699), .A2(new_n700), .A3(KEYINPUT94), .A4(new_n687), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(new_n649), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT31), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT95), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n496), .A2(new_n609), .A3(new_n706), .A4(new_n650), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n685), .A2(new_n696), .A3(new_n705), .A4(new_n707), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(G330), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  OR3_X1    g0510(.A1(new_n683), .A2(KEYINPUT96), .A3(new_n710), .ZN(new_n711));
  OAI21_X1  g0511(.A(KEYINPUT96), .B1(new_n683), .B2(new_n710), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n674), .B1(new_n713), .B2(G1), .ZN(G364));
  NOR2_X1   g0514(.A1(G13), .A2(G33), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(G20), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n652), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n331), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n671), .B1(G45), .B2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  XOR2_X1   g0521(.A(G355), .B(KEYINPUT97), .Z(new_n722));
  NOR2_X1   g0522(.A1(new_n221), .A2(new_n389), .ZN(new_n723));
  AOI22_X1  g0523(.A1(new_n722), .A2(new_n723), .B1(new_n573), .B2(new_n221), .ZN(new_n724));
  AOI21_X1  g0524(.A(G45), .B1(new_n228), .B2(G50), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n725), .B1(new_n245), .B2(G45), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n221), .A2(new_n265), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n724), .B1(new_n726), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n224), .B1(G20), .B2(new_n283), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n717), .A2(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n721), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(G20), .A2(G179), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT98), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n291), .A2(G200), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(G322), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g0538(.A1(G179), .A2(G200), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(G20), .A3(new_n291), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  AOI211_X1 g0541(.A(new_n265), .B(new_n738), .C1(G329), .C2(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n225), .B1(new_n739), .B2(G190), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n743), .A2(KEYINPUT102), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(KEYINPUT102), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n734), .A2(new_n291), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(G200), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n747), .A2(G294), .B1(new_n749), .B2(G311), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n291), .A2(new_n327), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n734), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g0553(.A(new_n742), .B(new_n750), .C1(new_n751), .C2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(G283), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n288), .A2(G179), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT99), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n757), .A2(new_n225), .A3(G190), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NOR3_X1   g0559(.A1(new_n757), .A2(new_n225), .A3(new_n291), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  OAI22_X1  g0561(.A1(new_n755), .A2(new_n759), .B1(new_n761), .B2(new_n587), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n734), .A2(new_n291), .A3(G200), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(KEYINPUT101), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n763), .A2(KEYINPUT101), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XNOR2_X1  g0568(.A(KEYINPUT33), .B(G317), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n754), .B(new_n762), .C1(new_n768), .C2(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n758), .A2(G107), .ZN(new_n771));
  OAI211_X1 g0571(.A(new_n771), .B(new_n265), .C1(new_n761), .C2(new_n534), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT100), .Z(new_n773));
  NOR2_X1   g0573(.A1(new_n746), .A2(new_n205), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n774), .B1(G77), .B2(new_n749), .ZN(new_n775));
  INV_X1    g0575(.A(new_n753), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT32), .ZN(new_n777));
  INV_X1    g0577(.A(G159), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n740), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n741), .A2(KEYINPUT32), .A3(G159), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n776), .A2(G50), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  OAI211_X1 g0581(.A(new_n775), .B(new_n781), .C1(new_n382), .C2(new_n736), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n782), .B1(G68), .B2(new_n768), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n770), .B1(new_n773), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n730), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n718), .B(new_n732), .C1(new_n784), .C2(new_n785), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n654), .A2(new_n721), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n653), .A2(G330), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(G396));
  NAND2_X1  g0589(.A1(new_n314), .A2(new_n650), .ZN(new_n790));
  MUX2_X1   g0590(.A(new_n300), .B(new_n650), .S(new_n310), .Z(new_n791));
  OAI21_X1  g0591(.A(new_n790), .B1(new_n791), .B2(new_n314), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n641), .A2(new_n650), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  AOI21_X1  g0595(.A(new_n793), .B1(new_n641), .B2(new_n650), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n720), .B1(new_n797), .B2(new_n710), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n710), .B2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n730), .A2(new_n715), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n720), .B1(G77), .B2(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT103), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n758), .A2(G68), .ZN(new_n804));
  INV_X1    g0604(.A(G132), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n265), .B1(new_n740), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(new_n747), .B2(G58), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n804), .B(new_n807), .C1(new_n761), .C2(new_n202), .ZN(new_n808));
  INV_X1    g0608(.A(new_n736), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n776), .B1(new_n809), .B2(G143), .ZN(new_n810));
  INV_X1    g0610(.A(new_n749), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n778), .B2(new_n811), .C1(new_n767), .C2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT34), .ZN(new_n814));
  AOI21_X1  g0614(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n265), .B1(new_n741), .B2(G311), .ZN(new_n817));
  INV_X1    g0617(.A(G294), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n817), .B1(new_n736), .B2(new_n818), .C1(new_n587), .C2(new_n753), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n774), .B(new_n819), .C1(G116), .C2(new_n749), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n768), .A2(G283), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n758), .A2(G87), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n760), .A2(G107), .ZN(new_n823));
  NAND4_X1  g0623(.A1(new_n820), .A2(new_n821), .A3(new_n822), .A4(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n816), .A2(new_n824), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n803), .B1(new_n825), .B2(new_n785), .C1(new_n793), .C2(new_n716), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n799), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G384));
  NAND2_X1  g0628(.A1(new_n463), .A2(new_n466), .ZN(new_n829));
  OAI211_X1 g0629(.A(G116), .B(new_n226), .C1(new_n829), .C2(KEYINPUT35), .ZN(new_n830));
  INV_X1    g0630(.A(KEYINPUT104), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n830), .A2(new_n831), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n829), .A2(KEYINPUT35), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n832), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  OR3_X1    g0636(.A1(new_n229), .A2(new_n267), .A3(new_n383), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n202), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n258), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n794), .A2(new_n790), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n402), .A2(new_n407), .ZN(new_n843));
  INV_X1    g0643(.A(new_n647), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n402), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT37), .ZN(new_n846));
  NAND4_X1  g0646(.A1(new_n843), .A2(new_n845), .A3(new_n846), .A4(new_n395), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  AOI21_X1  g0648(.A(KEYINPUT16), .B1(new_n392), .B2(new_n387), .ZN(new_n849));
  OAI21_X1  g0649(.A(KEYINPUT106), .B1(new_n849), .B2(new_n411), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT106), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n256), .C1(new_n414), .C2(KEYINPUT16), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n850), .A2(new_n393), .A3(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n406), .B1(new_n853), .B2(new_n351), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n853), .A2(new_n351), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n844), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n855), .A2(new_n857), .A3(new_n395), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n848), .B1(new_n858), .B2(KEYINPUT37), .ZN(new_n859));
  INV_X1    g0659(.A(new_n395), .ZN(new_n860));
  INV_X1    g0660(.A(KEYINPUT17), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI211_X1 g0662(.A(KEYINPUT75), .B(new_n861), .C1(new_n419), .C2(new_n368), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n399), .B1(new_n395), .B2(KEYINPUT17), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n862), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n421), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n857), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n842), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n647), .B1(new_n853), .B2(new_n351), .ZN(new_n869));
  NOR3_X1   g0669(.A1(new_n854), .A2(new_n869), .A3(new_n860), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n847), .B1(new_n870), .B2(new_n846), .ZN(new_n871));
  OAI21_X1  g0671(.A(new_n869), .B1(new_n401), .B2(new_n421), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n871), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n428), .A2(KEYINPUT105), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT105), .ZN(new_n876));
  OAI211_X1 g0676(.A(new_n876), .B(new_n346), .C1(new_n426), .C2(new_n427), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n346), .A2(new_n649), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n875), .A2(new_n348), .A3(new_n877), .A4(new_n878), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n613), .A2(new_n649), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n841), .A2(new_n874), .A3(new_n881), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n612), .A2(new_n844), .ZN(new_n883));
  INV_X1    g0683(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT107), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n874), .A2(KEYINPUT39), .ZN(new_n888));
  INV_X1    g0688(.A(KEYINPUT109), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n843), .A2(new_n845), .A3(new_n395), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(KEYINPUT37), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(new_n847), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT108), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n398), .A2(new_n400), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n894), .B1(new_n895), .B2(new_n862), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n894), .B(new_n862), .C1(new_n863), .C2(new_n864), .ZN(new_n897));
  INV_X1    g0697(.A(new_n897), .ZN(new_n898));
  OAI21_X1  g0698(.A(new_n612), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n845), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n893), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n889), .B1(new_n901), .B2(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n865), .A2(KEYINPUT108), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n903), .A2(new_n897), .ZN(new_n904));
  AOI21_X1  g0704(.A(new_n845), .B1(new_n904), .B2(new_n612), .ZN(new_n905));
  OAI211_X1 g0705(.A(KEYINPUT109), .B(new_n842), .C1(new_n905), .C2(new_n893), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n902), .A2(new_n873), .A3(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n888), .B1(new_n907), .B2(KEYINPUT39), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n649), .B1(new_n875), .B2(new_n877), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n882), .A2(KEYINPUT107), .A3(new_n884), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n887), .A2(new_n910), .A3(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n676), .A2(new_n429), .A3(new_n682), .ZN(new_n913));
  AND2_X1   g0713(.A1(new_n913), .A2(new_n616), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n912), .B(new_n914), .Z(new_n915));
  NAND3_X1  g0715(.A1(new_n702), .A2(KEYINPUT31), .A3(new_n649), .ZN(new_n916));
  NAND4_X1  g0716(.A1(new_n685), .A2(new_n707), .A3(new_n705), .A4(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n792), .B1(new_n879), .B2(new_n880), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n874), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT40), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(KEYINPUT110), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n919), .A2(KEYINPUT110), .A3(new_n920), .ZN(new_n924));
  AND3_X1   g0724(.A1(new_n917), .A2(KEYINPUT40), .A3(new_n918), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n923), .A2(new_n924), .B1(new_n907), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n926), .A2(new_n429), .A3(new_n917), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(G330), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n429), .B2(new_n917), .ZN(new_n929));
  OR2_X1    g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n915), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n258), .B2(new_n719), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n915), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n840), .B1(new_n932), .B2(new_n933), .ZN(G367));
  INV_X1    g0734(.A(KEYINPUT113), .ZN(new_n935));
  INV_X1    g0735(.A(new_n489), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n496), .B1(new_n936), .B2(new_n650), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n632), .A2(new_n649), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n664), .A2(new_n939), .A3(new_n661), .ZN(new_n940));
  XOR2_X1   g0740(.A(new_n940), .B(KEYINPUT42), .Z(new_n941));
  XOR2_X1   g0741(.A(new_n939), .B(KEYINPUT111), .Z(new_n942));
  AOI21_X1  g0742(.A(new_n632), .B1(new_n942), .B2(new_n608), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n941), .B1(new_n943), .B2(new_n649), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n619), .A2(new_n621), .A3(new_n649), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n635), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n946), .B1(new_n677), .B2(new_n945), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n947), .B(KEYINPUT43), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n949), .A2(KEYINPUT112), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT112), .ZN(new_n951));
  NAND3_X1  g0751(.A1(new_n944), .A2(new_n951), .A3(new_n948), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n947), .A2(KEYINPUT43), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n944), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n935), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  AOI211_X1 g0758(.A(KEYINPUT113), .B(new_n956), .C1(new_n950), .C2(new_n952), .ZN(new_n959));
  INV_X1    g0759(.A(new_n942), .ZN(new_n960));
  OAI22_X1  g0760(.A1(new_n958), .A2(new_n959), .B1(new_n662), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n952), .ZN(new_n962));
  AOI21_X1  g0762(.A(new_n951), .B1(new_n944), .B2(new_n948), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n957), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n964), .A2(KEYINPUT113), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n953), .A2(new_n935), .A3(new_n957), .ZN(new_n966));
  INV_X1    g0766(.A(new_n662), .ZN(new_n967));
  NAND4_X1  g0767(.A1(new_n965), .A2(new_n966), .A3(new_n967), .A4(new_n942), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n719), .A2(G45), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(G1), .ZN(new_n970));
  INV_X1    g0770(.A(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n939), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n666), .A2(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT44), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n973), .B(new_n974), .ZN(new_n975));
  NAND3_X1  g0775(.A1(new_n667), .A2(KEYINPUT45), .A3(new_n939), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT45), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n666), .B2(new_n972), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n967), .A2(KEYINPUT114), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n975), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n975), .B2(new_n979), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n664), .B(new_n661), .ZN(new_n984));
  XNOR2_X1  g0784(.A(new_n984), .B(new_n654), .ZN(new_n985));
  INV_X1    g0785(.A(new_n985), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n983), .A2(new_n986), .B1(new_n712), .B2(new_n711), .ZN(new_n987));
  XOR2_X1   g0787(.A(new_n669), .B(KEYINPUT41), .Z(new_n988));
  OAI21_X1  g0788(.A(new_n971), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g0789(.A1(new_n961), .A2(new_n968), .A3(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n731), .B1(new_n241), .B2(new_n728), .ZN(new_n991));
  INV_X1    g0791(.A(KEYINPUT68), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n303), .B(new_n992), .ZN(new_n993));
  AOI21_X1  g0793(.A(new_n991), .B1(new_n221), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(KEYINPUT115), .B(G317), .Z(new_n995));
  INV_X1    g0795(.A(G311), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n389), .B1(new_n740), .B2(new_n995), .C1(new_n753), .C2(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G303), .B2(new_n809), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n747), .A2(G107), .B1(new_n749), .B2(G283), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n759), .C2(new_n540), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT46), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n761), .B2(new_n573), .ZN(new_n1002));
  NAND3_X1  g0802(.A1(new_n760), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1003));
  OAI211_X1 g0803(.A(new_n1002), .B(new_n1003), .C1(new_n818), .C2(new_n767), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n746), .A2(new_n333), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n389), .B1(new_n741), .B2(G137), .ZN(new_n1006));
  INV_X1    g0806(.A(G143), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n736), .B2(new_n812), .C1(new_n1007), .C2(new_n753), .ZN(new_n1008));
  AOI211_X1 g0808(.A(new_n1005), .B(new_n1008), .C1(G50), .C2(new_n749), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n758), .A2(G77), .ZN(new_n1010));
  OAI211_X1 g0810(.A(new_n1009), .B(new_n1010), .C1(new_n382), .C2(new_n761), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n767), .A2(new_n778), .ZN(new_n1012));
  OAI22_X1  g0812(.A1(new_n1000), .A2(new_n1004), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(KEYINPUT116), .B(KEYINPUT47), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n785), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n721), .B(new_n994), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n717), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n947), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n990), .A2(new_n1019), .ZN(G387));
  NAND2_X1  g0820(.A1(new_n986), .A2(new_n970), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n661), .A2(new_n1018), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n728), .B1(new_n238), .B2(G45), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n1023), .B1(new_n672), .B2(new_n723), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n301), .A2(new_n202), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT50), .ZN(new_n1026));
  NOR2_X1   g0826(.A1(new_n333), .A2(new_n267), .ZN(new_n1027));
  NOR4_X1   g0827(.A1(new_n1026), .A2(G45), .A3(new_n1027), .A4(new_n672), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1024), .A2(new_n1028), .B1(G107), .B2(new_n220), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n721), .B1(new_n1029), .B2(new_n731), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n747), .A2(new_n993), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n809), .A2(G50), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n265), .B1(new_n740), .B2(new_n812), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1033), .B1(new_n776), .B2(G159), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n749), .A2(G68), .ZN(new_n1035));
  NAND4_X1  g0835(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OAI22_X1  g0836(.A1(new_n267), .A2(new_n761), .B1(new_n759), .B2(new_n205), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n1036), .B(new_n1037), .C1(new_n301), .C2(new_n768), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n389), .B1(new_n740), .B2(new_n751), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n776), .A2(G322), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n1040), .B1(new_n736), .B2(new_n995), .C1(new_n811), .C2(new_n587), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1041), .B1(new_n768), .B2(G311), .ZN(new_n1042));
  OR2_X1    g0842(.A1(new_n1042), .A2(KEYINPUT48), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1042), .A2(KEYINPUT48), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n760), .A2(G294), .B1(G283), .B2(new_n747), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1043), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT49), .ZN(new_n1047));
  NOR2_X1   g0847(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  AOI211_X1 g0848(.A(new_n1039), .B(new_n1048), .C1(G116), .C2(new_n758), .ZN(new_n1049));
  NAND2_X1  g0849(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1038), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1030), .B1(new_n1051), .B2(new_n785), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n713), .A2(new_n986), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n669), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n713), .A2(new_n986), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n1021), .B1(new_n1022), .B2(new_n1052), .C1(new_n1054), .C2(new_n1055), .ZN(G393));
  NOR2_X1   g0856(.A1(new_n248), .A2(new_n728), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n731), .B1(new_n220), .B2(new_n540), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n760), .A2(G283), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n747), .A2(G116), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n389), .B1(new_n740), .B2(new_n737), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n749), .B2(G294), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n771), .A2(new_n1059), .A3(new_n1060), .A4(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n1063), .ZN(new_n1064));
  AOI22_X1  g0864(.A1(G311), .A2(new_n809), .B1(new_n776), .B2(G317), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1065), .B(KEYINPUT52), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n768), .B2(G303), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n760), .A2(G68), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n749), .A2(new_n301), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n265), .B1(new_n740), .B2(new_n1007), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n1070), .B1(new_n747), .B2(G77), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n822), .A2(new_n1068), .A3(new_n1069), .A4(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(new_n1072), .ZN(new_n1073));
  OAI22_X1  g0873(.A1(new_n812), .A2(new_n753), .B1(new_n736), .B2(new_n778), .ZN(new_n1074));
  XOR2_X1   g0874(.A(new_n1074), .B(KEYINPUT51), .Z(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n768), .B2(G50), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(new_n1064), .A2(new_n1067), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n720), .B1(new_n1057), .B2(new_n1058), .C1(new_n1077), .C2(new_n785), .ZN(new_n1078));
  AOI21_X1  g0878(.A(new_n1078), .B1(new_n960), .B2(new_n717), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AND3_X1   g0880(.A1(new_n975), .A2(new_n967), .A3(new_n979), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n967), .B1(new_n975), .B2(new_n979), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1081), .A2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1080), .B1(new_n1083), .B2(new_n971), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1053), .ZN(new_n1085));
  AOI21_X1  g0885(.A(new_n670), .B1(new_n1085), .B2(new_n983), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1053), .A2(new_n1083), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(new_n1088), .ZN(G390));
  OR2_X1    g0889(.A1(new_n791), .A2(new_n314), .ZN(new_n1090));
  OAI211_X1 g0890(.A(new_n650), .B(new_n1090), .C1(new_n680), .C2(new_n681), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n790), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n909), .B1(new_n1092), .B2(new_n881), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n907), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n881), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(new_n794), .B2(new_n790), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1096), .A2(new_n909), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1094), .B1(new_n908), .B2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n917), .A2(G330), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(new_n918), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1098), .A2(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n710), .A2(new_n918), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1094), .B(new_n1104), .C1(new_n908), .C2(new_n1097), .ZN(new_n1105));
  NAND3_X1  g0905(.A1(new_n1103), .A2(new_n970), .A3(new_n1105), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT118), .Z(new_n1107));
  NAND2_X1  g0907(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1108));
  OAI21_X1  g0908(.A(KEYINPUT117), .B1(new_n617), .B2(new_n1099), .ZN(new_n1109));
  INV_X1    g0909(.A(KEYINPUT117), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1100), .A2(new_n1110), .A3(new_n429), .ZN(new_n1111));
  NAND4_X1  g0911(.A1(new_n913), .A2(new_n1109), .A3(new_n616), .A4(new_n1111), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n881), .B1(new_n710), .B2(new_n793), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n841), .B1(new_n1102), .B2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1095), .B1(new_n1099), .B2(new_n792), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n1104), .A2(new_n1115), .A3(new_n790), .A4(new_n1091), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1112), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1108), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1103), .A2(new_n1105), .A3(new_n1117), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1119), .A2(new_n669), .A3(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n720), .B1(new_n301), .B2(new_n801), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n760), .A2(G150), .ZN(new_n1123));
  XOR2_X1   g0923(.A(new_n1123), .B(KEYINPUT53), .Z(new_n1124));
  INV_X1    g0924(.A(G128), .ZN(new_n1125));
  NOR2_X1   g0925(.A1(new_n753), .A2(new_n1125), .ZN(new_n1126));
  AOI211_X1 g0926(.A(new_n389), .B(new_n1126), .C1(G125), .C2(new_n741), .ZN(new_n1127));
  XNOR2_X1  g0927(.A(KEYINPUT54), .B(G143), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n747), .A2(G159), .B1(new_n749), .B2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1127), .B(new_n1130), .C1(new_n805), .C2(new_n736), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G50), .B2(new_n758), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n768), .A2(G137), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1124), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n804), .B1(new_n818), .B2(new_n740), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT120), .ZN(new_n1136));
  AOI22_X1  g0936(.A1(G116), .A2(new_n809), .B1(new_n776), .B2(G283), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1137), .B1(new_n267), .B2(new_n746), .C1(new_n540), .C2(new_n811), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(new_n768), .B2(G107), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n265), .B1(new_n760), .B2(G87), .ZN(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT119), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1134), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1122), .B1(new_n1143), .B2(new_n730), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n908), .B2(new_n716), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1107), .A2(new_n1121), .A3(new_n1145), .ZN(G378));
  NAND2_X1  g0946(.A1(new_n923), .A2(new_n924), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n906), .A2(new_n873), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT90), .ZN(new_n1149));
  XNOR2_X1  g0949(.A(new_n421), .B(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(new_n903), .B2(new_n897), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n892), .B1(new_n1151), .B2(new_n845), .ZN(new_n1152));
  AOI21_X1  g0952(.A(KEYINPUT109), .B1(new_n1152), .B2(new_n842), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n925), .B1(new_n1148), .B2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n293), .A2(new_n285), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n264), .A2(new_n844), .ZN(new_n1156));
  XNOR2_X1  g0956(.A(new_n1155), .B(new_n1156), .ZN(new_n1157));
  XOR2_X1   g0957(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1159), .ZN(new_n1160));
  NAND4_X1  g0960(.A1(new_n1147), .A2(G330), .A3(new_n1154), .A4(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1160), .B1(new_n926), .B2(G330), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n912), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1164), .A2(KEYINPUT124), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n924), .ZN(new_n1166));
  AOI21_X1  g0966(.A(KEYINPUT110), .B1(new_n919), .B2(new_n920), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1154), .B(G330), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(new_n1159), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n886), .B(new_n883), .C1(new_n1096), .C2(new_n874), .ZN(new_n1170));
  AOI21_X1  g0970(.A(KEYINPUT107), .B1(new_n882), .B2(new_n884), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1169), .A2(new_n1172), .A3(new_n910), .A4(new_n1161), .ZN(new_n1173));
  INV_X1    g0973(.A(KEYINPUT124), .ZN(new_n1174));
  OAI211_X1 g0974(.A(new_n1174), .B(new_n912), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1165), .A2(new_n1173), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g0976(.A(KEYINPUT57), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n1112), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1177), .B1(new_n1120), .B2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n670), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1164), .A2(KEYINPUT122), .A3(new_n1173), .ZN(new_n1181));
  INV_X1    g0981(.A(KEYINPUT122), .ZN(new_n1182));
  OAI211_X1 g0982(.A(new_n1182), .B(new_n912), .C1(new_n1162), .C2(new_n1163), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1120), .A2(new_n1178), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1181), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n1177), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1180), .A2(new_n1186), .ZN(new_n1187));
  NAND3_X1  g0987(.A1(new_n1181), .A2(new_n970), .A3(new_n1183), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n721), .B1(new_n202), .B2(new_n800), .ZN(new_n1189));
  INV_X1    g0989(.A(G125), .ZN(new_n1190));
  OAI22_X1  g0990(.A1(new_n1190), .A2(new_n753), .B1(new_n736), .B2(new_n1125), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n746), .A2(new_n812), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n1191), .B(new_n1192), .C1(G137), .C2(new_n749), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n761), .B2(new_n1128), .C1(new_n767), .C2(new_n805), .ZN(new_n1194));
  OR2_X1    g0994(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1194), .A2(KEYINPUT59), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n758), .A2(G159), .ZN(new_n1197));
  AOI211_X1 g0997(.A(G33), .B(G41), .C1(new_n741), .C2(G124), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1195), .A2(new_n1196), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n389), .A2(new_n363), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n1200), .B1(G283), .B2(new_n741), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1201), .B1(new_n736), .B2(new_n206), .C1(new_n573), .C2(new_n753), .ZN(new_n1202));
  AOI211_X1 g1002(.A(new_n1005), .B(new_n1202), .C1(new_n993), .C2(new_n749), .ZN(new_n1203));
  AOI22_X1  g1003(.A1(G58), .A2(new_n758), .B1(new_n760), .B2(G77), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1203), .B(new_n1204), .C1(new_n205), .C2(new_n767), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1205), .ZN(new_n1206));
  OR2_X1    g1006(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1206), .A2(KEYINPUT58), .ZN(new_n1208));
  OAI211_X1 g1008(.A(new_n1200), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1209));
  AND4_X1   g1009(.A1(new_n1199), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1189), .B1(new_n785), .B2(new_n1210), .C1(new_n1160), .C2(new_n716), .ZN(new_n1211));
  XNOR2_X1  g1011(.A(new_n1211), .B(KEYINPUT121), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1188), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(KEYINPUT123), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1213), .A2(new_n1214), .ZN(new_n1215));
  AND2_X1   g1015(.A1(new_n1187), .A2(new_n1215), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1188), .A2(KEYINPUT123), .A3(new_n1212), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1216), .A2(new_n1217), .ZN(G375));
  AOI22_X1  g1018(.A1(new_n747), .A2(G50), .B1(new_n749), .B2(G150), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n265), .B1(new_n740), .B2(new_n1125), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n809), .B2(G137), .ZN(new_n1221));
  OAI211_X1 g1021(.A(new_n1219), .B(new_n1221), .C1(new_n805), .C2(new_n753), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n382), .A2(new_n759), .B1(new_n761), .B2(new_n778), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1222), .B(new_n1223), .C1(new_n768), .C2(new_n1129), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n389), .B1(new_n587), .B2(new_n740), .C1(new_n736), .C2(new_n755), .ZN(new_n1225));
  AOI21_X1  g1025(.A(new_n1225), .B1(G294), .B2(new_n776), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1226), .B(new_n1031), .C1(new_n206), .C2(new_n811), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1010), .B1(new_n761), .B2(new_n205), .ZN(new_n1228));
  AOI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(G116), .C2(new_n768), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n730), .B1(new_n1224), .B2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n721), .B1(new_n333), .B2(new_n800), .ZN(new_n1231));
  OAI211_X1 g1031(.A(new_n1230), .B(new_n1231), .C1(new_n881), .C2(new_n716), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1233), .B1(new_n1234), .B2(new_n970), .ZN(new_n1235));
  XOR2_X1   g1035(.A(new_n988), .B(KEYINPUT125), .Z(new_n1236));
  NAND2_X1  g1036(.A1(new_n1118), .A2(new_n1236), .ZN(new_n1237));
  NOR2_X1   g1037(.A1(new_n1234), .A2(new_n1178), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1235), .B1(new_n1237), .B2(new_n1238), .ZN(G381));
  AND3_X1   g1039(.A1(new_n1107), .A2(new_n1121), .A3(new_n1145), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1216), .A2(new_n1240), .A3(new_n1217), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n990), .A2(new_n1019), .A3(new_n1088), .ZN(new_n1242));
  OR3_X1    g1042(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1243));
  OR4_X1    g1043(.A1(G381), .A2(new_n1241), .A3(new_n1242), .A4(new_n1243), .ZN(G407));
  OAI211_X1 g1044(.A(G407), .B(G213), .C1(G343), .C2(new_n1241), .ZN(G409));
  NAND2_X1  g1045(.A1(G387), .A2(G390), .ZN(new_n1246));
  XNOR2_X1  g1046(.A(G393), .B(G396), .ZN(new_n1247));
  AND3_X1   g1047(.A1(new_n1246), .A2(new_n1242), .A3(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1247), .B1(new_n1246), .B2(new_n1242), .ZN(new_n1249));
  NOR2_X1   g1049(.A1(new_n1248), .A2(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1250), .ZN(new_n1251));
  NAND4_X1  g1051(.A1(new_n1187), .A2(new_n1215), .A3(G378), .A4(new_n1217), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1176), .A2(new_n970), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1236), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1253), .B(new_n1212), .C1(new_n1185), .C2(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1240), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1252), .A2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n648), .A2(G213), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1238), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1259), .A2(KEYINPUT60), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(new_n1259), .A2(KEYINPUT60), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n669), .B(new_n1118), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n1235), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1263), .A2(new_n827), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(G384), .A3(new_n1235), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1257), .A2(new_n1258), .A3(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(KEYINPUT126), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  NAND4_X1  g1070(.A1(new_n1257), .A2(KEYINPUT126), .A3(new_n1258), .A4(new_n1267), .ZN(new_n1271));
  AOI21_X1  g1071(.A(KEYINPUT62), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n648), .A2(G213), .A3(G2897), .ZN(new_n1274));
  AND3_X1   g1074(.A1(new_n1264), .A2(new_n1265), .A3(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1274), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1276));
  NOR2_X1   g1076(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT61), .B1(new_n1273), .B2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1268), .A2(KEYINPUT62), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1251), .B1(new_n1272), .B2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT63), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1270), .A2(new_n1282), .A3(new_n1271), .ZN(new_n1283));
  OR2_X1    g1083(.A1(new_n1268), .A2(new_n1282), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1283), .A2(new_n1284), .A3(new_n1278), .A4(new_n1250), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1281), .A2(new_n1285), .ZN(G405));
  NAND2_X1  g1086(.A1(G375), .A2(G378), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1287), .A2(new_n1241), .ZN(new_n1288));
  INV_X1    g1088(.A(KEYINPUT127), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1288), .A2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1266), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1247), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1242), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1088), .B1(new_n990), .B2(new_n1019), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1292), .B1(new_n1293), .B2(new_n1294), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1246), .A2(new_n1242), .A3(new_n1247), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1295), .A2(new_n1267), .A3(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1291), .A2(new_n1297), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1287), .A2(KEYINPUT127), .A3(new_n1241), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1290), .A2(new_n1298), .A3(new_n1299), .ZN(new_n1300));
  AOI21_X1  g1100(.A(new_n1298), .B1(new_n1290), .B2(new_n1299), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(G402));
endmodule


