

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586;

  XNOR2_X1 U321 ( .A(n405), .B(n404), .ZN(n406) );
  NOR2_X1 U322 ( .A1(n469), .A2(n468), .ZN(n471) );
  XNOR2_X1 U323 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U324 ( .A(n467), .B(n466), .ZN(n573) );
  XNOR2_X1 U325 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n466) );
  XNOR2_X1 U326 ( .A(n411), .B(n410), .ZN(n523) );
  XNOR2_X1 U327 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U328 ( .A(n401), .B(n400), .Z(n289) );
  XOR2_X1 U329 ( .A(G218GAT), .B(G106GAT), .Z(n290) );
  XOR2_X1 U330 ( .A(KEYINPUT2), .B(KEYINPUT3), .Z(n291) );
  AND2_X1 U331 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  INV_X1 U332 ( .A(KEYINPUT97), .ZN(n462) );
  XNOR2_X1 U333 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U334 ( .A(n465), .B(n464), .ZN(n469) );
  INV_X1 U335 ( .A(KEYINPUT98), .ZN(n470) );
  XNOR2_X1 U336 ( .A(n381), .B(KEYINPUT112), .ZN(n382) );
  XNOR2_X1 U337 ( .A(n383), .B(n382), .ZN(n394) );
  XNOR2_X1 U338 ( .A(n437), .B(n292), .ZN(n438) );
  XNOR2_X1 U339 ( .A(n327), .B(n326), .ZN(n328) );
  INV_X1 U340 ( .A(KEYINPUT92), .ZN(n404) );
  XNOR2_X1 U341 ( .A(n347), .B(KEYINPUT33), .ZN(n348) );
  XNOR2_X1 U342 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U343 ( .A(n444), .B(n290), .ZN(n445) );
  NOR2_X1 U344 ( .A1(n479), .A2(n478), .ZN(n490) );
  XNOR2_X1 U345 ( .A(n362), .B(n348), .ZN(n352) );
  XNOR2_X1 U346 ( .A(n451), .B(KEYINPUT55), .ZN(n452) );
  XNOR2_X1 U347 ( .A(n446), .B(n445), .ZN(n450) );
  XNOR2_X1 U348 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U349 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U350 ( .A(n358), .B(n357), .ZN(n578) );
  XNOR2_X1 U351 ( .A(n509), .B(KEYINPUT105), .ZN(n515) );
  XNOR2_X1 U352 ( .A(n309), .B(n410), .ZN(n533) );
  XNOR2_X1 U353 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U354 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n483) );
  XNOR2_X1 U355 ( .A(n458), .B(n457), .ZN(G1351GAT) );
  XNOR2_X1 U356 ( .A(n484), .B(n483), .ZN(G1328GAT) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(G190GAT), .ZN(n293) );
  XNOR2_X1 U358 ( .A(n293), .B(G134GAT), .ZN(n314) );
  XOR2_X1 U359 ( .A(n314), .B(KEYINPUT79), .Z(n295) );
  NAND2_X1 U360 ( .A1(G227GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U361 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U362 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n297) );
  XNOR2_X1 U363 ( .A(G15GAT), .B(G99GAT), .ZN(n296) );
  XNOR2_X1 U364 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U365 ( .A(n299), .B(n298), .Z(n304) );
  XNOR2_X1 U366 ( .A(G176GAT), .B(G71GAT), .ZN(n300) );
  XNOR2_X1 U367 ( .A(n300), .B(G120GAT), .ZN(n354) );
  XOR2_X1 U368 ( .A(KEYINPUT77), .B(KEYINPUT0), .Z(n302) );
  XNOR2_X1 U369 ( .A(G113GAT), .B(G127GAT), .ZN(n301) );
  XNOR2_X1 U370 ( .A(n302), .B(n301), .ZN(n428) );
  XNOR2_X1 U371 ( .A(n354), .B(n428), .ZN(n303) );
  XNOR2_X1 U372 ( .A(n304), .B(n303), .ZN(n309) );
  XOR2_X1 U373 ( .A(KEYINPUT80), .B(G183GAT), .Z(n306) );
  XNOR2_X1 U374 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n305) );
  XNOR2_X1 U375 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U376 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n307) );
  XNOR2_X1 U377 ( .A(n308), .B(n307), .ZN(n410) );
  XOR2_X1 U378 ( .A(KEYINPUT66), .B(G106GAT), .Z(n311) );
  XNOR2_X1 U379 ( .A(G99GAT), .B(G92GAT), .ZN(n310) );
  XNOR2_X1 U380 ( .A(n311), .B(n310), .ZN(n312) );
  XOR2_X1 U381 ( .A(G85GAT), .B(n312), .Z(n356) );
  XNOR2_X1 U382 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n313) );
  XNOR2_X1 U383 ( .A(n313), .B(KEYINPUT7), .ZN(n341) );
  XNOR2_X1 U384 ( .A(n314), .B(n341), .ZN(n320) );
  INV_X1 U385 ( .A(n320), .ZN(n318) );
  XNOR2_X1 U386 ( .A(KEYINPUT70), .B(KEYINPUT11), .ZN(n316) );
  AND2_X1 U387 ( .A1(G232GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U388 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U389 ( .A(n317), .B(KEYINPUT72), .ZN(n319) );
  NAND2_X1 U390 ( .A1(n318), .A2(n319), .ZN(n323) );
  INV_X1 U391 ( .A(n319), .ZN(n321) );
  NAND2_X1 U392 ( .A1(n321), .A2(n320), .ZN(n322) );
  NAND2_X1 U393 ( .A1(n323), .A2(n322), .ZN(n329) );
  XOR2_X1 U394 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n325) );
  XNOR2_X1 U395 ( .A(KEYINPUT69), .B(KEYINPUT9), .ZN(n324) );
  XOR2_X1 U396 ( .A(n325), .B(n324), .Z(n327) );
  XOR2_X1 U397 ( .A(G36GAT), .B(G218GAT), .Z(n401) );
  XOR2_X1 U398 ( .A(G50GAT), .B(G162GAT), .Z(n437) );
  XNOR2_X1 U399 ( .A(n401), .B(n437), .ZN(n326) );
  XNOR2_X1 U400 ( .A(n356), .B(n330), .ZN(n384) );
  XOR2_X1 U401 ( .A(G36GAT), .B(G50GAT), .Z(n332) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n331) );
  XNOR2_X1 U403 ( .A(n332), .B(n331), .ZN(n345) );
  XOR2_X1 U404 ( .A(G22GAT), .B(G113GAT), .Z(n334) );
  XNOR2_X1 U405 ( .A(KEYINPUT29), .B(G141GAT), .ZN(n333) );
  XNOR2_X1 U406 ( .A(n334), .B(n333), .ZN(n338) );
  XOR2_X1 U407 ( .A(KEYINPUT30), .B(G197GAT), .Z(n336) );
  XNOR2_X1 U408 ( .A(G169GAT), .B(G43GAT), .ZN(n335) );
  XNOR2_X1 U409 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U410 ( .A(n338), .B(n337), .Z(n343) );
  XOR2_X1 U411 ( .A(G1GAT), .B(G15GAT), .Z(n340) );
  XNOR2_X1 U412 ( .A(G8GAT), .B(KEYINPUT65), .ZN(n339) );
  XNOR2_X1 U413 ( .A(n340), .B(n339), .ZN(n365) );
  XNOR2_X1 U414 ( .A(n341), .B(n365), .ZN(n342) );
  XNOR2_X1 U415 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U416 ( .A(n345), .B(n344), .Z(n575) );
  INV_X1 U417 ( .A(n575), .ZN(n551) );
  XNOR2_X1 U418 ( .A(G57GAT), .B(G64GAT), .ZN(n346) );
  XNOR2_X1 U419 ( .A(n346), .B(KEYINPUT13), .ZN(n362) );
  AND2_X1 U420 ( .A1(G230GAT), .A2(G233GAT), .ZN(n347) );
  XOR2_X1 U421 ( .A(KEYINPUT68), .B(KEYINPUT31), .Z(n350) );
  XNOR2_X1 U422 ( .A(KEYINPUT32), .B(KEYINPUT67), .ZN(n349) );
  XOR2_X1 U423 ( .A(n350), .B(n349), .Z(n351) );
  XNOR2_X1 U424 ( .A(n352), .B(n351), .ZN(n358) );
  XNOR2_X1 U425 ( .A(G148GAT), .B(G204GAT), .ZN(n353) );
  XNOR2_X1 U426 ( .A(n353), .B(G78GAT), .ZN(n447) );
  XNOR2_X1 U427 ( .A(n354), .B(n447), .ZN(n355) );
  XNOR2_X1 U428 ( .A(KEYINPUT41), .B(n578), .ZN(n555) );
  NOR2_X1 U429 ( .A1(n551), .A2(n555), .ZN(n361) );
  XOR2_X1 U430 ( .A(KEYINPUT110), .B(KEYINPUT46), .Z(n359) );
  XNOR2_X1 U431 ( .A(KEYINPUT109), .B(n359), .ZN(n360) );
  XNOR2_X1 U432 ( .A(n361), .B(n360), .ZN(n378) );
  XOR2_X1 U433 ( .A(G22GAT), .B(G155GAT), .Z(n440) );
  XOR2_X1 U434 ( .A(n440), .B(n362), .Z(n364) );
  XNOR2_X1 U435 ( .A(G183GAT), .B(G211GAT), .ZN(n363) );
  XNOR2_X1 U436 ( .A(n364), .B(n363), .ZN(n369) );
  XOR2_X1 U437 ( .A(n365), .B(KEYINPUT12), .Z(n367) );
  NAND2_X1 U438 ( .A1(G231GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U439 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U440 ( .A(n369), .B(n368), .Z(n377) );
  XOR2_X1 U441 ( .A(KEYINPUT74), .B(KEYINPUT14), .Z(n371) );
  XNOR2_X1 U442 ( .A(KEYINPUT76), .B(KEYINPUT15), .ZN(n370) );
  XNOR2_X1 U443 ( .A(n371), .B(n370), .ZN(n375) );
  XOR2_X1 U444 ( .A(G78GAT), .B(KEYINPUT75), .Z(n373) );
  XNOR2_X1 U445 ( .A(G71GAT), .B(G127GAT), .ZN(n372) );
  XNOR2_X1 U446 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U448 ( .A(n377), .B(n376), .ZN(n581) );
  NOR2_X1 U449 ( .A1(n378), .A2(n581), .ZN(n379) );
  XNOR2_X1 U450 ( .A(n379), .B(KEYINPUT111), .ZN(n380) );
  NOR2_X1 U451 ( .A1(n384), .A2(n380), .ZN(n383) );
  INV_X1 U452 ( .A(KEYINPUT47), .ZN(n381) );
  INV_X1 U453 ( .A(KEYINPUT115), .ZN(n392) );
  INV_X1 U454 ( .A(n384), .ZN(n561) );
  XNOR2_X2 U455 ( .A(n561), .B(KEYINPUT73), .ZN(n544) );
  XNOR2_X1 U456 ( .A(KEYINPUT36), .B(n544), .ZN(n459) );
  NAND2_X1 U457 ( .A1(n459), .A2(n581), .ZN(n386) );
  XOR2_X1 U458 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n385) );
  XNOR2_X1 U459 ( .A(n386), .B(n385), .ZN(n387) );
  NOR2_X1 U460 ( .A1(n387), .A2(n578), .ZN(n389) );
  INV_X1 U461 ( .A(KEYINPUT114), .ZN(n388) );
  XNOR2_X1 U462 ( .A(n389), .B(n388), .ZN(n390) );
  NOR2_X1 U463 ( .A1(n575), .A2(n390), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n392), .B(n391), .ZN(n393) );
  NOR2_X1 U465 ( .A1(n394), .A2(n393), .ZN(n395) );
  XNOR2_X1 U466 ( .A(KEYINPUT48), .B(n395), .ZN(n531) );
  XOR2_X1 U467 ( .A(KEYINPUT90), .B(G64GAT), .Z(n397) );
  XNOR2_X1 U468 ( .A(KEYINPUT89), .B(G204GAT), .ZN(n396) );
  XNOR2_X1 U469 ( .A(n397), .B(n396), .ZN(n409) );
  XOR2_X1 U470 ( .A(KEYINPUT91), .B(G92GAT), .Z(n399) );
  XNOR2_X1 U471 ( .A(G8GAT), .B(G190GAT), .ZN(n398) );
  XNOR2_X1 U472 ( .A(n399), .B(n398), .ZN(n400) );
  NAND2_X1 U473 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U474 ( .A(n289), .B(n402), .ZN(n407) );
  XNOR2_X1 U475 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n403) );
  XNOR2_X1 U476 ( .A(n403), .B(G211GAT), .ZN(n448) );
  XNOR2_X1 U477 ( .A(G176GAT), .B(n448), .ZN(n405) );
  XNOR2_X1 U478 ( .A(n409), .B(n408), .ZN(n411) );
  NOR2_X1 U479 ( .A1(n531), .A2(n523), .ZN(n412) );
  XNOR2_X1 U480 ( .A(n412), .B(KEYINPUT54), .ZN(n435) );
  NAND2_X1 U481 ( .A1(G225GAT), .A2(G233GAT), .ZN(n418) );
  XOR2_X1 U482 ( .A(G57GAT), .B(G134GAT), .Z(n414) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G1GAT), .ZN(n413) );
  XNOR2_X1 U484 ( .A(n414), .B(n413), .ZN(n416) );
  XOR2_X1 U485 ( .A(G85GAT), .B(G162GAT), .Z(n415) );
  XNOR2_X1 U486 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U487 ( .A(n418), .B(n417), .ZN(n434) );
  XOR2_X1 U488 ( .A(KEYINPUT86), .B(KEYINPUT85), .Z(n420) );
  XNOR2_X1 U489 ( .A(KEYINPUT84), .B(KEYINPUT1), .ZN(n419) );
  XNOR2_X1 U490 ( .A(n420), .B(n419), .ZN(n432) );
  XOR2_X1 U491 ( .A(KEYINPUT88), .B(G148GAT), .Z(n422) );
  XNOR2_X1 U492 ( .A(G120GAT), .B(G155GAT), .ZN(n421) );
  XNOR2_X1 U493 ( .A(n422), .B(n421), .ZN(n426) );
  XOR2_X1 U494 ( .A(KEYINPUT87), .B(KEYINPUT4), .Z(n424) );
  XNOR2_X1 U495 ( .A(KEYINPUT6), .B(KEYINPUT5), .ZN(n423) );
  XNOR2_X1 U496 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U497 ( .A(n426), .B(n425), .Z(n430) );
  XNOR2_X1 U498 ( .A(G141GAT), .B(KEYINPUT83), .ZN(n427) );
  XNOR2_X1 U499 ( .A(n291), .B(n427), .ZN(n439) );
  XNOR2_X1 U500 ( .A(n428), .B(n439), .ZN(n429) );
  XNOR2_X1 U501 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U502 ( .A(n432), .B(n431), .Z(n433) );
  XNOR2_X1 U503 ( .A(n434), .B(n433), .ZN(n520) );
  NAND2_X1 U504 ( .A1(n435), .A2(n520), .ZN(n436) );
  XNOR2_X1 U505 ( .A(n436), .B(KEYINPUT64), .ZN(n574) );
  XOR2_X1 U506 ( .A(n441), .B(n440), .Z(n446) );
  XOR2_X1 U507 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n443) );
  XNOR2_X1 U508 ( .A(KEYINPUT82), .B(KEYINPUT24), .ZN(n442) );
  XNOR2_X1 U509 ( .A(n443), .B(n442), .ZN(n444) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U511 ( .A(n450), .B(n449), .ZN(n476) );
  NOR2_X1 U512 ( .A1(n574), .A2(n476), .ZN(n453) );
  INV_X1 U513 ( .A(KEYINPUT121), .ZN(n451) );
  NOR2_X2 U514 ( .A1(n533), .A2(n454), .ZN(n568) );
  NAND2_X1 U515 ( .A1(n568), .A2(n544), .ZN(n458) );
  XOR2_X1 U516 ( .A(KEYINPUT124), .B(KEYINPUT58), .Z(n456) );
  INV_X1 U517 ( .A(G190GAT), .ZN(n455) );
  NOR2_X1 U518 ( .A1(n551), .A2(n578), .ZN(n492) );
  NOR2_X1 U519 ( .A1(n533), .A2(n523), .ZN(n460) );
  XOR2_X1 U520 ( .A(KEYINPUT95), .B(n460), .Z(n461) );
  NOR2_X1 U521 ( .A1(n476), .A2(n461), .ZN(n465) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(KEYINPUT96), .Z(n463) );
  XNOR2_X1 U523 ( .A(KEYINPUT27), .B(n523), .ZN(n474) );
  NAND2_X1 U524 ( .A1(n476), .A2(n533), .ZN(n467) );
  NOR2_X1 U525 ( .A1(n474), .A2(n573), .ZN(n468) );
  XNOR2_X1 U526 ( .A(n471), .B(n470), .ZN(n472) );
  NAND2_X1 U527 ( .A1(n472), .A2(n520), .ZN(n473) );
  XNOR2_X1 U528 ( .A(n473), .B(KEYINPUT99), .ZN(n479) );
  NOR2_X1 U529 ( .A1(n520), .A2(n474), .ZN(n475) );
  XOR2_X1 U530 ( .A(KEYINPUT93), .B(n475), .Z(n550) );
  XOR2_X1 U531 ( .A(n476), .B(KEYINPUT28), .Z(n528) );
  NAND2_X1 U532 ( .A1(n550), .A2(n528), .ZN(n532) );
  XNOR2_X1 U533 ( .A(n533), .B(KEYINPUT81), .ZN(n477) );
  NOR2_X1 U534 ( .A1(n532), .A2(n477), .ZN(n478) );
  NOR2_X1 U535 ( .A1(n581), .A2(n490), .ZN(n480) );
  NAND2_X1 U536 ( .A1(n459), .A2(n480), .ZN(n481) );
  XNOR2_X1 U537 ( .A(KEYINPUT37), .B(n481), .ZN(n519) );
  NAND2_X1 U538 ( .A1(n492), .A2(n519), .ZN(n482) );
  XNOR2_X1 U539 ( .A(n482), .B(KEYINPUT38), .ZN(n506) );
  NOR2_X1 U540 ( .A1(n520), .A2(n506), .ZN(n484) );
  XOR2_X1 U541 ( .A(n555), .B(KEYINPUT104), .Z(n538) );
  NAND2_X1 U542 ( .A1(n538), .A2(n568), .ZN(n487) );
  XOR2_X1 U543 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n485) );
  XNOR2_X1 U544 ( .A(n485), .B(G176GAT), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1349GAT) );
  INV_X1 U546 ( .A(n581), .ZN(n559) );
  NOR2_X1 U547 ( .A1(n559), .A2(n544), .ZN(n488) );
  XOR2_X1 U548 ( .A(KEYINPUT16), .B(n488), .Z(n489) );
  NOR2_X1 U549 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U550 ( .A(KEYINPUT100), .B(n491), .ZN(n508) );
  NAND2_X1 U551 ( .A1(n492), .A2(n508), .ZN(n499) );
  NOR2_X1 U552 ( .A1(n520), .A2(n499), .ZN(n494) );
  XNOR2_X1 U553 ( .A(KEYINPUT34), .B(KEYINPUT101), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U555 ( .A(G1GAT), .B(n495), .ZN(G1324GAT) );
  NOR2_X1 U556 ( .A1(n523), .A2(n499), .ZN(n496) );
  XOR2_X1 U557 ( .A(G8GAT), .B(n496), .Z(G1325GAT) );
  NOR2_X1 U558 ( .A1(n533), .A2(n499), .ZN(n498) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(G1326GAT) );
  NOR2_X1 U561 ( .A1(n528), .A2(n499), .ZN(n500) );
  XOR2_X1 U562 ( .A(G22GAT), .B(n500), .Z(G1327GAT) );
  NOR2_X1 U563 ( .A1(n506), .A2(n523), .ZN(n501) );
  XOR2_X1 U564 ( .A(G36GAT), .B(n501), .Z(G1329GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n503) );
  XNOR2_X1 U566 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n502) );
  XNOR2_X1 U567 ( .A(n503), .B(n502), .ZN(n505) );
  NOR2_X1 U568 ( .A1(n533), .A2(n506), .ZN(n504) );
  XOR2_X1 U569 ( .A(n505), .B(n504), .Z(G1330GAT) );
  NOR2_X1 U570 ( .A1(n528), .A2(n506), .ZN(n507) );
  XOR2_X1 U571 ( .A(G50GAT), .B(n507), .Z(G1331GAT) );
  AND2_X1 U572 ( .A1(n538), .A2(n551), .ZN(n518) );
  AND2_X1 U573 ( .A1(n508), .A2(n518), .ZN(n509) );
  NOR2_X1 U574 ( .A1(n520), .A2(n515), .ZN(n510) );
  XOR2_X1 U575 ( .A(KEYINPUT42), .B(n510), .Z(n511) );
  XNOR2_X1 U576 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NOR2_X1 U577 ( .A1(n523), .A2(n515), .ZN(n512) );
  XOR2_X1 U578 ( .A(KEYINPUT106), .B(n512), .Z(n513) );
  XNOR2_X1 U579 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  NOR2_X1 U580 ( .A1(n533), .A2(n515), .ZN(n514) );
  XOR2_X1 U581 ( .A(G71GAT), .B(n514), .Z(G1334GAT) );
  NOR2_X1 U582 ( .A1(n528), .A2(n515), .ZN(n517) );
  XNOR2_X1 U583 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n516) );
  XNOR2_X1 U584 ( .A(n517), .B(n516), .ZN(G1335GAT) );
  NAND2_X1 U585 ( .A1(n519), .A2(n518), .ZN(n527) );
  NOR2_X1 U586 ( .A1(n520), .A2(n527), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G85GAT), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1336GAT) );
  NOR2_X1 U589 ( .A1(n523), .A2(n527), .ZN(n524) );
  XOR2_X1 U590 ( .A(KEYINPUT108), .B(n524), .Z(n525) );
  XNOR2_X1 U591 ( .A(G92GAT), .B(n525), .ZN(G1337GAT) );
  NOR2_X1 U592 ( .A1(n533), .A2(n527), .ZN(n526) );
  XOR2_X1 U593 ( .A(G99GAT), .B(n526), .Z(G1338GAT) );
  NOR2_X1 U594 ( .A1(n528), .A2(n527), .ZN(n529) );
  XOR2_X1 U595 ( .A(KEYINPUT44), .B(n529), .Z(n530) );
  XNOR2_X1 U596 ( .A(G106GAT), .B(n530), .ZN(G1339GAT) );
  NOR2_X1 U597 ( .A1(n531), .A2(n532), .ZN(n535) );
  INV_X1 U598 ( .A(n533), .ZN(n534) );
  NAND2_X1 U599 ( .A1(n535), .A2(n534), .ZN(n537) );
  NOR2_X1 U600 ( .A1(n551), .A2(n537), .ZN(n536) );
  XOR2_X1 U601 ( .A(G113GAT), .B(n536), .Z(G1340GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n540) );
  INV_X1 U603 ( .A(n537), .ZN(n545) );
  NAND2_X1 U604 ( .A1(n545), .A2(n538), .ZN(n539) );
  XNOR2_X1 U605 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n541), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n545), .A2(n581), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(KEYINPUT50), .ZN(n543) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n543), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT117), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U611 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U612 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U613 ( .A(G134GAT), .B(n548), .Z(G1343GAT) );
  NOR2_X1 U614 ( .A1(n531), .A2(n573), .ZN(n549) );
  NAND2_X1 U615 ( .A1(n550), .A2(n549), .ZN(n562) );
  NOR2_X1 U616 ( .A1(n551), .A2(n562), .ZN(n553) );
  XNOR2_X1 U617 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n552) );
  XNOR2_X1 U618 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U619 ( .A(G141GAT), .B(n554), .ZN(G1344GAT) );
  NOR2_X1 U620 ( .A1(n555), .A2(n562), .ZN(n557) );
  XNOR2_X1 U621 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n556) );
  XNOR2_X1 U622 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n558), .ZN(G1345GAT) );
  NOR2_X1 U624 ( .A1(n559), .A2(n562), .ZN(n560) );
  XOR2_X1 U625 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U626 ( .A1(n561), .A2(n562), .ZN(n563) );
  XOR2_X1 U627 ( .A(KEYINPUT120), .B(n563), .Z(n564) );
  XNOR2_X1 U628 ( .A(G162GAT), .B(n564), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n568), .A2(n575), .ZN(n566) );
  XOR2_X1 U630 ( .A(KEYINPUT122), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U631 ( .A(n566), .B(n565), .ZN(n567) );
  XNOR2_X1 U632 ( .A(n567), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n581), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U635 ( .A(KEYINPUT126), .B(KEYINPUT60), .Z(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n571), .B(n570), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(n572), .Z(n577) );
  NOR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n583) );
  NAND2_X1 U640 ( .A1(n583), .A2(n575), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n580) );
  NAND2_X1 U643 ( .A1(n583), .A2(n578), .ZN(n579) );
  XNOR2_X1 U644 ( .A(n580), .B(n579), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n583), .A2(n581), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U647 ( .A(KEYINPUT127), .B(KEYINPUT62), .Z(n585) );
  NAND2_X1 U648 ( .A1(n583), .A2(n459), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

