//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0 0 0 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n779,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n797, new_n798, new_n799, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n872, new_n873, new_n874, new_n875, new_n877, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n938, new_n939, new_n940, new_n941, new_n943, new_n944, new_n945,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT89), .B(G197gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XOR2_X1   g003(.A(KEYINPUT11), .B(G169gat), .Z(new_n205));
  XNOR2_X1  g004(.A(new_n204), .B(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(new_n206), .B(KEYINPUT12), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G15gat), .B(G22gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT91), .ZN(new_n210));
  INV_X1    g009(.A(G1gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(KEYINPUT91), .A3(G1gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT16), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n209), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(new_n213), .A3(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(G8gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(KEYINPUT14), .B(G29gat), .ZN(new_n219));
  INV_X1    g018(.A(G36gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G43gat), .B(G50gat), .ZN(new_n222));
  INV_X1    g021(.A(G29gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n223), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n224));
  NAND4_X1  g023(.A1(new_n221), .A2(KEYINPUT15), .A3(new_n222), .A4(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT90), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n222), .B(KEYINPUT15), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n221), .A2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n218), .A2(new_n226), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n226), .A2(new_n229), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n216), .B(G8gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n230), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G229gat), .A2(G233gat), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n235), .B(KEYINPUT13), .Z(new_n236));
  NAND2_X1  g035(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n231), .A2(KEYINPUT17), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT17), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n239), .B1(new_n226), .B2(new_n229), .ZN(new_n240));
  OR2_X1    g039(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n232), .B(KEYINPUT92), .ZN(new_n242));
  AOI22_X1  g041(.A1(new_n241), .A2(new_n242), .B1(new_n232), .B2(new_n231), .ZN(new_n243));
  AOI21_X1  g042(.A(KEYINPUT93), .B1(new_n243), .B2(new_n235), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT18), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n237), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n241), .A2(new_n242), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n235), .A3(new_n233), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT93), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n208), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n250), .A2(KEYINPUT18), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n244), .A2(new_n245), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n253), .A2(new_n254), .A3(new_n237), .A4(new_n207), .ZN(new_n255));
  AND2_X1   g054(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(G169gat), .ZN(new_n257));
  INV_X1    g056(.A(G176gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT69), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n259), .A2(KEYINPUT26), .ZN(new_n260));
  NAND2_X1  g059(.A1(G169gat), .A2(G176gat), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT65), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(KEYINPUT65), .A2(G169gat), .A3(G176gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(G169gat), .A2(G176gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT26), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n266), .A2(KEYINPUT69), .A3(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n265), .A3(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n270));
  INV_X1    g069(.A(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(G183gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT27), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT27), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n274), .A2(G183gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G190gat), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(KEYINPUT68), .B2(KEYINPUT28), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n271), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G183gat), .A2(G190gat), .ZN(new_n280));
  XNOR2_X1  g079(.A(KEYINPUT27), .B(G183gat), .ZN(new_n281));
  NOR2_X1   g080(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n282), .A2(G190gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n283), .A3(new_n270), .ZN(new_n284));
  NAND4_X1  g083(.A1(new_n269), .A2(new_n279), .A3(new_n280), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT70), .ZN(new_n286));
  INV_X1    g085(.A(new_n280), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n283), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n288), .B2(new_n271), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT70), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n289), .A2(new_n290), .A3(new_n269), .A4(new_n284), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n286), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT24), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n280), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g093(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n294), .B(new_n295), .C1(G183gat), .C2(G190gat), .ZN(new_n296));
  OR2_X1    g095(.A1(new_n266), .A2(KEYINPUT23), .ZN(new_n297));
  OR2_X1    g096(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n298));
  NAND2_X1  g097(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n298), .A2(KEYINPUT23), .A3(new_n257), .A4(new_n299), .ZN(new_n300));
  NAND4_X1  g099(.A1(new_n296), .A2(new_n265), .A3(new_n297), .A4(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT25), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(new_n264), .ZN(new_n304));
  AOI21_X1  g103(.A(KEYINPUT65), .B1(G169gat), .B2(G176gat), .ZN(new_n305));
  OAI22_X1  g104(.A1(new_n304), .A2(new_n305), .B1(KEYINPUT23), .B2(new_n266), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n257), .A2(new_n258), .A3(KEYINPUT23), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n307), .A2(KEYINPUT25), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT66), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n310), .A2(new_n311), .B1(new_n272), .B2(new_n277), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n294), .A2(KEYINPUT66), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n295), .A2(KEYINPUT67), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n312), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n309), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n303), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n292), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(G113gat), .ZN(new_n320));
  INV_X1    g119(.A(G120gat), .ZN(new_n321));
  AOI21_X1  g120(.A(KEYINPUT1), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n322), .B1(new_n320), .B2(new_n321), .ZN(new_n323));
  XNOR2_X1  g122(.A(G127gat), .B(G134gat), .ZN(new_n324));
  INV_X1    g123(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT71), .B(G113gat), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n322), .B(new_n324), .C1(new_n327), .C2(new_n321), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT72), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n329), .B1(new_n326), .B2(new_n328), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n319), .A2(new_n333), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n286), .A2(new_n291), .B1(new_n303), .B2(new_n317), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n335), .A2(new_n332), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n334), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(G227gat), .ZN(new_n338));
  INV_X1    g137(.A(G233gat), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g139(.A(KEYINPUT73), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  AND3_X1   g140(.A1(new_n292), .A2(new_n332), .A3(new_n318), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n332), .B1(new_n292), .B2(new_n318), .ZN(new_n343));
  OAI211_X1 g142(.A(KEYINPUT73), .B(new_n340), .C1(new_n342), .C2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT32), .B1(new_n341), .B2(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT33), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n347), .B1(new_n341), .B2(new_n345), .ZN(new_n348));
  XNOR2_X1  g147(.A(G15gat), .B(G43gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT76), .ZN(new_n350));
  XNOR2_X1  g149(.A(G71gat), .B(G99gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT74), .B(KEYINPUT75), .ZN(new_n353));
  XOR2_X1   g152(.A(new_n352), .B(new_n353), .Z(new_n354));
  NAND3_X1  g153(.A1(new_n346), .A2(new_n348), .A3(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT32), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n340), .B1(new_n342), .B2(new_n343), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT73), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n356), .B1(new_n359), .B2(new_n344), .ZN(new_n360));
  AOI21_X1  g159(.A(KEYINPUT33), .B1(new_n359), .B2(new_n344), .ZN(new_n361));
  INV_X1    g160(.A(new_n354), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n360), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT34), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n342), .A2(new_n343), .ZN(new_n365));
  INV_X1    g164(.A(new_n340), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n364), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NOR4_X1   g166(.A1(new_n342), .A2(new_n343), .A3(KEYINPUT34), .A4(new_n340), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AND3_X1   g168(.A1(new_n355), .A2(new_n363), .A3(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n371), .B1(new_n367), .B2(new_n368), .ZN(new_n372));
  OAI21_X1  g171(.A(KEYINPUT34), .B1(new_n337), .B2(new_n340), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n365), .A2(new_n364), .A3(new_n366), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n373), .A2(new_n374), .A3(KEYINPUT77), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n372), .A2(new_n375), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n376), .B1(new_n355), .B2(new_n363), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT36), .B1(new_n370), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n369), .ZN(new_n379));
  NOR3_X1   g178(.A1(new_n360), .A2(new_n361), .A3(new_n362), .ZN(new_n380));
  AOI221_X4 g179(.A(new_n356), .B1(KEYINPUT33), .B2(new_n354), .C1(new_n359), .C2(new_n344), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n379), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT36), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n355), .A2(new_n363), .A3(new_n369), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  AND2_X1   g184(.A1(new_n378), .A2(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT88), .ZN(new_n387));
  NAND2_X1  g186(.A1(G226gat), .A2(G233gat), .ZN(new_n388));
  INV_X1    g187(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(KEYINPUT29), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n319), .A2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT78), .ZN(new_n392));
  XNOR2_X1  g191(.A(G197gat), .B(G204gat), .ZN(new_n393));
  INV_X1    g192(.A(G211gat), .ZN(new_n394));
  INV_X1    g193(.A(G218gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n393), .B1(KEYINPUT22), .B2(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(G211gat), .B(G218gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n397), .B(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n318), .A2(new_n389), .A3(new_n285), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n391), .A2(new_n392), .A3(new_n399), .A4(new_n400), .ZN(new_n401));
  INV_X1    g200(.A(new_n390), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n399), .B(new_n400), .C1(new_n335), .C2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n406));
  INV_X1    g205(.A(new_n285), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n303), .B2(new_n317), .ZN(new_n408));
  OAI211_X1 g207(.A(new_n406), .B(new_n388), .C1(new_n408), .C2(KEYINPUT29), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT29), .B1(new_n318), .B2(new_n285), .ZN(new_n410));
  OAI21_X1  g209(.A(KEYINPUT79), .B1(new_n410), .B2(new_n389), .ZN(new_n411));
  INV_X1    g210(.A(new_n398), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n397), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n319), .A2(new_n389), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n409), .A2(new_n411), .A3(new_n413), .A4(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n405), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT80), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT80), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n405), .A2(new_n418), .A3(new_n415), .ZN(new_n419));
  XOR2_X1   g218(.A(G64gat), .B(G92gat), .Z(new_n420));
  XNOR2_X1  g219(.A(G8gat), .B(G36gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n420), .B(new_n421), .ZN(new_n422));
  XNOR2_X1  g221(.A(new_n422), .B(KEYINPUT81), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n417), .A2(new_n419), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g223(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n425));
  NOR2_X1   g224(.A1(new_n403), .A2(KEYINPUT78), .ZN(new_n426));
  OAI211_X1 g225(.A(new_n415), .B(new_n422), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n427), .A2(KEYINPUT30), .ZN(new_n428));
  INV_X1    g227(.A(KEYINPUT30), .ZN(new_n429));
  NAND4_X1  g228(.A1(new_n405), .A2(new_n429), .A3(new_n415), .A4(new_n422), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n428), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n424), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n326), .A2(new_n328), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n433), .A2(KEYINPUT72), .ZN(new_n434));
  INV_X1    g233(.A(G155gat), .ZN(new_n435));
  INV_X1    g234(.A(G162gat), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(G155gat), .A2(G162gat), .ZN(new_n438));
  AND2_X1   g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n440));
  XNOR2_X1  g239(.A(G141gat), .B(G148gat), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n439), .B(new_n440), .C1(KEYINPUT2), .C2(new_n441), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n439), .B1(KEYINPUT2), .B2(new_n441), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n438), .B1(new_n437), .B2(KEYINPUT2), .ZN(new_n444));
  INV_X1    g243(.A(G141gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G148gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n446), .A2(KEYINPUT83), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT83), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n448), .A2(new_n445), .A3(G148gat), .ZN(new_n449));
  INV_X1    g248(.A(G148gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(G141gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n447), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g251(.A1(new_n443), .A2(KEYINPUT82), .B1(new_n444), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n326), .A2(new_n328), .A3(new_n329), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n442), .A3(new_n453), .A4(new_n454), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT4), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n452), .A2(new_n444), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT2), .B1(new_n451), .B2(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n437), .A2(new_n438), .ZN(new_n460));
  OAI21_X1  g259(.A(KEYINPUT82), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n442), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT3), .ZN(new_n464));
  NAND4_X1  g263(.A1(new_n442), .A2(new_n458), .A3(new_n461), .A4(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n465), .A3(new_n433), .ZN(new_n466));
  INV_X1    g265(.A(new_n462), .ZN(new_n467));
  AND2_X1   g266(.A1(new_n324), .A2(new_n322), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT71), .B(G113gat), .Z(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(G120gat), .ZN(new_n470));
  AOI22_X1  g269(.A1(new_n468), .A2(new_n470), .B1(new_n323), .B2(new_n325), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n467), .A2(KEYINPUT4), .A3(new_n471), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n457), .A2(new_n466), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(G225gat), .A2(G233gat), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n453), .A2(new_n471), .A3(new_n442), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n433), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n479), .A2(new_n475), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT39), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n476), .A2(new_n482), .ZN(new_n483));
  XOR2_X1   g282(.A(G1gat), .B(G29gat), .Z(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT0), .ZN(new_n485));
  XNOR2_X1  g284(.A(G57gat), .B(G85gat), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n485), .B(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(new_n487), .B(KEYINPUT87), .Z(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n473), .A2(new_n481), .A3(new_n475), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n483), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT40), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT5), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n494), .B1(new_n479), .B2(new_n475), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n462), .A2(KEYINPUT4), .A3(new_n433), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n455), .B2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n466), .A2(new_n474), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n495), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n471), .B1(new_n462), .B2(KEYINPUT3), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n475), .B1(new_n500), .B2(new_n465), .ZN(new_n501));
  NAND4_X1  g300(.A1(new_n501), .A2(new_n457), .A3(new_n494), .A4(new_n472), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n499), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(new_n488), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n483), .A2(new_n489), .A3(KEYINPUT40), .A4(new_n490), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n493), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n432), .A2(new_n506), .ZN(new_n507));
  INV_X1    g306(.A(G228gat), .ZN(new_n508));
  NOR2_X1   g307(.A1(new_n508), .A2(new_n339), .ZN(new_n509));
  INV_X1    g308(.A(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  XNOR2_X1  g311(.A(G78gat), .B(G106gat), .ZN(new_n513));
  XNOR2_X1  g312(.A(new_n512), .B(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT3), .B1(new_n413), .B2(new_n516), .ZN(new_n517));
  OAI22_X1  g316(.A1(new_n517), .A2(new_n467), .B1(KEYINPUT85), .B2(new_n509), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n413), .B1(new_n516), .B2(new_n465), .ZN(new_n519));
  OAI21_X1  g318(.A(G22gat), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g319(.A(new_n464), .B1(new_n399), .B2(KEYINPUT29), .ZN(new_n521));
  AOI22_X1  g320(.A1(new_n521), .A2(new_n462), .B1(new_n511), .B2(new_n510), .ZN(new_n522));
  INV_X1    g321(.A(G22gat), .ZN(new_n523));
  INV_X1    g322(.A(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G50gat), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n520), .A2(new_n525), .A3(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n527), .B1(new_n520), .B2(new_n525), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n515), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n518), .A2(new_n519), .A3(G22gat), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n523), .B1(new_n522), .B2(new_n524), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n526), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n520), .A2(new_n525), .A3(new_n527), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n533), .A2(new_n514), .A3(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n530), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n507), .A2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT37), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n405), .A2(new_n539), .A3(new_n415), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT38), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n423), .A2(new_n541), .ZN(new_n542));
  AOI22_X1  g341(.A1(new_n319), .A2(new_n390), .B1(new_n408), .B2(new_n389), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n539), .B1(new_n543), .B2(new_n413), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n409), .A2(new_n411), .A3(new_n399), .A4(new_n414), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n542), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n540), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT6), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n499), .A2(new_n487), .A3(new_n502), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n504), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n487), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n503), .A2(KEYINPUT6), .A3(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n547), .A2(new_n550), .A3(new_n552), .A4(new_n427), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n417), .A2(KEYINPUT37), .A3(new_n419), .ZN(new_n554));
  INV_X1    g353(.A(new_n422), .ZN(new_n555));
  NAND3_X1  g354(.A1(new_n554), .A2(new_n555), .A3(new_n540), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n553), .B1(new_n556), .B2(KEYINPUT38), .ZN(new_n557));
  OAI21_X1  g356(.A(new_n387), .B1(new_n538), .B2(new_n557), .ZN(new_n558));
  AND3_X1   g357(.A1(new_n405), .A2(new_n418), .A3(new_n415), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n418), .B1(new_n405), .B2(new_n415), .ZN(new_n560));
  NOR3_X1   g359(.A1(new_n559), .A2(new_n560), .A3(new_n539), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n540), .A2(new_n555), .ZN(new_n562));
  OAI21_X1  g361(.A(KEYINPUT38), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n553), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n536), .B1(new_n432), .B2(new_n506), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(KEYINPUT88), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n549), .A2(KEYINPUT84), .A3(new_n548), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n503), .A2(new_n551), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT84), .B1(new_n549), .B2(new_n548), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n552), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(new_n424), .A3(new_n431), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT86), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n536), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n530), .A2(KEYINPUT86), .A3(new_n535), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n573), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n386), .A2(new_n558), .A3(new_n567), .A4(new_n578), .ZN(new_n579));
  OAI211_X1 g378(.A(new_n372), .B(new_n375), .C1(new_n380), .C2(new_n381), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n580), .A2(new_n537), .A3(new_n384), .ZN(new_n581));
  OAI21_X1  g380(.A(KEYINPUT35), .B1(new_n581), .B2(new_n573), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n369), .B1(new_n355), .B2(new_n363), .ZN(new_n583));
  NOR2_X1   g382(.A1(new_n370), .A2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n432), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n550), .A2(new_n552), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n536), .A2(KEYINPUT35), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .A4(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n256), .B1(new_n579), .B2(new_n589), .ZN(new_n590));
  OR2_X1    g389(.A1(G57gat), .A2(G64gat), .ZN(new_n591));
  NAND2_X1  g390(.A1(G57gat), .A2(G64gat), .ZN(new_n592));
  AND2_X1   g391(.A1(G71gat), .A2(G78gat), .ZN(new_n593));
  OAI211_X1 g392(.A(new_n591), .B(new_n592), .C1(new_n593), .C2(KEYINPUT9), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(KEYINPUT94), .B2(new_n593), .ZN(new_n595));
  XNOR2_X1  g394(.A(G71gat), .B(G78gat), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n595), .B(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT21), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(G231gat), .A2(G233gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n601), .B(G127gat), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n597), .A2(KEYINPUT95), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(KEYINPUT21), .A3(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n218), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n602), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(new_n435), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n607), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  INV_X1    g412(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(G85gat), .A2(G92gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(KEYINPUT7), .ZN(new_n616));
  NAND2_X1  g415(.A1(G99gat), .A2(G106gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT8), .ZN(new_n618));
  OAI211_X1 g417(.A(new_n616), .B(new_n618), .C1(G85gat), .C2(G92gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G99gat), .B(G106gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n622), .B1(new_n238), .B2(new_n240), .ZN(new_n623));
  AND2_X1   g422(.A1(G232gat), .A2(G233gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(new_n231), .A2(new_n621), .B1(KEYINPUT41), .B2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n614), .B1(new_n623), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT96), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n623), .A2(new_n614), .A3(new_n625), .ZN(new_n630));
  NOR2_X1   g429(.A1(new_n624), .A2(KEYINPUT41), .ZN(new_n631));
  XNOR2_X1  g430(.A(G134gat), .B(G162gat), .ZN(new_n632));
  XOR2_X1   g431(.A(new_n631), .B(new_n632), .Z(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n630), .B(new_n634), .C1(new_n626), .C2(new_n627), .ZN(new_n635));
  OAI21_X1  g434(.A(KEYINPUT97), .B1(new_n629), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n623), .A2(new_n625), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(new_n613), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(KEYINPUT96), .ZN(new_n639));
  AND2_X1   g438(.A1(new_n630), .A2(new_n634), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n639), .A2(new_n640), .A3(new_n641), .A4(new_n628), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n634), .B1(new_n638), .B2(new_n630), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n643), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT98), .B1(new_n612), .B2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(new_n611), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n607), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT98), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n644), .B1(new_n636), .B2(new_n642), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n649), .A2(new_n650), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(G230gat), .A2(G233gat), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(new_n620), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n597), .B1(KEYINPUT99), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(new_n621), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n620), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n622), .B1(new_n597), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT10), .ZN(new_n662));
  NAND3_X1  g461(.A1(new_n658), .A2(new_n661), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n604), .A4(new_n621), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n655), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n654), .B1(new_n658), .B2(new_n661), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT100), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(KEYINPUT100), .B(new_n670), .C1(new_n665), .C2(new_n666), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n653), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n590), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n676), .A2(new_n572), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT101), .B(G1gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(G1324gat));
  INV_X1    g478(.A(new_n676), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n217), .B1(new_n680), .B2(new_n432), .ZN(new_n681));
  XNOR2_X1  g480(.A(KEYINPUT16), .B(G8gat), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n676), .A2(new_n585), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g482(.A(KEYINPUT42), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(KEYINPUT42), .B2(new_n683), .ZN(G1325gat));
  AOI21_X1  g484(.A(G15gat), .B1(new_n680), .B2(new_n584), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT102), .ZN(new_n687));
  INV_X1    g486(.A(new_n386), .ZN(new_n688));
  AND2_X1   g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n687), .B1(new_n680), .B2(new_n689), .ZN(G1326gat));
  NAND2_X1  g489(.A1(new_n680), .A2(new_n577), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT103), .ZN(new_n692));
  XNOR2_X1  g491(.A(KEYINPUT43), .B(G22gat), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n692), .B(new_n693), .ZN(G1327gat));
  INV_X1    g493(.A(KEYINPUT106), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n651), .A2(new_n695), .ZN(new_n696));
  AOI211_X1 g495(.A(KEYINPUT106), .B(new_n644), .C1(new_n636), .C2(new_n642), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g497(.A1(new_n698), .A2(KEYINPUT44), .ZN(new_n699));
  AND3_X1   g498(.A1(new_n565), .A2(KEYINPUT88), .A3(new_n566), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n378), .A2(new_n578), .A3(new_n385), .ZN(new_n701));
  AOI21_X1  g500(.A(KEYINPUT88), .B1(new_n565), .B2(new_n566), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n582), .A2(new_n588), .ZN(new_n704));
  OAI211_X1 g503(.A(KEYINPUT107), .B(new_n699), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT44), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n651), .B1(new_n579), .B2(new_n589), .ZN(new_n707));
  OAI21_X1  g506(.A(new_n705), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n579), .A2(new_n589), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT107), .B1(new_n709), .B2(new_n699), .ZN(new_n710));
  OR2_X1    g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n612), .A2(KEYINPUT104), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT104), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n649), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NOR3_X1   g514(.A1(new_n715), .A2(new_n256), .A3(new_n674), .ZN(new_n716));
  XNOR2_X1  g515(.A(new_n716), .B(KEYINPUT105), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n711), .A2(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n572), .ZN(new_n719));
  AOI21_X1  g518(.A(new_n223), .B1(new_n718), .B2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n649), .A2(new_n651), .A3(new_n674), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n590), .A2(new_n721), .ZN(new_n722));
  INV_X1    g521(.A(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n723), .A2(new_n223), .A3(new_n719), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT45), .ZN(new_n725));
  INV_X1    g524(.A(new_n725), .ZN(new_n726));
  OR3_X1    g525(.A1(new_n720), .A2(new_n726), .A3(KEYINPUT108), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT108), .B1(new_n720), .B2(new_n726), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(G1328gat));
  INV_X1    g528(.A(KEYINPUT109), .ZN(new_n730));
  AOI21_X1  g529(.A(G36gat), .B1(new_n730), .B2(KEYINPUT46), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n723), .A2(new_n432), .A3(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n730), .A2(KEYINPUT46), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n732), .B(new_n733), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n718), .A2(new_n432), .ZN(new_n735));
  OAI21_X1  g534(.A(new_n734), .B1(new_n735), .B2(new_n220), .ZN(G1329gat));
  INV_X1    g535(.A(G43gat), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n718), .B2(new_n688), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT47), .ZN(new_n739));
  INV_X1    g538(.A(new_n584), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n722), .A2(G43gat), .A3(new_n740), .ZN(new_n741));
  OR3_X1    g540(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n739), .B1(new_n738), .B2(new_n741), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1330gat));
  NAND2_X1  g543(.A1(new_n718), .A2(new_n536), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(G50gat), .ZN(new_n746));
  INV_X1    g545(.A(new_n577), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n722), .A2(G50gat), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n746), .A2(KEYINPUT48), .A3(new_n749), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n577), .B(new_n717), .C1(new_n708), .C2(new_n710), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(G50gat), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT110), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n748), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n751), .A2(KEYINPUT110), .A3(G50gat), .ZN(new_n755));
  AOI211_X1 g554(.A(KEYINPUT111), .B(KEYINPUT48), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT111), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n752), .A2(new_n753), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n755), .A3(new_n749), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n757), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n750), .B1(new_n756), .B2(new_n761), .ZN(G1331gat));
  NAND2_X1  g561(.A1(new_n252), .A2(new_n255), .ZN(new_n763));
  INV_X1    g562(.A(new_n674), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n653), .A2(new_n763), .A3(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n709), .A2(new_n765), .ZN(new_n766));
  INV_X1    g565(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(new_n719), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g568(.A1(new_n766), .A2(new_n585), .ZN(new_n770));
  NOR2_X1   g569(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n771));
  AND2_X1   g570(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n770), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n770), .B2(new_n771), .ZN(G1333gat));
  NOR3_X1   g573(.A1(new_n766), .A2(G71gat), .A3(new_n740), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n767), .A2(new_n688), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n775), .B1(G71gat), .B2(new_n776), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g577(.A1(new_n767), .A2(new_n577), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n779), .B(G78gat), .ZN(G1335gat));
  NAND3_X1  g579(.A1(new_n707), .A2(new_n256), .A3(new_n612), .ZN(new_n781));
  OR2_X1    g580(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(KEYINPUT51), .ZN(new_n783));
  AND3_X1   g582(.A1(new_n782), .A2(new_n674), .A3(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(G85gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n784), .A2(new_n785), .A3(new_n719), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n763), .A2(new_n649), .A3(new_n764), .ZN(new_n787));
  AND2_X1   g586(.A1(new_n711), .A2(new_n787), .ZN(new_n788));
  AND2_X1   g587(.A1(new_n788), .A2(new_n719), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n786), .B1(new_n789), .B2(new_n785), .ZN(G1336gat));
  NOR2_X1   g589(.A1(new_n585), .A2(G92gat), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n432), .B(new_n787), .C1(new_n708), .C2(new_n710), .ZN(new_n792));
  AOI22_X1  g591(.A1(new_n784), .A2(new_n791), .B1(G92gat), .B2(new_n792), .ZN(new_n793));
  AOI21_X1  g592(.A(KEYINPUT112), .B1(new_n792), .B2(G92gat), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n794), .A2(KEYINPUT52), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n793), .B(new_n795), .ZN(G1337gat));
  INV_X1    g595(.A(G99gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n784), .A2(new_n797), .A3(new_n584), .ZN(new_n798));
  AND2_X1   g597(.A1(new_n788), .A2(new_n688), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n799), .B2(new_n797), .ZN(G1338gat));
  INV_X1    g599(.A(G106gat), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n788), .B2(new_n577), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n537), .A2(G106gat), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n802), .B1(new_n784), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT53), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n801), .B1(new_n788), .B2(new_n536), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n784), .A2(new_n803), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n805), .ZN(new_n808));
  OAI22_X1  g607(.A1(new_n804), .A2(new_n805), .B1(new_n806), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n663), .A2(new_n664), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n654), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n663), .A2(new_n655), .A3(new_n664), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n811), .A2(KEYINPUT54), .A3(new_n812), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT54), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n670), .B1(new_n665), .B2(new_n814), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT55), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  OR3_X1    g617(.A1(new_n665), .A2(new_n666), .A3(new_n671), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n813), .A2(KEYINPUT55), .A3(new_n815), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n821), .B1(new_n252), .B2(new_n255), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n235), .B1(new_n247), .B2(new_n233), .ZN(new_n824));
  INV_X1    g623(.A(new_n236), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n230), .A2(new_n233), .A3(new_n825), .ZN(new_n826));
  INV_X1    g625(.A(KEYINPUT113), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n827), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n823), .B(new_n206), .C1(new_n824), .C2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(new_n828), .B(new_n829), .C1(new_n243), .C2(new_n235), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(new_n206), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT114), .ZN(new_n834));
  AND4_X1   g633(.A1(new_n255), .A2(new_n674), .A3(new_n831), .A4(new_n834), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT115), .B1(new_n822), .B2(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT115), .ZN(new_n837));
  INV_X1    g636(.A(new_n831), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n823), .B1(new_n832), .B2(new_n206), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n840), .A2(new_n255), .A3(new_n674), .ZN(new_n841));
  OAI211_X1 g640(.A(new_n837), .B(new_n841), .C1(new_n256), .C2(new_n821), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n836), .A2(new_n842), .A3(new_n698), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n820), .A2(new_n819), .ZN(new_n844));
  AOI21_X1  g643(.A(KEYINPUT55), .B1(new_n813), .B2(new_n815), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n840), .A3(new_n255), .ZN(new_n847));
  NOR3_X1   g646(.A1(new_n847), .A2(new_n696), .A3(new_n697), .ZN(new_n848));
  INV_X1    g647(.A(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n715), .B1(new_n843), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n647), .A2(new_n652), .A3(new_n256), .A4(new_n764), .ZN(new_n851));
  INV_X1    g650(.A(new_n851), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n850), .A2(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n432), .A2(new_n572), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n853), .A2(new_n855), .ZN(new_n856));
  INV_X1    g655(.A(new_n581), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  INV_X1    g657(.A(new_n858), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n327), .A3(new_n763), .ZN(new_n860));
  NOR2_X1   g659(.A1(new_n740), .A2(new_n577), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT116), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g663(.A(KEYINPUT116), .B1(new_n856), .B2(new_n861), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n864), .A2(new_n256), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n860), .B1(new_n866), .B2(new_n320), .ZN(G1340gat));
  AOI21_X1  g666(.A(G120gat), .B1(new_n859), .B2(new_n674), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n864), .A2(new_n865), .ZN(new_n869));
  NOR2_X1   g668(.A1(new_n764), .A2(new_n321), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(G1341gat));
  NOR3_X1   g670(.A1(new_n858), .A2(KEYINPUT117), .A3(new_n612), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(G127gat), .ZN(new_n873));
  OAI21_X1  g672(.A(KEYINPUT117), .B1(new_n858), .B2(new_n612), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n715), .A2(G127gat), .ZN(new_n875));
  AOI22_X1  g674(.A1(new_n873), .A2(new_n874), .B1(new_n869), .B2(new_n875), .ZN(G1342gat));
  NAND2_X1  g675(.A1(new_n869), .A2(new_n646), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n877), .A2(G134gat), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n853), .A2(new_n572), .ZN(new_n880));
  NOR4_X1   g679(.A1(new_n581), .A2(new_n651), .A3(G134gat), .A4(new_n432), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(KEYINPUT118), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n882), .A2(KEYINPUT118), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n879), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OR3_X1    g684(.A1(new_n883), .A2(new_n884), .A3(new_n879), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n878), .A2(new_n885), .A3(new_n886), .ZN(G1343gat));
  NOR2_X1   g686(.A1(new_n688), .A2(new_n855), .ZN(new_n888));
  INV_X1    g687(.A(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT57), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n747), .A2(new_n890), .ZN(new_n891));
  INV_X1    g690(.A(new_n891), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n818), .A2(KEYINPUT119), .A3(new_n819), .A4(new_n820), .ZN(new_n893));
  INV_X1    g692(.A(KEYINPUT119), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n844), .B2(new_n845), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n763), .A2(new_n893), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n646), .B1(new_n896), .B2(new_n841), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n612), .B1(new_n897), .B2(new_n848), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n852), .B1(new_n898), .B2(KEYINPUT120), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT120), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n900), .B(new_n612), .C1(new_n897), .C2(new_n848), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n892), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  OAI21_X1  g701(.A(new_n536), .B1(new_n850), .B2(new_n852), .ZN(new_n903));
  AOI22_X1  g702(.A1(new_n902), .A2(KEYINPUT121), .B1(new_n903), .B2(new_n890), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n899), .A2(new_n901), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n891), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT121), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n889), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n445), .B1(new_n909), .B2(new_n763), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n688), .A2(new_n537), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT122), .Z(new_n912));
  NAND2_X1  g711(.A1(new_n856), .A2(new_n912), .ZN(new_n913));
  NOR3_X1   g712(.A1(new_n913), .A2(G141gat), .A3(new_n256), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT58), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n904), .A2(new_n908), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n916), .A2(new_n763), .A3(new_n888), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G141gat), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT58), .ZN(new_n919));
  INV_X1    g718(.A(new_n914), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n915), .A2(new_n921), .ZN(G1344gat));
  INV_X1    g721(.A(new_n913), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n923), .A2(new_n450), .A3(new_n674), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT59), .B(new_n450), .C1(new_n909), .C2(new_n674), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT59), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n852), .A2(KEYINPUT123), .ZN(new_n927));
  NOR2_X1   g726(.A1(new_n847), .A2(new_n651), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n612), .B1(new_n897), .B2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT123), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n851), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n747), .A2(KEYINPUT57), .ZN(new_n933));
  AOI22_X1  g732(.A1(new_n903), .A2(KEYINPUT57), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n934), .A2(new_n674), .A3(new_n888), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n926), .B1(new_n935), .B2(G148gat), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n924), .B1(new_n925), .B2(new_n936), .ZN(G1345gat));
  INV_X1    g736(.A(new_n909), .ZN(new_n938));
  INV_X1    g737(.A(new_n715), .ZN(new_n939));
  OAI21_X1  g738(.A(G155gat), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n923), .A2(new_n435), .A3(new_n649), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1346gat));
  OAI21_X1  g741(.A(G162gat), .B1(new_n938), .B2(new_n698), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n651), .A2(G162gat), .A3(new_n432), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n880), .A2(new_n912), .A3(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n943), .A2(new_n945), .ZN(G1347gat));
  NOR2_X1   g745(.A1(new_n585), .A2(new_n719), .ZN(new_n947));
  INV_X1    g746(.A(new_n947), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n853), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n857), .ZN(new_n950));
  INV_X1    g749(.A(new_n950), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n951), .A2(new_n257), .A3(new_n763), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(new_n861), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n954), .A2(new_n763), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n955), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n956));
  INV_X1    g755(.A(new_n956), .ZN(new_n957));
  AOI21_X1  g756(.A(KEYINPUT124), .B1(new_n955), .B2(G169gat), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n952), .B1(new_n957), .B2(new_n958), .ZN(G1348gat));
  AOI21_X1  g758(.A(G176gat), .B1(new_n951), .B2(new_n674), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n764), .B1(new_n298), .B2(new_n299), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n960), .B1(new_n954), .B2(new_n961), .ZN(G1349gat));
  OAI21_X1  g761(.A(G183gat), .B1(new_n953), .B2(new_n939), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n649), .A2(new_n281), .ZN(new_n964));
  OAI21_X1  g763(.A(new_n963), .B1(new_n950), .B2(new_n964), .ZN(new_n965));
  XNOR2_X1  g764(.A(new_n965), .B(KEYINPUT60), .ZN(G1350gat));
  NOR2_X1   g765(.A1(new_n696), .A2(new_n697), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n951), .A2(new_n277), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n954), .A2(new_n646), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n970));
  NAND3_X1  g769(.A1(new_n969), .A2(new_n970), .A3(G190gat), .ZN(new_n971));
  INV_X1    g770(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n970), .B1(new_n969), .B2(G190gat), .ZN(new_n973));
  OAI21_X1  g772(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(G1351gat));
  OR2_X1    g773(.A1(new_n850), .A2(new_n852), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n975), .A2(new_n911), .A3(new_n947), .ZN(new_n976));
  NOR2_X1   g775(.A1(new_n256), .A2(G197gat), .ZN(new_n977));
  INV_X1    g776(.A(new_n977), .ZN(new_n978));
  OR3_X1    g777(.A1(new_n976), .A2(KEYINPUT125), .A3(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(KEYINPUT125), .B1(new_n976), .B2(new_n978), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n688), .A2(new_n948), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n934), .A2(new_n763), .A3(new_n982), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G197gat), .ZN(new_n984));
  NAND2_X1  g783(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n985), .A2(KEYINPUT126), .ZN(new_n986));
  INV_X1    g785(.A(KEYINPUT126), .ZN(new_n987));
  NAND3_X1  g786(.A1(new_n981), .A2(new_n987), .A3(new_n984), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n986), .A2(new_n988), .ZN(G1352gat));
  NOR3_X1   g788(.A1(new_n976), .A2(G204gat), .A3(new_n764), .ZN(new_n990));
  XNOR2_X1  g789(.A(new_n990), .B(KEYINPUT62), .ZN(new_n991));
  INV_X1    g790(.A(G204gat), .ZN(new_n992));
  INV_X1    g791(.A(new_n934), .ZN(new_n993));
  INV_X1    g792(.A(new_n982), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n993), .A2(new_n764), .A3(new_n994), .ZN(new_n995));
  OAI21_X1  g794(.A(new_n991), .B1(new_n992), .B2(new_n995), .ZN(G1353gat));
  INV_X1    g795(.A(new_n976), .ZN(new_n997));
  NAND3_X1  g796(.A1(new_n997), .A2(new_n394), .A3(new_n649), .ZN(new_n998));
  NAND4_X1  g797(.A1(new_n934), .A2(KEYINPUT127), .A3(new_n649), .A4(new_n982), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n999), .A2(G211gat), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n903), .A2(KEYINPUT57), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n932), .A2(new_n933), .ZN(new_n1002));
  NAND4_X1  g801(.A1(new_n1001), .A2(new_n649), .A3(new_n1002), .A4(new_n982), .ZN(new_n1003));
  INV_X1    g802(.A(KEYINPUT127), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  AND4_X1   g805(.A1(KEYINPUT63), .A2(new_n1005), .A3(G211gat), .A4(new_n999), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  NAND3_X1  g807(.A1(new_n997), .A2(new_n395), .A3(new_n967), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n993), .A2(new_n651), .A3(new_n994), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1009), .B1(new_n1010), .B2(new_n395), .ZN(G1355gat));
endmodule


