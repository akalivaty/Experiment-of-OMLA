//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 1 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:42 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT64), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G134), .ZN(new_n193));
  INV_X1    g007(.A(G137), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(KEYINPUT11), .ZN(new_n195));
  AND3_X1   g009(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(KEYINPUT11), .A3(G134), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT11), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G137), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  OAI21_X1  g014(.A(G131), .B1(new_n196), .B2(new_n200), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n193), .A3(new_n195), .ZN(new_n202));
  INV_X1    g016(.A(G131), .ZN(new_n203));
  NAND4_X1  g017(.A1(new_n202), .A2(new_n203), .A3(new_n197), .A4(new_n199), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n201), .A2(new_n204), .ZN(new_n205));
  XNOR2_X1  g019(.A(new_n205), .B(KEYINPUT80), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  OAI211_X1 g022(.A(new_n207), .B(G146), .C1(new_n208), .C2(KEYINPUT1), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n208), .A2(new_n210), .A3(G143), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT79), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n208), .A2(KEYINPUT1), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n207), .A2(G146), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(KEYINPUT65), .ZN(new_n219));
  XNOR2_X1  g033(.A(G143), .B(G146), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(new_n215), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT79), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n212), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n214), .A2(new_n223), .A3(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G107), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G104), .ZN(new_n228));
  INV_X1    g042(.A(G104), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(G107), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n228), .A2(new_n230), .A3(KEYINPUT78), .ZN(new_n231));
  OAI211_X1 g045(.A(new_n231), .B(G101), .C1(KEYINPUT78), .C2(new_n228), .ZN(new_n232));
  OAI21_X1  g046(.A(KEYINPUT3), .B1(new_n229), .B2(G107), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(new_n227), .A3(G104), .ZN(new_n235));
  INV_X1    g049(.A(G101), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n233), .A2(new_n235), .A3(new_n236), .A4(new_n230), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n226), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n216), .A2(new_n217), .A3(KEYINPUT0), .A4(G128), .ZN(new_n242));
  XNOR2_X1  g056(.A(KEYINPUT0), .B(G128), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n242), .B1(new_n220), .B2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n233), .A2(new_n235), .A3(new_n230), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT4), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n246), .A2(new_n247), .A3(G101), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n246), .A2(G101), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n237), .A2(KEYINPUT4), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n245), .B(new_n248), .C1(new_n249), .C2(new_n250), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n221), .B1(new_n220), .B2(new_n215), .ZN(new_n252));
  AND4_X1   g066(.A1(new_n221), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n213), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n238), .A2(KEYINPUT10), .A3(new_n254), .ZN(new_n255));
  NAND4_X1  g069(.A1(new_n206), .A2(new_n241), .A3(new_n251), .A4(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n205), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n232), .A2(new_n237), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n212), .B1(new_n219), .B2(new_n222), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n257), .B1(new_n239), .B2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT12), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT12), .ZN(new_n263));
  AOI211_X1 g077(.A(new_n263), .B(new_n257), .C1(new_n239), .C2(new_n260), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n256), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G227), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n267), .B(KEYINPUT77), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(new_n212), .B(KEYINPUT79), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n258), .B1(new_n271), .B2(new_n223), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n255), .B(new_n251), .C1(new_n272), .C2(KEYINPUT10), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n270), .B1(new_n274), .B2(new_n206), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n205), .ZN(new_n276));
  AOI22_X1  g090(.A1(new_n265), .A2(new_n270), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(G469), .B1(new_n277), .B2(G902), .ZN(new_n278));
  INV_X1    g092(.A(new_n260), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n205), .B1(new_n279), .B2(new_n272), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n263), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n261), .A2(KEYINPUT12), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n275), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n276), .A2(new_n256), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n270), .ZN(new_n286));
  AOI21_X1  g100(.A(G902), .B1(new_n284), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(KEYINPUT81), .B(G469), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n189), .B1(new_n278), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G952), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n291), .A2(KEYINPUT98), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(KEYINPUT98), .ZN(new_n293));
  AOI21_X1  g107(.A(G953), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(G234), .A2(G237), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XOR2_X1   g110(.A(new_n296), .B(KEYINPUT99), .Z(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  XNOR2_X1  g112(.A(KEYINPUT21), .B(G898), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n295), .A2(G902), .A3(G953), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n298), .B1(new_n299), .B2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(G478), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n304), .A2(KEYINPUT15), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  INV_X1    g120(.A(G122), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(G116), .ZN(new_n308));
  INV_X1    g122(.A(G116), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G122), .ZN(new_n310));
  AOI21_X1  g124(.A(KEYINPUT92), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n308), .A2(new_n310), .A3(KEYINPUT92), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(G107), .ZN(new_n314));
  INV_X1    g128(.A(new_n313), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n227), .B1(new_n315), .B2(new_n311), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n191), .A2(new_n193), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n208), .A2(G143), .ZN(new_n319));
  NOR2_X1   g133(.A1(new_n207), .A2(G128), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT95), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n207), .A2(G128), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n208), .A2(G143), .ZN(new_n323));
  INV_X1    g137(.A(KEYINPUT95), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  AOI22_X1  g140(.A1(new_n314), .A2(new_n316), .B1(new_n318), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n319), .B1(KEYINPUT13), .B2(new_n323), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT93), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n190), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT13), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n322), .B1(new_n320), .B2(new_n331), .ZN(new_n332));
  OAI211_X1 g146(.A(new_n332), .B(KEYINPUT93), .C1(new_n331), .C2(new_n322), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT94), .ZN(new_n334));
  AND3_X1   g148(.A1(new_n330), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n334), .B1(new_n330), .B2(new_n333), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n327), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n309), .A2(KEYINPUT14), .A3(G122), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n308), .A2(new_n310), .ZN(new_n339));
  OAI211_X1 g153(.A(G107), .B(new_n338), .C1(new_n339), .C2(KEYINPUT14), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT96), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n326), .A2(new_n318), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n321), .A2(new_n317), .A3(new_n325), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n316), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(new_n187), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G217), .A3(new_n266), .ZN(new_n348));
  INV_X1    g162(.A(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n337), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n337), .B2(new_n346), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n306), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT97), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT97), .ZN(new_n354));
  OAI211_X1 g168(.A(new_n354), .B(new_n306), .C1(new_n350), .C2(new_n351), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n305), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n355), .A2(new_n305), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(G237), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n359), .A2(new_n266), .A3(G214), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n207), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n359), .A2(new_n266), .A3(G143), .A4(G214), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(KEYINPUT18), .ZN(new_n364));
  OAI21_X1  g178(.A(new_n363), .B1(new_n364), .B2(new_n203), .ZN(new_n365));
  NAND4_X1  g179(.A1(new_n361), .A2(KEYINPUT18), .A3(G131), .A4(new_n362), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(G140), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(G125), .ZN(new_n369));
  INV_X1    g183(.A(G125), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(G140), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G146), .ZN(new_n373));
  XNOR2_X1  g187(.A(G125), .B(G140), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(new_n210), .ZN(new_n375));
  INV_X1    g189(.A(KEYINPUT86), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n373), .B2(new_n375), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n367), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n368), .A3(G125), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n381), .B1(new_n372), .B2(new_n380), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(new_n210), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n374), .A2(KEYINPUT16), .ZN(new_n384));
  AOI21_X1  g198(.A(G146), .B1(new_n384), .B2(new_n381), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT90), .B1(new_n383), .B2(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n203), .B1(new_n361), .B2(new_n362), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n382), .A2(new_n210), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n384), .A2(G146), .A3(new_n381), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n386), .A2(new_n388), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n363), .A2(G131), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n361), .A2(new_n203), .A3(new_n362), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n397), .A2(KEYINPUT91), .B1(KEYINPUT17), .B2(new_n387), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n379), .B1(new_n393), .B2(new_n398), .ZN(new_n399));
  XOR2_X1   g213(.A(G113), .B(G122), .Z(new_n400));
  XOR2_X1   g214(.A(KEYINPUT87), .B(G104), .Z(new_n401));
  XNOR2_X1  g215(.A(new_n400), .B(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT89), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n402), .B(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n405), .B(new_n379), .C1(new_n393), .C2(new_n398), .ZN(new_n406));
  AOI21_X1  g220(.A(G902), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(G475), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT88), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n394), .A2(new_n396), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n374), .A2(KEYINPUT19), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n374), .A2(KEYINPUT19), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n210), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n411), .A2(new_n391), .A3(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n379), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n410), .B1(new_n416), .B2(new_n402), .ZN(new_n417));
  INV_X1    g231(.A(new_n402), .ZN(new_n418));
  AOI211_X1 g232(.A(KEYINPUT88), .B(new_n418), .C1(new_n379), .C2(new_n415), .ZN(new_n419));
  OAI21_X1  g233(.A(new_n406), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(G475), .A2(G902), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT20), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n420), .A2(new_n424), .A3(new_n421), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n409), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n290), .A2(new_n303), .A3(new_n358), .A4(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT85), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n245), .A2(G125), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT82), .B(G224), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n266), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT7), .ZN(new_n432));
  OAI211_X1 g246(.A(new_n429), .B(new_n432), .C1(G125), .C2(new_n259), .ZN(new_n433));
  OAI21_X1  g247(.A(new_n429), .B1(G125), .B2(new_n259), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n434), .A2(KEYINPUT7), .A3(new_n431), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT5), .ZN(new_n436));
  INV_X1    g250(.A(G119), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n436), .A2(new_n437), .A3(G116), .ZN(new_n438));
  XOR2_X1   g252(.A(G116), .B(G119), .Z(new_n439));
  OAI211_X1 g253(.A(G113), .B(new_n438), .C1(new_n439), .C2(new_n436), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT2), .B(G113), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(G116), .B(G119), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n440), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n258), .ZN(new_n446));
  NAND4_X1  g260(.A1(new_n440), .A2(new_n232), .A3(new_n444), .A4(new_n237), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  XOR2_X1   g263(.A(new_n449), .B(KEYINPUT8), .Z(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT83), .B1(new_n448), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT83), .ZN(new_n453));
  AOI211_X1 g267(.A(new_n453), .B(new_n450), .C1(new_n446), .C2(new_n447), .ZN(new_n454));
  OAI211_X1 g268(.A(new_n433), .B(new_n435), .C1(new_n452), .C2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT84), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n439), .A2(new_n441), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n444), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(new_n248), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n249), .A2(new_n250), .ZN(new_n461));
  OAI211_X1 g275(.A(new_n447), .B(new_n449), .C1(new_n460), .C2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n447), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n444), .A2(new_n440), .B1(new_n232), .B2(new_n237), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n451), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n453), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n448), .A2(KEYINPUT83), .A3(new_n451), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g282(.A1(new_n435), .A2(new_n433), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(KEYINPUT84), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n457), .A2(new_n462), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(new_n434), .B(new_n431), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n447), .B1(new_n460), .B2(new_n461), .ZN(new_n473));
  INV_X1    g287(.A(new_n449), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n475), .A2(KEYINPUT6), .A3(new_n462), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n473), .A2(new_n477), .A3(new_n474), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n472), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n479), .A2(new_n306), .ZN(new_n480));
  OAI21_X1  g294(.A(G210), .B1(G237), .B2(G902), .ZN(new_n481));
  AND3_X1   g295(.A1(new_n471), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n481), .B1(new_n471), .B2(new_n480), .ZN(new_n483));
  NOR2_X1   g297(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g298(.A(G214), .B1(G237), .B2(G902), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n428), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n471), .A2(new_n480), .ZN(new_n488));
  INV_X1    g302(.A(new_n481), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n471), .A2(new_n480), .A3(new_n481), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(KEYINPUT85), .A3(new_n485), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n427), .B1(new_n487), .B2(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT76), .ZN(new_n495));
  INV_X1    g309(.A(new_n375), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n383), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT23), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n437), .B2(G128), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n208), .A2(KEYINPUT23), .A3(G119), .ZN(new_n500));
  OAI211_X1 g314(.A(new_n499), .B(new_n500), .C1(G119), .C2(new_n208), .ZN(new_n501));
  XNOR2_X1  g315(.A(G119), .B(G128), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  OAI22_X1  g317(.A1(new_n501), .A2(G110), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n497), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n389), .A2(new_n391), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n501), .A2(G110), .B1(new_n502), .B2(new_n503), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n266), .A2(G221), .A3(G234), .ZN(new_n510));
  XNOR2_X1  g324(.A(new_n510), .B(KEYINPUT74), .ZN(new_n511));
  XNOR2_X1  g325(.A(KEYINPUT22), .B(G137), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n495), .B1(new_n509), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g329(.A1(new_n497), .A2(new_n504), .B1(new_n506), .B2(new_n507), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n516), .A2(KEYINPUT76), .A3(new_n513), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n509), .A2(KEYINPUT75), .A3(new_n514), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT75), .ZN(new_n519));
  OAI21_X1  g333(.A(new_n519), .B1(new_n516), .B2(new_n513), .ZN(new_n520));
  AOI22_X1  g334(.A1(new_n515), .A2(new_n517), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT25), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n521), .A2(new_n522), .A3(new_n306), .ZN(new_n523));
  INV_X1    g337(.A(G234), .ZN(new_n524));
  OAI21_X1  g338(.A(G217), .B1(new_n524), .B2(G902), .ZN(new_n525));
  XNOR2_X1  g339(.A(new_n525), .B(KEYINPUT72), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT73), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n523), .A2(new_n527), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n522), .B1(new_n521), .B2(new_n306), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g344(.A(new_n521), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n526), .A2(new_n306), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(G472), .A2(G902), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n203), .B1(G134), .B2(G137), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n317), .B2(G137), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n204), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT67), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n204), .A2(KEYINPUT67), .A3(new_n537), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n540), .A2(new_n541), .A3(new_n254), .ZN(new_n542));
  INV_X1    g356(.A(new_n459), .ZN(new_n543));
  INV_X1    g357(.A(new_n204), .ZN(new_n544));
  INV_X1    g358(.A(new_n200), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n203), .B1(new_n545), .B2(new_n202), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n245), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n542), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n359), .A2(new_n266), .A3(G210), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n549), .B(KEYINPUT27), .ZN(new_n550));
  XNOR2_X1  g364(.A(KEYINPUT26), .B(G101), .ZN(new_n551));
  XNOR2_X1  g365(.A(new_n550), .B(new_n551), .ZN(new_n552));
  AND3_X1   g366(.A1(new_n548), .A2(KEYINPUT69), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(KEYINPUT69), .B1(new_n548), .B2(new_n552), .ZN(new_n554));
  OR2_X1    g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT31), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT30), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n259), .A2(new_n538), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n244), .B1(new_n201), .B2(new_n204), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT66), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n542), .A2(KEYINPUT30), .A3(new_n547), .ZN(new_n563));
  OAI211_X1 g377(.A(KEYINPUT66), .B(new_n557), .C1(new_n558), .C2(new_n559), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n562), .A2(new_n459), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n565), .A2(KEYINPUT68), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n565), .A2(KEYINPUT68), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n555), .B(new_n556), .C1(new_n566), .C2(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT71), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n553), .A2(new_n554), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n254), .A2(new_n204), .A3(new_n537), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n547), .ZN(new_n572));
  AOI21_X1  g386(.A(KEYINPUT66), .B1(new_n572), .B2(new_n557), .ZN(new_n573));
  INV_X1    g387(.A(new_n564), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT68), .ZN(new_n576));
  NAND4_X1  g390(.A1(new_n575), .A2(new_n576), .A3(new_n459), .A4(new_n563), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n565), .A2(KEYINPUT68), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n570), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT71), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n579), .A2(new_n580), .A3(new_n556), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n569), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT70), .B1(new_n579), .B2(new_n556), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n555), .B1(new_n566), .B2(new_n567), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT70), .ZN(new_n585));
  NAND3_X1  g399(.A1(new_n584), .A2(new_n585), .A3(KEYINPUT31), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n548), .B(KEYINPUT28), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n572), .A2(new_n459), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n552), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n583), .A2(new_n586), .A3(new_n591), .ZN(new_n592));
  OAI211_X1 g406(.A(KEYINPUT32), .B(new_n535), .C1(new_n582), .C2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n589), .A2(new_n590), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n548), .B1(new_n566), .B2(new_n567), .ZN(new_n595));
  AOI211_X1 g409(.A(KEYINPUT29), .B(new_n594), .C1(new_n590), .C2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n542), .A2(new_n547), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n459), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n587), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n552), .A2(KEYINPUT29), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n306), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n596), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n593), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n569), .A2(new_n581), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n604), .A2(new_n583), .A3(new_n586), .A4(new_n591), .ZN(new_n605));
  AOI21_X1  g419(.A(KEYINPUT32), .B1(new_n605), .B2(new_n535), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n494), .B(new_n534), .C1(new_n603), .C2(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n607), .B(G101), .ZN(G3));
  OAI21_X1  g422(.A(new_n306), .B1(new_n582), .B2(new_n592), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n609), .A2(G472), .B1(new_n535), .B2(new_n605), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n610), .A2(new_n534), .A3(new_n290), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT100), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n486), .B1(new_n482), .B2(KEYINPUT101), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT101), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n490), .A2(new_n614), .A3(new_n491), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n613), .A2(new_n615), .A3(new_n303), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n352), .A2(G478), .ZN(new_n617));
  INV_X1    g431(.A(new_n351), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT33), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n337), .A2(new_n346), .A3(new_n349), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n618), .A2(new_n619), .A3(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(KEYINPUT33), .B1(new_n350), .B2(new_n351), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(G478), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(G478), .A2(G902), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n617), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n426), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT102), .ZN(new_n627));
  OR2_X1    g441(.A1(new_n626), .A2(KEYINPUT102), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n616), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n612), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT103), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  AND3_X1   g447(.A1(new_n420), .A2(new_n424), .A3(new_n421), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n424), .B1(new_n420), .B2(new_n421), .ZN(new_n635));
  OAI22_X1  g449(.A1(new_n634), .A2(new_n635), .B1(new_n408), .B2(new_n407), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n358), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n616), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n612), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT35), .B(G107), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G9));
  NOR2_X1   g456(.A1(new_n514), .A2(KEYINPUT36), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n509), .ZN(new_n644));
  INV_X1    g458(.A(new_n532), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n528), .B2(new_n529), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n647), .A2(new_n358), .A3(new_n303), .A4(new_n426), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n648), .B1(new_n487), .B2(new_n493), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n610), .A2(new_n290), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT37), .B(G110), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G12));
  OAI21_X1  g466(.A(new_n535), .B1(new_n582), .B2(new_n592), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT32), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n655), .A2(new_n593), .A3(new_n602), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n485), .B1(new_n491), .B2(new_n614), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n484), .B2(new_n614), .ZN(new_n658));
  INV_X1    g472(.A(new_n647), .ZN(new_n659));
  INV_X1    g473(.A(G900), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n298), .B1(new_n660), .B2(new_n301), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n658), .A2(new_n662), .A3(new_n290), .A4(new_n637), .ZN(new_n663));
  INV_X1    g477(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n656), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G128), .ZN(G30));
  AOI21_X1  g480(.A(new_n552), .B1(new_n598), .B2(new_n548), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n306), .B1(new_n579), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(G472), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n655), .A2(new_n593), .A3(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n659), .A2(new_n485), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n358), .A2(new_n426), .ZN(new_n674));
  AOI21_X1  g488(.A(KEYINPUT104), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n673), .A2(KEYINPUT104), .A3(new_n674), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n492), .B(KEYINPUT38), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NOR3_X1   g492(.A1(new_n671), .A2(new_n675), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(KEYINPUT105), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n661), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n290), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT106), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n679), .A2(KEYINPUT105), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT107), .B(G143), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G45));
  INV_X1    g503(.A(new_n658), .ZN(new_n690));
  INV_X1    g504(.A(new_n661), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n290), .A2(new_n647), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n626), .ZN(new_n693));
  NOR3_X1   g507(.A1(new_n690), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n656), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G146), .ZN(G48));
  AOI22_X1  g510(.A1(new_n283), .A2(new_n275), .B1(new_n285), .B2(new_n270), .ZN(new_n697));
  OAI21_X1  g511(.A(G469), .B1(new_n697), .B2(G902), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n289), .A2(new_n698), .A3(new_n188), .ZN(new_n699));
  INV_X1    g513(.A(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n534), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n629), .B(new_n702), .C1(new_n603), .C2(new_n606), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT108), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT108), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n656), .A2(new_n705), .A3(new_n629), .A4(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n704), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(KEYINPUT41), .B(G113), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G15));
  OAI211_X1 g523(.A(new_n639), .B(new_n702), .C1(new_n603), .C2(new_n606), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G116), .ZN(G18));
  NAND2_X1  g525(.A1(new_n658), .A2(new_n699), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n712), .A2(new_n648), .ZN(new_n713));
  OAI21_X1  g527(.A(new_n713), .B1(new_n606), .B2(new_n603), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  INV_X1    g529(.A(new_n535), .ZN(new_n716));
  AOI22_X1  g530(.A1(new_n584), .A2(KEYINPUT31), .B1(new_n599), .B2(new_n590), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n716), .B1(new_n604), .B2(new_n717), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n718), .B1(new_n609), .B2(G472), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n613), .A2(new_n615), .A3(new_n674), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n720), .A2(new_n302), .A3(new_n700), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n719), .A2(new_n721), .A3(new_n534), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NOR3_X1   g537(.A1(new_n426), .A2(new_n625), .A3(new_n661), .ZN(new_n724));
  AND4_X1   g538(.A1(new_n615), .A2(new_n724), .A3(new_n613), .A4(new_n699), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n719), .A2(new_n647), .A3(new_n725), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G125), .ZN(G27));
  INV_X1    g541(.A(KEYINPUT111), .ZN(new_n728));
  AOI21_X1  g542(.A(new_n728), .B1(new_n653), .B2(new_n654), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n603), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n606), .A2(new_n728), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n701), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n733), .B1(new_n277), .B2(G469), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n277), .A2(new_n733), .A3(G469), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(G469), .A2(G902), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT109), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n739), .B1(new_n287), .B2(new_n288), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n189), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n492), .A2(new_n486), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n741), .A2(new_n724), .A3(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  AND2_X1   g559(.A1(new_n741), .A2(new_n742), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n656), .A2(new_n534), .A3(new_n724), .A4(new_n746), .ZN(new_n747));
  AOI22_X1  g561(.A1(new_n732), .A2(new_n745), .B1(new_n747), .B2(new_n744), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(new_n203), .ZN(G33));
  NOR2_X1   g563(.A1(new_n638), .A2(new_n661), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n656), .A2(new_n534), .A3(new_n746), .A4(new_n750), .ZN(new_n751));
  XNOR2_X1  g565(.A(new_n751), .B(G134), .ZN(G36));
  INV_X1    g566(.A(KEYINPUT112), .ZN(new_n753));
  INV_X1    g567(.A(G469), .ZN(new_n754));
  INV_X1    g568(.A(new_n277), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT45), .ZN(new_n756));
  AOI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n757), .B1(new_n756), .B2(new_n755), .ZN(new_n758));
  INV_X1    g572(.A(new_n739), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  INV_X1    g574(.A(new_n760), .ZN(new_n761));
  OAI21_X1  g575(.A(new_n753), .B1(new_n761), .B2(KEYINPUT46), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n763));
  NAND3_X1  g577(.A1(new_n760), .A2(KEYINPUT112), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(KEYINPUT46), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n762), .A2(new_n289), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n766), .A2(new_n188), .ZN(new_n767));
  INV_X1    g581(.A(new_n767), .ZN(new_n768));
  INV_X1    g582(.A(new_n610), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n636), .A2(new_n625), .ZN(new_n770));
  INV_X1    g584(.A(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT43), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n772), .A2(KEYINPUT113), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  XNOR2_X1  g588(.A(KEYINPUT113), .B(KEYINPUT43), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n774), .B1(new_n771), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n769), .A2(new_n647), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT44), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n681), .A2(new_n768), .A3(new_n742), .A4(new_n779), .ZN(new_n780));
  OR2_X1    g594(.A1(new_n777), .A2(new_n778), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G137), .ZN(G39));
  INV_X1    g597(.A(KEYINPUT47), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n767), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n766), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n742), .A2(new_n701), .A3(new_n724), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n656), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  AND2_X1   g605(.A1(new_n776), .A2(new_n298), .ZN(new_n792));
  AND2_X1   g606(.A1(new_n719), .A2(new_n534), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n742), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  AND2_X1   g610(.A1(new_n289), .A2(new_n698), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n797), .A2(new_n189), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n796), .B1(new_n787), .B2(new_n798), .ZN(new_n799));
  NOR3_X1   g613(.A1(new_n677), .A2(new_n485), .A3(new_n700), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n792), .A2(new_n793), .A3(new_n800), .ZN(new_n801));
  XOR2_X1   g615(.A(new_n801), .B(KEYINPUT50), .Z(new_n802));
  NOR4_X1   g616(.A1(new_n795), .A2(new_n701), .A3(new_n700), .A4(new_n297), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n671), .A2(new_n426), .A3(new_n625), .A4(new_n803), .ZN(new_n804));
  AOI211_X1 g618(.A(new_n659), .B(new_n718), .C1(new_n609), .C2(G472), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n795), .A2(new_n700), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n792), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AND2_X1   g621(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n799), .A2(new_n802), .A3(new_n808), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT51), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n799), .A2(new_n802), .A3(KEYINPUT51), .A4(new_n808), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n628), .A2(new_n627), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n671), .A2(new_n813), .A3(new_n803), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n294), .C1(new_n794), .C2(new_n712), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n732), .A2(new_n792), .A3(new_n806), .ZN(new_n816));
  OR2_X1    g630(.A1(new_n816), .A2(KEYINPUT48), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(KEYINPUT48), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n815), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n811), .A2(new_n812), .A3(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT118), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n820), .B(new_n821), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n593), .A2(new_n602), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n823), .B1(new_n728), .B2(new_n606), .ZN(new_n824));
  INV_X1    g638(.A(new_n731), .ZN(new_n825));
  OAI211_X1 g639(.A(new_n534), .B(new_n745), .C1(new_n824), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n747), .A2(new_n744), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(new_n743), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n805), .A2(KEYINPUT114), .A3(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT114), .ZN(new_n831));
  INV_X1    g645(.A(new_n718), .ZN(new_n832));
  AND3_X1   g646(.A1(new_n583), .A2(new_n586), .A3(new_n591), .ZN(new_n833));
  AOI21_X1  g647(.A(G902), .B1(new_n833), .B2(new_n604), .ZN(new_n834));
  INV_X1    g648(.A(G472), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n647), .B(new_n832), .C1(new_n834), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n831), .B1(new_n836), .B2(new_n743), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n830), .A2(new_n837), .ZN(new_n838));
  INV_X1    g652(.A(new_n358), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n692), .A2(new_n839), .A3(new_n636), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n656), .A2(new_n742), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n751), .A2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n828), .A2(new_n838), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g657(.A(new_n303), .B1(new_n637), .B2(new_n626), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n844), .B1(new_n487), .B2(new_n493), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n610), .A2(new_n845), .A3(new_n534), .A4(new_n290), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n846), .A2(new_n607), .A3(new_n710), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n714), .A2(new_n722), .A3(new_n650), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n849), .A2(new_n707), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n843), .A2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(new_n720), .ZN(new_n852));
  INV_X1    g666(.A(new_n736), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n740), .B1(new_n853), .B2(new_n734), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n646), .B(new_n691), .C1(new_n528), .C2(new_n529), .ZN(new_n855));
  INV_X1    g669(.A(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n854), .A2(new_n856), .A3(KEYINPUT116), .A4(new_n188), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n852), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT116), .B1(new_n741), .B2(new_n856), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n670), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n861), .A2(new_n695), .A3(new_n665), .A4(new_n726), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  XNOR2_X1  g677(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n851), .A2(KEYINPUT53), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g679(.A(KEYINPUT114), .B1(new_n805), .B2(new_n829), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n836), .A2(new_n831), .A3(new_n743), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n751), .B(new_n841), .C1(new_n866), .C2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n869), .A2(new_n707), .A3(new_n828), .A4(new_n849), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT115), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n663), .B1(new_n823), .B2(new_n655), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n609), .A2(G472), .ZN(new_n873));
  AND4_X1   g687(.A1(new_n873), .A2(new_n647), .A3(new_n725), .A4(new_n832), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n871), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n665), .A2(KEYINPUT115), .A3(new_n726), .ZN(new_n876));
  AOI22_X1  g690(.A1(new_n860), .A2(new_n670), .B1(new_n656), .B2(new_n694), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n875), .A2(KEYINPUT52), .A3(new_n876), .A4(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n862), .A2(new_n863), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT117), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT117), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n878), .A2(new_n879), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n870), .B1(new_n881), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n865), .B1(new_n884), .B2(KEYINPUT53), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(KEYINPUT54), .ZN(new_n886));
  INV_X1    g700(.A(new_n883), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n882), .B1(new_n878), .B2(new_n879), .ZN(new_n888));
  OAI211_X1 g702(.A(new_n851), .B(KEYINPUT53), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT54), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT53), .ZN(new_n891));
  XNOR2_X1  g705(.A(new_n862), .B(KEYINPUT52), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n891), .B1(new_n870), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n890), .A3(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n886), .A2(new_n894), .ZN(new_n895));
  OAI22_X1  g709(.A1(new_n822), .A2(new_n895), .B1(G952), .B2(G953), .ZN(new_n896));
  XNOR2_X1  g710(.A(new_n797), .B(KEYINPUT49), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n189), .A2(new_n486), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n897), .A2(new_n534), .A3(new_n771), .A4(new_n898), .ZN(new_n899));
  OR2_X1    g713(.A1(new_n899), .A2(new_n677), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n670), .B2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n266), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n889), .A2(new_n893), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G902), .ZN(new_n905));
  INV_X1    g719(.A(G210), .ZN(new_n906));
  NOR2_X1   g720(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n476), .A2(new_n478), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n908), .B(new_n472), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT55), .Z(new_n910));
  OR2_X1    g724(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n903), .B1(new_n907), .B2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n907), .A2(KEYINPUT119), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT119), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n915), .B1(new_n905), .B2(new_n906), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n913), .A2(new_n914), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n912), .B1(new_n917), .B2(new_n910), .ZN(G51));
  NOR2_X1   g732(.A1(new_n905), .A2(new_n758), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n748), .A2(new_n868), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n846), .A2(new_n607), .A3(new_n710), .ZN(new_n921));
  AND3_X1   g735(.A1(new_n714), .A2(new_n650), .A3(new_n722), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n707), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n920), .A2(new_n923), .A3(KEYINPUT53), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n924), .B1(new_n883), .B2(new_n881), .ZN(new_n925));
  AOI21_X1  g739(.A(KEYINPUT53), .B1(new_n851), .B2(new_n864), .ZN(new_n926));
  OAI21_X1  g740(.A(KEYINPUT54), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n927), .A2(new_n894), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n739), .B(KEYINPUT57), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n697), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n919), .B1(new_n930), .B2(KEYINPUT120), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n932));
  INV_X1    g746(.A(new_n929), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n927), .B2(new_n894), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n932), .B1(new_n934), .B2(new_n697), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n902), .B1(new_n931), .B2(new_n935), .ZN(G54));
  AND2_X1   g750(.A1(KEYINPUT58), .A2(G475), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n904), .A2(G902), .A3(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(new_n420), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n902), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND4_X1  g754(.A1(new_n904), .A2(G902), .A3(new_n420), .A4(new_n937), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n940), .B1(KEYINPUT121), .B2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n942), .B1(KEYINPUT121), .B2(new_n941), .ZN(G60));
  XOR2_X1   g757(.A(new_n624), .B(KEYINPUT59), .Z(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n886), .B2(new_n894), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n621), .A2(new_n622), .ZN(new_n946));
  INV_X1    g760(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g761(.A(KEYINPUT122), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n944), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n851), .B1(new_n887), .B2(new_n888), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n950), .A2(new_n891), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n890), .B1(new_n951), .B2(new_n865), .ZN(new_n952));
  INV_X1    g766(.A(new_n894), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n949), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT122), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n954), .A2(new_n955), .A3(new_n946), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n946), .A2(new_n944), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n902), .B1(new_n928), .B2(new_n957), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n948), .A2(new_n956), .A3(new_n958), .ZN(G63));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XOR2_X1   g774(.A(new_n960), .B(KEYINPUT60), .Z(new_n961));
  NAND2_X1  g775(.A1(new_n904), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n962), .A2(new_n531), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n904), .A2(new_n644), .A3(new_n961), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n963), .A2(new_n903), .A3(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(KEYINPUT61), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G66));
  INV_X1    g781(.A(new_n430), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n968), .B2(new_n299), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n969), .B1(new_n923), .B2(G953), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n908), .B1(G898), .B2(new_n266), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n971), .B(KEYINPUT123), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n970), .B(new_n972), .ZN(G69));
  AOI21_X1  g787(.A(new_n266), .B1(G227), .B2(G900), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n575), .A2(new_n563), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n412), .A2(new_n413), .ZN(new_n977));
  XOR2_X1   g791(.A(new_n976), .B(new_n977), .Z(new_n978));
  AND3_X1   g792(.A1(new_n768), .A2(new_n681), .A3(new_n852), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n780), .A2(new_n781), .B1(new_n979), .B2(new_n732), .ZN(new_n980));
  AND2_X1   g794(.A1(new_n790), .A2(new_n751), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n875), .A2(new_n876), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n982), .A2(new_n695), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  NAND4_X1  g798(.A1(new_n980), .A2(new_n981), .A3(new_n828), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(new_n266), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n660), .A2(G953), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n987), .B(KEYINPUT125), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n978), .B1(new_n986), .B2(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n984), .B1(new_n686), .B2(new_n685), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT124), .B1(new_n991), .B2(KEYINPUT62), .ZN(new_n992));
  OAI211_X1 g806(.A(KEYINPUT124), .B(KEYINPUT62), .C1(new_n687), .C2(new_n983), .ZN(new_n993));
  INV_X1    g807(.A(new_n993), .ZN(new_n994));
  OR2_X1    g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n638), .A2(new_n693), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n795), .A2(new_n682), .ZN(new_n997));
  NAND4_X1  g811(.A1(new_n656), .A2(new_n534), .A3(new_n996), .A4(new_n997), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n782), .A2(new_n790), .A3(new_n998), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n687), .A2(new_n983), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n999), .B1(new_n1000), .B2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(G953), .B1(new_n995), .B2(new_n1002), .ZN(new_n1003));
  INV_X1    g817(.A(new_n978), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n975), .B(new_n990), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n1002), .B1(new_n992), .B2(new_n994), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1004), .B1(new_n1006), .B2(new_n266), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n974), .B1(new_n1007), .B2(new_n989), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n1005), .A2(new_n1008), .ZN(G72));
  NAND2_X1  g823(.A1(new_n595), .A2(new_n552), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n995), .A2(new_n923), .A3(new_n1002), .ZN(new_n1011));
  XNOR2_X1  g825(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1012));
  NOR2_X1   g826(.A1(new_n835), .A2(new_n306), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1010), .B1(new_n1011), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1014), .B1(new_n985), .B2(new_n850), .ZN(new_n1016));
  NOR2_X1   g830(.A1(new_n595), .A2(new_n552), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n902), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n885), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n595), .A2(new_n590), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1014), .B1(new_n1020), .B2(new_n579), .ZN(new_n1021));
  XNOR2_X1  g835(.A(new_n1021), .B(KEYINPUT127), .ZN(new_n1022));
  OAI21_X1  g836(.A(new_n1018), .B1(new_n1019), .B2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g837(.A1(new_n1015), .A2(new_n1023), .ZN(G57));
endmodule


