//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 1 1 0 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:04 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n757, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(G137), .ZN(new_n191));
  INV_X1    g005(.A(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n192), .A2(KEYINPUT11), .A3(G134), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n191), .A3(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G131), .ZN(new_n195));
  INV_X1    g009(.A(G131), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n190), .A2(new_n193), .A3(new_n196), .A4(new_n191), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n199), .A2(KEYINPUT65), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT65), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n202), .A3(G143), .ZN(new_n203));
  INV_X1    g017(.A(G143), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G143), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G146), .ZN(new_n208));
  NAND4_X1  g022(.A1(new_n203), .A2(new_n208), .A3(KEYINPUT0), .A4(G128), .ZN(new_n209));
  XOR2_X1   g023(.A(KEYINPUT0), .B(G128), .Z(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n205), .B2(new_n207), .ZN(new_n211));
  AOI21_X1  g025(.A(G143), .B1(new_n200), .B2(new_n202), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n198), .A2(new_n209), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT68), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n198), .A2(KEYINPUT68), .A3(new_n209), .A4(new_n213), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT2), .B(G113), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT67), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT2), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(G113), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n223), .A2(new_n225), .A3(new_n220), .ZN(new_n226));
  XNOR2_X1  g040(.A(G116), .B(G119), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n221), .A2(new_n226), .B1(KEYINPUT66), .B2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n227), .A2(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n223), .A2(new_n225), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT67), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n219), .A2(new_n220), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n228), .A2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT1), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n203), .A2(new_n208), .A3(new_n236), .A4(G128), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n211), .A2(new_n212), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  AOI21_X1  g053(.A(new_n239), .B1(new_n203), .B2(KEYINPUT1), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n237), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n191), .ZN(new_n242));
  NOR2_X1   g056(.A1(new_n189), .A2(G137), .ZN(new_n243));
  OAI21_X1  g057(.A(G131), .B1(new_n242), .B2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n241), .A2(new_n244), .A3(new_n197), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n218), .A2(new_n235), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(KEYINPUT69), .B(G237), .ZN(new_n247));
  INV_X1    g061(.A(G953), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(G210), .A3(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(new_n249), .B(KEYINPUT27), .ZN(new_n250));
  XNOR2_X1  g064(.A(KEYINPUT26), .B(G101), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n250), .B(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT30), .ZN(new_n253));
  AND3_X1   g067(.A1(new_n245), .A2(new_n253), .A3(new_n214), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n213), .A2(new_n209), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT68), .B1(new_n255), .B2(new_n198), .ZN(new_n256));
  INV_X1    g070(.A(new_n217), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n245), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n254), .B1(new_n258), .B2(KEYINPUT30), .ZN(new_n259));
  OAI211_X1 g073(.A(new_n246), .B(new_n252), .C1(new_n259), .C2(new_n235), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT70), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n245), .A2(new_n253), .A3(new_n214), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n244), .A2(new_n197), .ZN(new_n263));
  XNOR2_X1  g077(.A(KEYINPUT65), .B(G146), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n236), .B1(new_n264), .B2(G143), .ZN(new_n265));
  OAI22_X1  g079(.A1(new_n265), .A2(new_n239), .B1(new_n211), .B2(new_n212), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n263), .B1(new_n266), .B2(new_n237), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n216), .B2(new_n217), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n262), .B1(new_n268), .B2(new_n253), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n269), .A2(new_n234), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT70), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n270), .A2(new_n271), .A3(new_n246), .A4(new_n252), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n261), .A2(KEYINPUT31), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n252), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n245), .A2(new_n235), .A3(new_n214), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT28), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(new_n235), .B1(new_n245), .B2(new_n214), .ZN(new_n278));
  INV_X1    g092(.A(new_n278), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n276), .B1(new_n246), .B2(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(KEYINPUT71), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n277), .B1(new_n280), .B2(new_n281), .ZN(new_n282));
  AOI21_X1  g096(.A(new_n278), .B1(new_n268), .B2(new_n235), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n283), .A2(KEYINPUT71), .A3(new_n276), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n274), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  AOI211_X1 g099(.A(new_n234), .B(new_n267), .C1(new_n216), .C2(new_n217), .ZN(new_n286));
  AOI211_X1 g100(.A(new_n274), .B(new_n286), .C1(new_n269), .C2(new_n234), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT31), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n285), .A2(new_n289), .ZN(new_n290));
  OAI21_X1  g104(.A(new_n187), .B1(new_n273), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT32), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n187), .ZN(new_n294));
  OAI21_X1  g108(.A(KEYINPUT71), .B1(new_n283), .B2(new_n276), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n281), .B(KEYINPUT28), .C1(new_n286), .C2(new_n278), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n295), .A2(new_n296), .A3(new_n277), .ZN(new_n297));
  AOI22_X1  g111(.A1(new_n297), .A2(new_n274), .B1(new_n287), .B2(new_n288), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n261), .A2(KEYINPUT31), .A3(new_n272), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(KEYINPUT32), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n270), .A2(new_n246), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(new_n274), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT29), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n303), .B(new_n304), .C1(new_n297), .C2(new_n274), .ZN(new_n305));
  INV_X1    g119(.A(G902), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n235), .B1(new_n218), .B2(new_n245), .ZN(new_n307));
  OAI21_X1  g121(.A(KEYINPUT28), .B1(new_n286), .B2(new_n307), .ZN(new_n308));
  NAND4_X1  g122(.A1(new_n308), .A2(KEYINPUT29), .A3(new_n252), .A4(new_n277), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G472), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n293), .A2(new_n301), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT23), .ZN(new_n313));
  INV_X1    g127(.A(G119), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n313), .B1(new_n314), .B2(G128), .ZN(new_n315));
  OAI21_X1  g129(.A(KEYINPUT72), .B1(new_n314), .B2(G128), .ZN(new_n316));
  XNOR2_X1  g130(.A(new_n315), .B(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G119), .B(G128), .ZN(new_n318));
  XOR2_X1   g132(.A(KEYINPUT24), .B(G110), .Z(new_n319));
  OAI22_X1  g133(.A1(new_n317), .A2(G110), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  XNOR2_X1  g134(.A(G125), .B(G140), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n323), .A2(KEYINPUT16), .A3(G140), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(G146), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n264), .A2(new_n321), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n320), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g141(.A(G146), .B1(new_n322), .B2(new_n324), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT74), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n325), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n330), .B1(new_n329), .B2(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n319), .A2(new_n318), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT73), .ZN(new_n333));
  OAI21_X1  g147(.A(G110), .B1(new_n317), .B2(new_n333), .ZN(new_n334));
  OR2_X1    g148(.A1(new_n315), .A2(new_n316), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n315), .A2(new_n316), .ZN(new_n336));
  AOI21_X1  g150(.A(KEYINPUT73), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n332), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n327), .B1(new_n331), .B2(new_n338), .ZN(new_n339));
  XNOR2_X1  g153(.A(KEYINPUT22), .B(G137), .ZN(new_n340));
  AND3_X1   g154(.A1(new_n248), .A2(G221), .A3(G234), .ZN(new_n341));
  XOR2_X1   g155(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n339), .A2(new_n343), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n327), .B(new_n342), .C1(new_n331), .C2(new_n338), .ZN(new_n345));
  AND2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G217), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n347), .B1(G234), .B2(new_n306), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n348), .A2(G902), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n349), .B(KEYINPUT75), .Z(new_n350));
  INV_X1    g164(.A(new_n350), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n346), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT76), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT76), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n346), .A2(new_n354), .A3(new_n351), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(new_n348), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n344), .A2(new_n306), .A3(new_n345), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT25), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND4_X1  g174(.A1(new_n344), .A2(KEYINPUT25), .A3(new_n306), .A4(new_n345), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n357), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  OR3_X1    g176(.A1(new_n356), .A2(KEYINPUT77), .A3(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT77), .B1(new_n356), .B2(new_n362), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n312), .A2(KEYINPUT78), .A3(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT78), .B1(new_n312), .B2(new_n365), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(new_n198), .ZN(new_n369));
  XNOR2_X1  g183(.A(G104), .B(G107), .ZN(new_n370));
  INV_X1    g184(.A(G101), .ZN(new_n371));
  OAI21_X1  g185(.A(KEYINPUT82), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G104), .ZN(new_n373));
  OAI21_X1  g187(.A(KEYINPUT3), .B1(new_n373), .B2(G107), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT3), .ZN(new_n375));
  INV_X1    g189(.A(G107), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(G104), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n373), .A2(G107), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n374), .A2(new_n377), .A3(new_n371), .A4(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT82), .ZN(new_n380));
  NOR2_X1   g194(.A1(new_n373), .A2(G107), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n376), .A2(G104), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n380), .B(G101), .C1(new_n381), .C2(new_n382), .ZN(new_n383));
  AND3_X1   g197(.A1(new_n372), .A2(new_n379), .A3(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT64), .B(G143), .ZN(new_n385));
  OAI21_X1  g199(.A(KEYINPUT1), .B1(new_n385), .B2(G146), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n386), .A2(G128), .B1(new_n203), .B2(new_n208), .ZN(new_n387));
  OAI21_X1  g201(.A(new_n237), .B1(new_n387), .B2(KEYINPUT83), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n203), .A2(new_n208), .ZN(new_n389));
  NOR2_X1   g203(.A1(new_n211), .A2(new_n236), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n389), .B(KEYINPUT83), .C1(new_n390), .C2(new_n239), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n384), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n241), .A2(new_n384), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n369), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT84), .B1(new_n396), .B2(KEYINPUT12), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT84), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT12), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT83), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n206), .A2(G143), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n204), .A2(KEYINPUT64), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n199), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n239), .B1(new_n403), .B2(KEYINPUT1), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n203), .A2(new_n208), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n400), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n237), .A3(new_n391), .ZN(new_n407));
  AOI21_X1  g221(.A(new_n394), .B1(new_n407), .B2(new_n384), .ZN(new_n408));
  OAI211_X1 g222(.A(new_n398), .B(new_n399), .C1(new_n408), .C2(new_n369), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n396), .A2(KEYINPUT12), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n397), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT10), .ZN(new_n412));
  INV_X1    g226(.A(new_n384), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n412), .ZN(new_n414));
  AOI22_X1  g228(.A1(new_n393), .A2(new_n412), .B1(new_n241), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n374), .A2(new_n377), .A3(new_n378), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(G101), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n417), .A2(KEYINPUT4), .A3(new_n379), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT80), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  NAND4_X1  g234(.A1(new_n417), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n379), .ZN(new_n421));
  INV_X1    g235(.A(new_n417), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n420), .A2(new_n255), .A3(new_n421), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT81), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI22_X1  g241(.A1(new_n418), .A2(new_n419), .B1(new_n422), .B2(new_n423), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n428), .A2(KEYINPUT81), .A3(new_n255), .A4(new_n421), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n415), .A2(new_n430), .A3(new_n369), .ZN(new_n431));
  XNOR2_X1  g245(.A(G110), .B(G140), .ZN(new_n432));
  AND2_X1   g246(.A1(new_n248), .A2(G227), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n411), .A2(new_n431), .A3(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n431), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n369), .B1(new_n415), .B2(new_n430), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n434), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n436), .B2(new_n439), .ZN(new_n440));
  XOR2_X1   g254(.A(KEYINPUT87), .B(G469), .Z(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT85), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n411), .A2(new_n444), .A3(new_n431), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n444), .B1(new_n411), .B2(new_n431), .ZN(new_n446));
  XOR2_X1   g260(.A(new_n434), .B(KEYINPUT79), .Z(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  NOR3_X1   g262(.A1(new_n445), .A2(new_n446), .A3(new_n448), .ZN(new_n449));
  AND3_X1   g263(.A1(new_n431), .A2(KEYINPUT86), .A3(new_n435), .ZN(new_n450));
  AOI21_X1  g264(.A(KEYINPUT86), .B1(new_n431), .B2(new_n435), .ZN(new_n451));
  NOR3_X1   g265(.A1(new_n450), .A2(new_n451), .A3(new_n438), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n306), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n443), .B1(new_n453), .B2(G469), .ZN(new_n454));
  INV_X1    g268(.A(G221), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT9), .B(G234), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n455), .B1(new_n457), .B2(new_n306), .ZN(new_n458));
  OAI21_X1  g272(.A(KEYINPUT88), .B1(new_n454), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n411), .A2(new_n431), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n448), .B1(new_n460), .B2(KEYINPUT85), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n411), .A2(new_n444), .A3(new_n431), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n452), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(G469), .B1(new_n463), .B2(G902), .ZN(new_n464));
  AOI21_X1  g278(.A(new_n458), .B1(new_n464), .B2(new_n442), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT88), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NOR3_X1   g281(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  AND2_X1   g283(.A1(KEYINPUT69), .A2(G237), .ZN(new_n470));
  NOR2_X1   g284(.A1(KEYINPUT69), .A2(G237), .ZN(new_n471));
  OAI211_X1 g285(.A(G214), .B(new_n248), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n385), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n247), .A2(G143), .A3(G214), .A4(new_n248), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT18), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n476), .B1(new_n477), .B2(new_n196), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n326), .B1(new_n199), .B2(new_n321), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n475), .A2(G131), .ZN(new_n480));
  OAI211_X1 g294(.A(new_n478), .B(new_n479), .C1(new_n477), .C2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(KEYINPUT92), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n475), .A2(KEYINPUT92), .A3(G131), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n483), .A2(new_n484), .B1(new_n196), .B2(new_n476), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n321), .A2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT19), .ZN(new_n488));
  INV_X1    g302(.A(new_n264), .ZN(new_n489));
  OAI21_X1  g303(.A(new_n325), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(new_n481), .B1(new_n485), .B2(new_n490), .ZN(new_n491));
  XNOR2_X1  g305(.A(G113), .B(G122), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(new_n373), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n476), .A2(new_n196), .ZN(new_n496));
  INV_X1    g310(.A(KEYINPUT17), .ZN(new_n497));
  AOI21_X1  g311(.A(KEYINPUT92), .B1(new_n475), .B2(G131), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n482), .B(new_n196), .C1(new_n473), .C2(new_n474), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n496), .B(new_n497), .C1(new_n498), .C2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n483), .A2(KEYINPUT17), .A3(new_n484), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n500), .A2(new_n501), .A3(new_n331), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n502), .A2(new_n493), .A3(new_n481), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n469), .B1(new_n495), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n495), .A2(new_n503), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT94), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g321(.A1(G475), .A2(G902), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n495), .A2(new_n503), .A3(KEYINPUT94), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n504), .B1(new_n510), .B2(KEYINPUT20), .ZN(new_n511));
  INV_X1    g325(.A(G475), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n502), .A2(new_n481), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n494), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n503), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n512), .B1(new_n515), .B2(new_n306), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(G234), .A2(G237), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n518), .A2(G952), .A3(new_n248), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT21), .B(G898), .Z(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(G902), .A3(G953), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n519), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  XOR2_X1   g336(.A(new_n522), .B(KEYINPUT98), .Z(new_n523));
  INV_X1    g337(.A(KEYINPUT97), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n385), .A2(G128), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n239), .A2(G143), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(KEYINPUT13), .A3(new_n526), .ZN(new_n527));
  OAI211_X1 g341(.A(new_n527), .B(G134), .C1(KEYINPUT13), .C2(new_n525), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n525), .A2(new_n189), .A3(new_n526), .ZN(new_n529));
  INV_X1    g343(.A(G122), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n530), .A2(G116), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n531), .A2(KEYINPUT95), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT95), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(G116), .B2(new_n530), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G116), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n536), .A2(G122), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n535), .A2(new_n376), .A3(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n376), .B1(new_n535), .B2(new_n537), .ZN(new_n540));
  OAI211_X1 g354(.A(new_n528), .B(new_n529), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n525), .A2(new_n526), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(G134), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(new_n529), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n537), .A2(KEYINPUT14), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n530), .A2(KEYINPUT14), .A3(G116), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n545), .B(new_n546), .C1(new_n532), .C2(new_n534), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT96), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n547), .A2(new_n548), .A3(G107), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n548), .B1(new_n547), .B2(G107), .ZN(new_n550));
  OAI211_X1 g364(.A(new_n544), .B(new_n538), .C1(new_n549), .C2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n524), .B1(new_n541), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n541), .A2(new_n551), .A3(new_n524), .ZN(new_n554));
  NOR3_X1   g368(.A1(new_n456), .A2(new_n347), .A3(G953), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n553), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n555), .ZN(new_n557));
  INV_X1    g371(.A(new_n554), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n557), .B1(new_n558), .B2(new_n552), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n556), .A2(new_n559), .A3(new_n306), .ZN(new_n560));
  INV_X1    g374(.A(G478), .ZN(new_n561));
  NOR2_X1   g375(.A1(new_n561), .A2(KEYINPUT15), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n562), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n556), .A2(new_n559), .A3(new_n306), .A4(new_n564), .ZN(new_n565));
  AND2_X1   g379(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n517), .A2(new_n523), .A3(new_n566), .ZN(new_n567));
  OAI21_X1  g381(.A(G214), .B1(G237), .B2(G902), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT90), .ZN(new_n569));
  NAND4_X1  g383(.A1(new_n420), .A2(new_n234), .A3(new_n421), .A4(new_n424), .ZN(new_n570));
  OR3_X1    g384(.A1(new_n536), .A2(KEYINPUT5), .A3(G119), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT89), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n222), .B1(new_n227), .B2(KEYINPUT5), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n572), .A2(new_n573), .B1(new_n227), .B2(new_n230), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n384), .ZN(new_n575));
  XNOR2_X1  g389(.A(G110), .B(G122), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n577), .A2(KEYINPUT6), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n576), .B1(new_n570), .B2(new_n575), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n569), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n579), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n581), .A2(KEYINPUT90), .A3(KEYINPUT6), .A4(new_n577), .ZN(new_n582));
  OR2_X1    g396(.A1(new_n255), .A2(new_n323), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n266), .A2(new_n323), .A3(new_n237), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n248), .A2(G224), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT91), .Z(new_n586));
  AND3_X1   g400(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n583), .B2(new_n584), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT6), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n579), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n580), .A2(new_n582), .A3(new_n589), .A4(new_n591), .ZN(new_n592));
  XOR2_X1   g406(.A(new_n576), .B(KEYINPUT8), .Z(new_n593));
  OR2_X1    g407(.A1(new_n574), .A2(new_n384), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n593), .B1(new_n594), .B2(new_n575), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n583), .A2(new_n584), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n585), .A2(KEYINPUT7), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n583), .A2(new_n584), .A3(new_n597), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n595), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  AOI21_X1  g415(.A(G902), .B1(new_n601), .B2(new_n577), .ZN(new_n602));
  OAI21_X1  g416(.A(G210), .B1(G237), .B2(G902), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n592), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n603), .B1(new_n592), .B2(new_n602), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n568), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n567), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n459), .A2(new_n467), .A3(new_n608), .ZN(new_n609));
  NOR2_X1   g423(.A1(new_n368), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n371), .ZN(G3));
  AOI211_X1 g425(.A(KEYINPUT88), .B(new_n458), .C1(new_n464), .C2(new_n442), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n460), .A2(KEYINPUT85), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n613), .A2(new_n462), .A3(new_n447), .ZN(new_n614));
  OR3_X1    g428(.A1(new_n450), .A2(new_n451), .A3(new_n438), .ZN(new_n615));
  AOI21_X1  g429(.A(G902), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(G469), .ZN(new_n617));
  OAI21_X1  g431(.A(new_n442), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n458), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n466), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n612), .A2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n516), .ZN(new_n622));
  AND2_X1   g436(.A1(new_n510), .A2(KEYINPUT20), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n622), .B1(new_n623), .B2(new_n504), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n556), .A2(new_n559), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT33), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND4_X1  g442(.A1(new_n556), .A2(new_n559), .A3(new_n625), .A4(KEYINPUT33), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(G478), .A3(new_n306), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n560), .A2(new_n561), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n624), .A2(new_n633), .ZN(new_n634));
  OAI211_X1 g448(.A(new_n568), .B(new_n523), .C1(new_n604), .C2(new_n605), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(KEYINPUT99), .A2(G472), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n298), .A2(new_n299), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n637), .B1(new_n638), .B2(new_n306), .ZN(new_n639));
  INV_X1    g453(.A(new_n637), .ZN(new_n640));
  AOI211_X1 g454(.A(G902), .B(new_n640), .C1(new_n298), .C2(new_n299), .ZN(new_n641));
  OR2_X1    g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n363), .A2(new_n364), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g458(.A1(new_n621), .A2(new_n636), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g459(.A(new_n645), .B(G104), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NOR2_X1   g462(.A1(new_n566), .A2(new_n516), .ZN(new_n649));
  AND2_X1   g463(.A1(new_n507), .A2(new_n509), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n468), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n510), .A2(KEYINPUT102), .A3(KEYINPUT20), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g467(.A(KEYINPUT102), .B1(new_n510), .B2(KEYINPUT20), .ZN(new_n654));
  OAI21_X1  g468(.A(new_n649), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n655), .A2(new_n635), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n621), .A2(new_n644), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(new_n376), .ZN(new_n658));
  XNOR2_X1  g472(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G9));
  INV_X1    g474(.A(new_n339), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT36), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n661), .B1(new_n662), .B2(new_n342), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n339), .A2(KEYINPUT36), .A3(new_n343), .ZN(new_n664));
  NOR3_X1   g478(.A1(new_n663), .A2(new_n664), .A3(new_n350), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n362), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n642), .A2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n459), .A2(new_n467), .A3(new_n667), .A4(new_n608), .ZN(new_n668));
  XOR2_X1   g482(.A(KEYINPUT37), .B(G110), .Z(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G12));
  INV_X1    g484(.A(new_n666), .ZN(new_n671));
  AND3_X1   g485(.A1(new_n312), .A2(new_n607), .A3(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n519), .B(KEYINPUT104), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n673), .B1(G900), .B2(new_n521), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT105), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n649), .B(new_n676), .C1(new_n653), .C2(new_n654), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n672), .A2(new_n459), .A3(new_n467), .A4(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(G128), .ZN(G30));
  XOR2_X1   g494(.A(new_n675), .B(KEYINPUT39), .Z(new_n681));
  NAND3_X1  g495(.A1(new_n459), .A2(new_n467), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  OAI21_X1  g497(.A(new_n274), .B1(new_n286), .B2(new_n307), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n261), .A2(new_n272), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(new_n306), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n686), .A2(G472), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n293), .A2(new_n301), .A3(new_n687), .ZN(new_n688));
  NOR2_X1   g502(.A1(new_n604), .A2(new_n605), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT38), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n568), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n362), .A2(new_n692), .A3(new_n665), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n563), .A2(new_n565), .ZN(new_n694));
  OAI211_X1 g508(.A(new_n693), .B(new_n694), .C1(new_n511), .C2(new_n516), .ZN(new_n695));
  INV_X1    g509(.A(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n688), .A2(new_n691), .A3(new_n696), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n697), .B(KEYINPUT106), .ZN(new_n698));
  INV_X1    g512(.A(KEYINPUT40), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n459), .A2(new_n467), .A3(new_n699), .A4(new_n681), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n683), .A2(new_n698), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(new_n385), .Z(G45));
  AND3_X1   g516(.A1(new_n624), .A2(new_n633), .A3(new_n676), .ZN(new_n703));
  AND4_X1   g517(.A1(new_n312), .A2(new_n703), .A3(new_n607), .A4(new_n671), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(new_n459), .A3(new_n467), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G146), .ZN(G48));
  XNOR2_X1  g520(.A(new_n300), .B(new_n292), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n643), .B1(new_n707), .B2(new_n311), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n440), .A2(new_n617), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n709), .A2(new_n619), .A3(new_n442), .ZN(new_n710));
  INV_X1    g524(.A(new_n710), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n708), .A2(new_n636), .A3(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT41), .B(G113), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G15));
  NAND3_X1  g528(.A1(new_n708), .A2(new_n656), .A3(new_n711), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G116), .ZN(G18));
  AND3_X1   g530(.A1(new_n312), .A2(new_n567), .A3(new_n671), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n710), .A2(new_n606), .ZN(new_n718));
  AND2_X1   g532(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n314), .ZN(G21));
  NAND2_X1  g534(.A1(new_n308), .A2(new_n277), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(new_n274), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n289), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n187), .B1(new_n273), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n356), .A2(new_n362), .ZN(new_n725));
  AOI21_X1  g539(.A(G902), .B1(new_n298), .B2(new_n299), .ZN(new_n726));
  INV_X1    g540(.A(G472), .ZN(new_n727));
  OAI211_X1 g541(.A(new_n724), .B(new_n725), .C1(new_n726), .C2(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT107), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n638), .A2(new_n306), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(G472), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n732), .A2(KEYINPUT107), .A3(new_n725), .A4(new_n724), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n624), .A2(new_n607), .A3(new_n694), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n709), .A2(new_n619), .A3(new_n442), .A4(new_n523), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n734), .A2(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(new_n530), .ZN(G24));
  NAND3_X1  g553(.A1(new_n624), .A2(new_n633), .A3(new_n676), .ZN(new_n740));
  OAI211_X1 g554(.A(new_n724), .B(new_n671), .C1(new_n726), .C2(new_n727), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n718), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G125), .ZN(G27));
  NOR3_X1   g558(.A1(new_n604), .A2(new_n605), .A3(new_n692), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n465), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n703), .A2(new_n312), .A3(new_n725), .ZN(new_n747));
  OAI21_X1  g561(.A(KEYINPUT42), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n689), .A2(new_n568), .ZN(new_n749));
  AOI211_X1 g563(.A(new_n458), .B(new_n749), .C1(new_n464), .C2(new_n442), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n740), .A2(KEYINPUT42), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n750), .A2(new_n708), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n196), .ZN(G33));
  INV_X1    g568(.A(KEYINPUT108), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n677), .B(new_n755), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n756), .A2(new_n708), .A3(new_n750), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G134), .ZN(G36));
  OAI21_X1  g572(.A(new_n671), .B1(new_n639), .B2(new_n641), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(KEYINPUT111), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n761));
  OAI211_X1 g575(.A(new_n761), .B(new_n671), .C1(new_n639), .C2(new_n641), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT110), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT43), .B1(new_n517), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n633), .A2(new_n517), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OAI211_X1 g580(.A(new_n633), .B(new_n517), .C1(new_n763), .C2(KEYINPUT43), .ZN(new_n767));
  AOI22_X1  g581(.A1(new_n760), .A2(new_n762), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n745), .B1(new_n768), .B2(KEYINPUT44), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n760), .A2(new_n762), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n766), .A2(new_n767), .ZN(new_n771));
  AND3_X1   g585(.A1(new_n770), .A2(KEYINPUT44), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n681), .A2(new_n619), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n617), .A2(new_n306), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(G469), .B1(new_n463), .B2(KEYINPUT45), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT45), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n449), .A2(new_n778), .A3(new_n452), .ZN(new_n779));
  OAI211_X1 g593(.A(KEYINPUT46), .B(new_n776), .C1(new_n777), .C2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT109), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n408), .A2(new_n399), .A3(new_n369), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n399), .B1(new_n408), .B2(new_n369), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n783), .B1(KEYINPUT84), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n437), .B1(new_n785), .B2(new_n409), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n447), .B1(new_n786), .B2(new_n444), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n615), .B1(new_n787), .B2(new_n445), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n778), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n463), .A2(KEYINPUT45), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n789), .A2(G469), .A3(new_n790), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(KEYINPUT109), .A3(KEYINPUT46), .A4(new_n776), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n776), .B1(new_n777), .B2(new_n779), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n443), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n774), .B1(new_n793), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n773), .A2(new_n797), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  AOI21_X1  g613(.A(new_n617), .B1(new_n788), .B2(new_n778), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n775), .B1(new_n800), .B2(new_n790), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT109), .B1(new_n801), .B2(KEYINPUT46), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n780), .A2(new_n781), .ZN(new_n803));
  OAI21_X1  g617(.A(new_n796), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n619), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(KEYINPUT47), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n458), .B1(new_n793), .B2(new_n796), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT47), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NOR4_X1   g623(.A1(new_n312), .A2(new_n365), .A3(new_n740), .A4(new_n749), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n809), .A3(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G140), .ZN(G42));
  NAND4_X1  g626(.A1(new_n678), .A2(new_n312), .A3(new_n607), .A4(new_n671), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n813), .A2(new_n612), .A3(new_n620), .ZN(new_n814));
  INV_X1    g628(.A(new_n743), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n735), .ZN(new_n817));
  XOR2_X1   g631(.A(new_n675), .B(KEYINPUT116), .Z(new_n818));
  NOR2_X1   g632(.A1(new_n671), .A2(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n465), .A2(new_n817), .A3(new_n688), .A4(new_n819), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n816), .A2(KEYINPUT52), .A3(new_n705), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n705), .A2(new_n820), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n679), .A2(new_n743), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n822), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n821), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT113), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n750), .A2(new_n742), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n465), .A2(new_n312), .A3(new_n365), .A4(new_n745), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n677), .B(KEYINPUT108), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n694), .A2(new_n516), .A3(new_n675), .ZN(new_n832));
  OAI211_X1 g646(.A(new_n745), .B(new_n832), .C1(new_n653), .C2(new_n654), .ZN(new_n833));
  INV_X1    g647(.A(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n834), .A2(new_n312), .A3(new_n671), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n612), .A2(new_n835), .A3(new_n620), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n827), .B1(new_n831), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n835), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n838), .A2(new_n459), .A3(new_n467), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(new_n757), .A3(KEYINPUT113), .A4(new_n828), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n837), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n517), .A2(new_n694), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n635), .B1(new_n634), .B2(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n459), .A2(new_n467), .A3(new_n644), .A4(new_n843), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n668), .B(new_n844), .C1(new_n368), .C2(new_n609), .ZN(new_n845));
  AOI22_X1  g659(.A1(new_n717), .A2(new_n718), .B1(new_n734), .B2(new_n737), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n708), .B(new_n711), .C1(new_n636), .C2(new_n656), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n846), .A2(new_n748), .A3(new_n752), .A4(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n845), .A2(new_n848), .ZN(new_n849));
  NAND4_X1  g663(.A1(new_n826), .A2(KEYINPUT53), .A3(new_n841), .A4(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n849), .A2(new_n841), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n853), .A2(KEYINPUT117), .A3(KEYINPUT53), .A4(new_n826), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n849), .A2(new_n841), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT115), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n858), .B1(new_n814), .B2(new_n815), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n679), .A2(KEYINPUT115), .A3(new_n743), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n820), .A2(KEYINPUT52), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n859), .A2(new_n705), .A3(new_n860), .A4(new_n861), .ZN(new_n862));
  AOI22_X1  g676(.A1(new_n856), .A2(new_n857), .B1(new_n825), .B2(new_n862), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n849), .A2(new_n841), .A3(KEYINPUT114), .ZN(new_n864));
  AOI21_X1  g678(.A(KEYINPUT53), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g679(.A(KEYINPUT54), .B1(new_n855), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n826), .A2(new_n841), .A3(new_n849), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n825), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n866), .A2(new_n873), .ZN(new_n874));
  NOR3_X1   g688(.A1(new_n688), .A2(new_n643), .A3(new_n519), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n710), .A2(new_n749), .ZN(new_n876));
  AND2_X1   g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n517), .A3(new_n632), .A4(new_n631), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n673), .B1(new_n766), .B2(new_n767), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n876), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n741), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n879), .A2(new_n734), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NOR3_X1   g697(.A1(new_n691), .A2(new_n710), .A3(new_n568), .ZN(new_n884));
  AND2_X1   g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  OR2_X1    g699(.A1(new_n885), .A2(KEYINPUT50), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(KEYINPUT50), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n881), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n882), .A2(new_n749), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n807), .B(KEYINPUT47), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n709), .A2(new_n458), .A3(new_n442), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n889), .B1(new_n890), .B2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT51), .B1(new_n888), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n725), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n707), .B2(new_n311), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n879), .A2(new_n896), .A3(new_n876), .ZN(new_n897));
  XNOR2_X1  g711(.A(KEYINPUT119), .B(KEYINPUT48), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n897), .A2(KEYINPUT119), .A3(KEYINPUT48), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n883), .A2(new_n718), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n248), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(new_n634), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n902), .B1(new_n877), .B2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n900), .A2(new_n901), .A3(new_n904), .ZN(new_n905));
  NOR3_X1   g719(.A1(new_n894), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n893), .A2(KEYINPUT51), .A3(new_n888), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n907), .A2(KEYINPUT118), .ZN(new_n909));
  NAND3_X1  g723(.A1(new_n906), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n874), .A2(new_n910), .B1(G952), .B2(G953), .ZN(new_n911));
  NOR4_X1   g725(.A1(new_n765), .A2(new_n895), .A3(new_n458), .A4(new_n692), .ZN(new_n912));
  XNOR2_X1  g726(.A(new_n912), .B(KEYINPUT112), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n709), .A2(new_n442), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT49), .ZN(new_n915));
  OR4_X1    g729(.A1(new_n691), .A2(new_n913), .A3(new_n688), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n911), .A2(new_n916), .ZN(G75));
  NOR2_X1   g731(.A1(new_n248), .A2(G952), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n306), .B1(new_n869), .B2(new_n871), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT56), .B1(new_n920), .B2(G210), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n580), .A2(new_n582), .A3(new_n591), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n589), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n919), .B1(new_n921), .B2(new_n924), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n924), .B2(new_n921), .ZN(G51));
  AND3_X1   g740(.A1(new_n853), .A2(KEYINPUT53), .A3(new_n870), .ZN(new_n927));
  AOI21_X1  g741(.A(KEYINPUT53), .B1(new_n853), .B2(new_n826), .ZN(new_n928));
  OAI21_X1  g742(.A(KEYINPUT54), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n929), .A2(KEYINPUT120), .A3(new_n873), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n869), .A2(new_n871), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT120), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n931), .A2(new_n932), .A3(KEYINPUT54), .ZN(new_n933));
  XNOR2_X1  g747(.A(new_n775), .B(KEYINPUT57), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n436), .A2(new_n439), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n920), .A2(new_n790), .A3(new_n800), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n918), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND2_X1  g753(.A1(KEYINPUT58), .A2(G475), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n920), .A2(new_n650), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n650), .B1(new_n920), .B2(new_n941), .ZN(new_n943));
  NOR3_X1   g757(.A1(new_n942), .A2(new_n943), .A3(new_n918), .ZN(G60));
  XOR2_X1   g758(.A(new_n630), .B(KEYINPUT121), .Z(new_n945));
  NAND2_X1  g759(.A1(G478), .A2(G902), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT59), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n930), .A2(new_n933), .A3(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n949), .A2(new_n919), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n874), .B2(new_n947), .ZN(new_n951));
  NOR2_X1   g765(.A1(new_n950), .A2(new_n951), .ZN(G63));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT122), .ZN(new_n955));
  NAND2_X1  g769(.A1(G217), .A2(G902), .ZN(new_n956));
  XNOR2_X1  g770(.A(new_n956), .B(KEYINPUT60), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n957), .B1(new_n869), .B2(new_n871), .ZN(new_n958));
  OR2_X1    g772(.A1(new_n663), .A2(new_n664), .ZN(new_n959));
  INV_X1    g773(.A(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n919), .B1(new_n958), .B2(new_n346), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n954), .B(new_n955), .C1(new_n962), .C2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n957), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n931), .A2(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(new_n346), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n918), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n968), .A2(KEYINPUT122), .A3(new_n953), .A4(new_n961), .ZN(new_n969));
  AND2_X1   g783(.A1(new_n964), .A2(new_n969), .ZN(G66));
  NAND3_X1  g784(.A1(new_n520), .A2(G224), .A3(G953), .ZN(new_n971));
  INV_X1    g785(.A(new_n845), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n846), .A2(new_n847), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n971), .B1(new_n974), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n922), .B1(G898), .B2(new_n248), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n975), .B(new_n976), .Z(G69));
  XNOR2_X1  g791(.A(new_n259), .B(new_n488), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n979), .B1(G900), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(new_n774), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n896), .A2(new_n817), .ZN(new_n982));
  AND4_X1   g796(.A1(KEYINPUT123), .A2(new_n804), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(KEYINPUT123), .B1(new_n797), .B2(new_n982), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  AND3_X1   g799(.A1(new_n859), .A2(new_n705), .A3(new_n860), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n757), .A2(new_n748), .A3(new_n752), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n987), .B1(new_n773), .B2(new_n797), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n985), .A2(new_n811), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n980), .B1(new_n989), .B2(G953), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n701), .A2(new_n859), .A3(new_n705), .A4(new_n860), .ZN(new_n991));
  INV_X1    g805(.A(KEYINPUT62), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  AOI22_X1  g807(.A1(new_n824), .A2(new_n858), .B1(new_n621), .B2(new_n704), .ZN(new_n994));
  NAND4_X1  g808(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n701), .A4(new_n860), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n682), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n749), .B1(new_n634), .B2(new_n842), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n997), .B(new_n998), .C1(new_n367), .C2(new_n366), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n770), .A2(new_n771), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT44), .ZN(new_n1001));
  NAND2_X1  g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n768), .A2(KEYINPUT44), .ZN(new_n1003));
  NAND3_X1  g817(.A1(new_n1002), .A2(new_n745), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n804), .A2(new_n981), .ZN(new_n1005));
  OAI21_X1  g819(.A(new_n999), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1006), .B1(new_n890), .B2(new_n810), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n996), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g822(.A(KEYINPUT124), .B(new_n990), .C1(new_n1008), .C2(new_n978), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n248), .B1(G227), .B2(G900), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OR2_X1    g825(.A1(new_n1008), .A2(new_n978), .ZN(new_n1012));
  AOI21_X1  g826(.A(KEYINPUT124), .B1(new_n1012), .B2(new_n990), .ZN(new_n1013));
  XNOR2_X1  g827(.A(new_n1011), .B(new_n1013), .ZN(G72));
  INV_X1    g828(.A(KEYINPUT127), .ZN(new_n1015));
  NAND2_X1  g829(.A1(G472), .A2(G902), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT63), .Z(new_n1017));
  OAI21_X1  g831(.A(new_n1017), .B1(new_n989), .B2(new_n974), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1018), .A2(KEYINPUT126), .ZN(new_n1019));
  INV_X1    g833(.A(KEYINPUT126), .ZN(new_n1020));
  OAI211_X1 g834(.A(new_n1020), .B(new_n1017), .C1(new_n989), .C2(new_n974), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n302), .A2(new_n252), .ZN(new_n1022));
  NAND3_X1  g836(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1017), .ZN(new_n1024));
  AND2_X1   g838(.A1(new_n261), .A2(new_n272), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(new_n303), .ZN(new_n1026));
  OAI21_X1  g840(.A(new_n1026), .B1(new_n855), .B2(new_n865), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1023), .A2(new_n919), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n974), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n996), .A2(new_n1007), .A3(new_n1029), .ZN(new_n1030));
  NAND3_X1  g844(.A1(new_n1030), .A2(KEYINPUT125), .A3(new_n1017), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n274), .B1(new_n270), .B2(new_n246), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g847(.A(KEYINPUT125), .B1(new_n1030), .B2(new_n1017), .ZN(new_n1034));
  NOR2_X1   g848(.A1(new_n1033), .A2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g849(.A(new_n1015), .B1(new_n1028), .B2(new_n1035), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n856), .A2(new_n857), .ZN(new_n1037));
  NAND3_X1  g851(.A1(new_n1037), .A2(new_n864), .A3(new_n870), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n1038), .A2(new_n868), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n1039), .A2(new_n852), .A3(new_n854), .ZN(new_n1040));
  AOI21_X1  g854(.A(new_n918), .B1(new_n1040), .B2(new_n1026), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n1030), .A2(new_n1017), .ZN(new_n1042));
  INV_X1    g856(.A(KEYINPUT125), .ZN(new_n1043));
  NAND2_X1  g857(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1044), .A2(new_n1031), .A3(new_n1032), .ZN(new_n1045));
  NAND4_X1  g859(.A1(new_n1041), .A2(new_n1045), .A3(KEYINPUT127), .A4(new_n1023), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1036), .A2(new_n1046), .ZN(G57));
endmodule


