//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 0 0 0 0 0 1 0 1 0 1 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:49 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n840, new_n841,
    new_n843, new_n844, new_n846, new_n847, new_n848, new_n849, new_n850,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n908, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n952, new_n953, new_n954, new_n955, new_n957, new_n958, new_n959,
    new_n960, new_n962, new_n963;
  XNOR2_X1  g000(.A(KEYINPUT31), .B(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT3), .ZN(new_n205));
  XNOR2_X1  g004(.A(G197gat), .B(G204gat), .ZN(new_n206));
  INV_X1    g005(.A(G211gat), .ZN(new_n207));
  INV_X1    g006(.A(G218gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g008(.A(new_n206), .B1(KEYINPUT22), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(G211gat), .B(G218gat), .ZN(new_n211));
  XNOR2_X1  g010(.A(new_n210), .B(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(new_n205), .B1(new_n212), .B2(KEYINPUT29), .ZN(new_n213));
  NAND2_X1  g012(.A1(G155gat), .A2(G162gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT2), .ZN(new_n215));
  OR2_X1    g014(.A1(G141gat), .A2(G148gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(G141gat), .A2(G148gat), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n215), .A2(new_n216), .A3(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT76), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n214), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(G155gat), .B(G162gat), .ZN(new_n222));
  INV_X1    g021(.A(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n218), .A2(new_n222), .A3(new_n220), .ZN(new_n225));
  NAND3_X1  g024(.A1(new_n213), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AND3_X1   g025(.A1(new_n218), .A2(new_n222), .A3(new_n220), .ZN(new_n227));
  AOI21_X1  g026(.A(new_n222), .B1(new_n218), .B2(new_n220), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n205), .B1(new_n227), .B2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n212), .B1(new_n230), .B2(KEYINPUT29), .ZN(new_n231));
  INV_X1    g030(.A(G50gat), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n226), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n232), .B1(new_n226), .B2(new_n231), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n204), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(new_n235), .ZN(new_n237));
  INV_X1    g036(.A(new_n204), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n237), .A2(new_n233), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(G78gat), .B(G106gat), .ZN(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n236), .A2(new_n239), .A3(new_n241), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT78), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n225), .A3(KEYINPUT3), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT1), .ZN(new_n250));
  INV_X1    g049(.A(G113gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n251), .A2(G120gat), .ZN(new_n252));
  INV_X1    g051(.A(G120gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n253), .A2(G113gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n250), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G127gat), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G127gat), .A2(G134gat), .ZN(new_n259));
  AND2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT69), .B1(new_n251), .B2(G120gat), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT69), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n263), .A2(new_n253), .A3(G113gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n251), .A2(G120gat), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT1), .B1(new_n258), .B2(new_n259), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n261), .A2(new_n268), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n229), .A2(new_n249), .A3(new_n269), .ZN(new_n270));
  AOI22_X1  g069(.A1(new_n255), .A2(new_n260), .B1(new_n266), .B2(new_n267), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n271), .B(new_n272), .C1(new_n228), .C2(new_n227), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n224), .A2(new_n225), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n272), .B1(new_n275), .B2(new_n271), .ZN(new_n276));
  OAI211_X1 g075(.A(new_n248), .B(new_n270), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT5), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n269), .A2(new_n224), .A3(new_n225), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n271), .B1(new_n228), .B2(new_n227), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n248), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n277), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(KEYINPUT77), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n277), .A2(new_n283), .A3(new_n286), .ZN(new_n287));
  OR2_X1    g086(.A1(new_n277), .A2(KEYINPUT5), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n285), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  XNOR2_X1  g088(.A(G1gat), .B(G29gat), .ZN(new_n290));
  INV_X1    g089(.A(G85gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n290), .B(new_n291), .ZN(new_n292));
  XNOR2_X1  g091(.A(KEYINPUT0), .B(G57gat), .ZN(new_n293));
  XOR2_X1   g092(.A(new_n292), .B(new_n293), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n296));
  INV_X1    g095(.A(new_n294), .ZN(new_n297));
  NAND4_X1  g096(.A1(new_n285), .A2(new_n288), .A3(new_n297), .A4(new_n287), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n295), .A2(new_n296), .A3(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n289), .A2(KEYINPUT6), .A3(new_n294), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(G226gat), .A2(G233gat), .ZN(new_n302));
  INV_X1    g101(.A(new_n302), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(KEYINPUT29), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT25), .ZN(new_n305));
  AND3_X1   g104(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n307));
  NOR2_X1   g106(.A1(G183gat), .A2(G190gat), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(G169gat), .ZN(new_n310));
  INV_X1    g109(.A(G176gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n310), .A2(new_n311), .A3(KEYINPUT23), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(G169gat), .B2(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G169gat), .A2(G176gat), .ZN(new_n315));
  NAND3_X1  g114(.A1(new_n312), .A2(new_n314), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n305), .B1(new_n309), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT64), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g118(.A(KEYINPUT64), .B(new_n305), .C1(new_n309), .C2(new_n316), .ZN(new_n320));
  AND4_X1   g119(.A1(KEYINPUT25), .A2(new_n312), .A3(new_n314), .A4(new_n315), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n307), .B(KEYINPUT65), .ZN(new_n322));
  INV_X1    g121(.A(new_n306), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT66), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n324), .ZN(new_n325));
  OAI21_X1  g124(.A(KEYINPUT66), .B1(G183gat), .B2(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n323), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n321), .B1(new_n322), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n319), .A2(new_n320), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT28), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n330), .A2(G190gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  NOR2_X1   g132(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT68), .ZN(new_n335));
  NOR3_X1   g134(.A1(new_n333), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337));
  INV_X1    g136(.A(G183gat), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(KEYINPUT68), .B1(new_n339), .B2(new_n332), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n331), .B1(new_n336), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(G190gat), .B1(new_n339), .B2(new_n332), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT67), .B1(new_n342), .B2(KEYINPUT28), .ZN(new_n343));
  INV_X1    g142(.A(G190gat), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n344), .B1(new_n333), .B2(new_n334), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT67), .ZN(new_n346));
  NAND3_X1  g145(.A1(new_n345), .A2(new_n346), .A3(new_n330), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n341), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n315), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n310), .A2(new_n311), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n349), .B1(KEYINPUT26), .B2(new_n350), .ZN(new_n351));
  OR2_X1    g150(.A1(new_n350), .A2(KEYINPUT26), .ZN(new_n352));
  AOI22_X1  g151(.A1(new_n351), .A2(new_n352), .B1(G183gat), .B2(G190gat), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n348), .A2(new_n353), .ZN(new_n354));
  AND3_X1   g153(.A1(new_n329), .A2(KEYINPUT74), .A3(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT74), .B1(new_n329), .B2(new_n354), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n304), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n329), .A2(new_n354), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n359), .A2(new_n303), .ZN(new_n360));
  AND3_X1   g159(.A1(new_n357), .A2(new_n212), .A3(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT74), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n329), .A2(new_n354), .A3(KEYINPUT74), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n303), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n358), .A2(new_n304), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n212), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  XNOR2_X1  g166(.A(G8gat), .B(G36gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(G64gat), .B(G92gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n361), .A2(new_n367), .A3(new_n370), .ZN(new_n371));
  XOR2_X1   g170(.A(new_n370), .B(KEYINPUT75), .Z(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n212), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n355), .A2(new_n356), .A3(new_n302), .ZN(new_n375));
  INV_X1    g174(.A(new_n366), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n374), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n357), .A2(new_n212), .A3(new_n360), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(KEYINPUT30), .B1(new_n371), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n370), .ZN(new_n381));
  NAND3_X1  g180(.A1(new_n377), .A2(new_n378), .A3(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT30), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AND4_X1   g183(.A1(new_n247), .A2(new_n301), .A3(new_n380), .A4(new_n384), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n372), .B1(new_n361), .B2(new_n367), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n383), .B1(new_n386), .B2(new_n382), .ZN(new_n387));
  AND2_X1   g186(.A1(new_n382), .A2(new_n383), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n247), .B1(new_n389), .B2(new_n301), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n246), .B1(new_n385), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n380), .A2(new_n384), .ZN(new_n392));
  OAI21_X1  g191(.A(KEYINPUT39), .B1(new_n281), .B2(new_n282), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT79), .ZN(new_n394));
  OR2_X1    g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n393), .A2(new_n394), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n274), .A2(new_n276), .ZN(new_n397));
  AND2_X1   g196(.A1(new_n397), .A2(new_n270), .ZN(new_n398));
  OAI211_X1 g197(.A(new_n395), .B(new_n396), .C1(new_n398), .C2(new_n248), .ZN(new_n399));
  AOI21_X1  g198(.A(new_n248), .B1(new_n397), .B2(new_n270), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT39), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n294), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n399), .A2(KEYINPUT40), .A3(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n295), .ZN(new_n404));
  AOI21_X1  g203(.A(KEYINPUT40), .B1(new_n399), .B2(new_n402), .ZN(new_n405));
  NOR3_X1   g204(.A1(new_n403), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n246), .B1(new_n392), .B2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n408));
  NAND3_X1  g207(.A1(new_n377), .A2(new_n408), .A3(new_n378), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n212), .B1(new_n375), .B2(new_n376), .ZN(new_n410));
  NAND3_X1  g209(.A1(new_n357), .A2(new_n374), .A3(new_n360), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n410), .A2(KEYINPUT37), .A3(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n373), .A2(KEYINPUT38), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT80), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  NAND4_X1  g215(.A1(new_n409), .A2(new_n412), .A3(new_n416), .A4(new_n413), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  AND2_X1   g217(.A1(new_n299), .A2(new_n300), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n418), .A2(new_n419), .A3(new_n382), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT38), .ZN(new_n421));
  INV_X1    g220(.A(new_n409), .ZN(new_n422));
  OAI21_X1  g221(.A(KEYINPUT37), .B1(new_n361), .B2(new_n367), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n370), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n422), .B1(new_n424), .B2(KEYINPUT81), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT81), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n423), .A2(new_n426), .A3(new_n370), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n421), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n407), .B1(new_n420), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT71), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n358), .A2(new_n271), .ZN(new_n431));
  NAND2_X1  g230(.A1(G227gat), .A2(G233gat), .ZN(new_n432));
  AOI21_X1  g231(.A(new_n269), .B1(new_n329), .B2(new_n354), .ZN(new_n433));
  NOR3_X1   g232(.A1(new_n431), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT32), .ZN(new_n435));
  XNOR2_X1  g234(.A(G15gat), .B(G43gat), .ZN(new_n436));
  XNOR2_X1  g235(.A(G71gat), .B(G99gat), .ZN(new_n437));
  XOR2_X1   g236(.A(new_n436), .B(new_n437), .Z(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n435), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  OAI21_X1  g240(.A(new_n430), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n359), .A2(new_n269), .ZN(new_n443));
  INV_X1    g242(.A(new_n432), .ZN(new_n444));
  INV_X1    g243(.A(new_n433), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n443), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n446), .A2(KEYINPUT71), .A3(new_n440), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n442), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n439), .A2(new_n435), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n446), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n438), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n448), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT34), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n453), .B1(new_n432), .B2(KEYINPUT72), .ZN(new_n454));
  INV_X1    g253(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n443), .A2(new_n445), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n455), .B1(new_n456), .B2(new_n432), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n432), .B(new_n455), .C1(new_n431), .C2(new_n433), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n452), .A2(new_n461), .ZN(new_n462));
  AOI22_X1  g261(.A1(new_n442), .A2(new_n447), .B1(new_n450), .B2(new_n438), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n463), .A2(new_n460), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n462), .A2(KEYINPUT36), .A3(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT73), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n466), .B1(new_n463), .B2(new_n460), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n462), .A2(new_n464), .ZN(new_n468));
  AOI21_X1  g267(.A(new_n467), .B1(new_n468), .B2(new_n466), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n469), .B2(KEYINPUT36), .ZN(new_n470));
  AND3_X1   g269(.A1(new_n391), .A2(new_n429), .A3(new_n470), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n452), .A2(new_n461), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n463), .A2(new_n460), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n466), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n467), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT35), .ZN(new_n477));
  NAND4_X1  g276(.A1(new_n389), .A2(new_n477), .A3(new_n301), .A4(new_n245), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  OAI21_X1  g278(.A(KEYINPUT78), .B1(new_n419), .B2(new_n392), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n389), .A2(new_n247), .A3(new_n301), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n468), .A2(new_n246), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n480), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n479), .B1(KEYINPUT35), .B2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT82), .B1(new_n471), .B2(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G134gat), .B(G162gat), .Z(new_n486));
  AND2_X1   g285(.A1(G232gat), .A2(G233gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n487), .A2(KEYINPUT41), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n486), .B(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G43gat), .B(G50gat), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n490), .A2(KEYINPUT83), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT83), .ZN(new_n492));
  INV_X1    g291(.A(G43gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(G50gat), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n232), .A2(G43gat), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n492), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g295(.A1(new_n491), .A2(new_n496), .A3(KEYINPUT15), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT14), .ZN(new_n498));
  INV_X1    g297(.A(G29gat), .ZN(new_n499));
  INV_X1    g298(.A(G36gat), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n502));
  AOI22_X1  g301(.A1(new_n501), .A2(new_n502), .B1(G29gat), .B2(G36gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(KEYINPUT84), .B(KEYINPUT15), .ZN(new_n504));
  OAI21_X1  g303(.A(new_n503), .B1(new_n490), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT85), .B1(new_n497), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n491), .A2(new_n496), .A3(KEYINPUT15), .ZN(new_n507));
  OR2_X1    g306(.A1(new_n507), .A2(new_n503), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT85), .ZN(new_n509));
  OR2_X1    g308(.A1(new_n490), .A2(new_n504), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n507), .A2(new_n509), .A3(new_n510), .A4(new_n503), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n506), .A2(new_n508), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT17), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT17), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n506), .A2(new_n508), .A3(new_n514), .A4(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G99gat), .B(G106gat), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  NOR2_X1   g317(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g318(.A1(G85gat), .A2(G92gat), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(G92gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n291), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(G99gat), .A2(G106gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n524), .A2(KEYINPUT8), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n521), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(KEYINPUT91), .A2(KEYINPUT7), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n528), .A2(new_n519), .A3(new_n520), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n518), .B1(new_n526), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT91), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT7), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND4_X1  g332(.A1(new_n533), .A2(G85gat), .A3(G92gat), .A4(new_n527), .ZN(new_n534));
  AOI22_X1  g333(.A1(KEYINPUT8), .A2(new_n524), .B1(new_n291), .B2(new_n522), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n534), .A2(new_n517), .A3(new_n521), .A4(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n530), .A2(KEYINPUT92), .A3(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT92), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n538), .B(new_n518), .C1(new_n526), .C2(new_n529), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT94), .ZN(new_n543));
  NAND3_X1  g342(.A1(new_n537), .A2(KEYINPUT93), .A3(new_n539), .ZN(new_n544));
  AND3_X1   g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  AOI21_X1  g344(.A(new_n543), .B1(new_n542), .B2(new_n544), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n516), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n547), .A2(KEYINPUT95), .ZN(new_n548));
  XOR2_X1   g347(.A(G190gat), .B(G218gat), .Z(new_n549));
  INV_X1    g348(.A(KEYINPUT95), .ZN(new_n550));
  OAI211_X1 g349(.A(new_n516), .B(new_n550), .C1(new_n545), .C2(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n487), .A2(KEYINPUT41), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n542), .A2(new_n544), .ZN(new_n553));
  INV_X1    g352(.A(new_n512), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n548), .A2(new_n549), .A3(new_n551), .A4(new_n556), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT96), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n555), .B1(new_n547), .B2(KEYINPUT95), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT96), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n559), .A2(new_n560), .A3(new_n549), .A4(new_n551), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n558), .A2(new_n561), .A3(KEYINPUT97), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n549), .B1(new_n559), .B2(new_n551), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(KEYINPUT97), .B1(new_n558), .B2(new_n561), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n489), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n558), .A2(new_n561), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n489), .B1(new_n563), .B2(KEYINPUT98), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n568), .B(new_n569), .C1(KEYINPUT98), .C2(new_n563), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n567), .A2(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(G8gat), .ZN(new_n572));
  XNOR2_X1  g371(.A(G15gat), .B(G22gat), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT16), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(G1gat), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n575), .B2(KEYINPUT86), .ZN(new_n576));
  OAI21_X1  g375(.A(new_n575), .B1(G1gat), .B2(new_n573), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n576), .B(new_n577), .ZN(new_n578));
  OR2_X1    g377(.A1(G57gat), .A2(G64gat), .ZN(new_n579));
  NAND2_X1  g378(.A1(G57gat), .A2(G64gat), .ZN(new_n580));
  NAND2_X1  g379(.A1(G71gat), .A2(G78gat), .ZN(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  OAI211_X1 g381(.A(new_n579), .B(new_n580), .C1(new_n582), .C2(KEYINPUT9), .ZN(new_n583));
  NAND2_X1  g382(.A1(KEYINPUT89), .A2(KEYINPUT9), .ZN(new_n584));
  OR2_X1    g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n583), .A2(new_n581), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  OR2_X1    g385(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n585), .A2(new_n581), .A3(new_n584), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n587), .A2(new_n579), .A3(new_n580), .A4(new_n588), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n586), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n578), .B1(KEYINPUT21), .B2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n591), .B(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(G127gat), .B(G155gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n594), .B(KEYINPUT20), .Z(new_n595));
  XNOR2_X1  g394(.A(new_n593), .B(new_n595), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n590), .A2(KEYINPUT21), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(new_n338), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n599), .B(new_n207), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n597), .B(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  OR2_X1    g401(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n596), .A2(new_n602), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT99), .B1(new_n571), .B2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT99), .ZN(new_n608));
  NAND4_X1  g407(.A1(new_n567), .A2(new_n608), .A3(new_n570), .A4(new_n605), .ZN(new_n609));
  AND2_X1   g408(.A1(new_n607), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n483), .A2(KEYINPUT35), .ZN(new_n611));
  INV_X1    g410(.A(new_n479), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT82), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n391), .A2(new_n429), .A3(new_n470), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n578), .B1(new_n513), .B2(new_n515), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n512), .A2(new_n578), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G229gat), .A2(G233gat), .ZN(new_n620));
  XOR2_X1   g419(.A(new_n620), .B(KEYINPUT87), .Z(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT18), .B1(new_n619), .B2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT18), .ZN(new_n624));
  NOR4_X1   g423(.A1(new_n617), .A2(new_n618), .A3(new_n624), .A4(new_n621), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n512), .A2(new_n578), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n618), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g426(.A(KEYINPUT88), .B(KEYINPUT13), .Z(new_n628));
  XNOR2_X1  g427(.A(new_n621), .B(new_n628), .ZN(new_n629));
  NOR2_X1   g428(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n623), .A2(new_n625), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G113gat), .B(G141gat), .ZN(new_n632));
  INV_X1    g431(.A(G197gat), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT11), .B(G169gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT12), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n631), .B(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT100), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n590), .A2(new_n640), .A3(new_n530), .A4(new_n536), .ZN(new_n641));
  NAND4_X1  g440(.A1(new_n530), .A2(new_n586), .A3(new_n589), .A4(new_n536), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT100), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n586), .A2(new_n589), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n537), .A2(new_n644), .A3(new_n539), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n641), .A2(new_n643), .A3(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(G230gat), .A2(G233gat), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n649), .B(KEYINPUT101), .Z(new_n650));
  NAND4_X1  g449(.A1(new_n542), .A2(KEYINPUT10), .A3(new_n544), .A4(new_n590), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT10), .ZN(new_n652));
  NAND4_X1  g451(.A1(new_n641), .A2(new_n643), .A3(new_n645), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n647), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n650), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n657), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n650), .A2(new_n661), .A3(new_n655), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n639), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n485), .A2(new_n610), .A3(new_n616), .A4(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT102), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n666), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n419), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n670), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  NAND3_X1  g471(.A1(new_n669), .A2(new_n392), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n572), .B1(new_n669), .B2(new_n392), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT42), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n673), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n673), .ZN(new_n677));
  AOI21_X1  g476(.A(KEYINPUT103), .B1(new_n677), .B2(KEYINPUT42), .ZN(new_n678));
  INV_X1    g477(.A(KEYINPUT103), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n673), .A2(new_n679), .A3(new_n675), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n676), .B1(new_n678), .B2(new_n680), .ZN(G1325gat));
  NOR2_X1   g480(.A1(new_n476), .A2(G15gat), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n669), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(G15gat), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n470), .B1(new_n667), .B2(new_n668), .ZN(new_n685));
  OAI21_X1  g484(.A(new_n683), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT104), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n686), .B(new_n687), .ZN(G1326gat));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT105), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n690), .B1(new_n669), .B2(new_n246), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  AOI211_X1 g491(.A(KEYINPUT105), .B(new_n245), .C1(new_n667), .C2(new_n668), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n689), .B1(new_n692), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n689), .ZN(new_n696));
  NOR3_X1   g495(.A1(new_n691), .A2(new_n693), .A3(new_n696), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n695), .A2(new_n697), .ZN(G1327gat));
  AND2_X1   g497(.A1(new_n567), .A2(new_n570), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n605), .ZN(new_n700));
  NAND4_X1  g499(.A1(new_n485), .A2(new_n616), .A3(new_n664), .A4(new_n700), .ZN(new_n701));
  NOR3_X1   g500(.A1(new_n701), .A2(G29gat), .A3(new_n301), .ZN(new_n702));
  XOR2_X1   g501(.A(new_n702), .B(KEYINPUT45), .Z(new_n703));
  NAND3_X1  g502(.A1(new_n485), .A2(new_n571), .A3(new_n616), .ZN(new_n704));
  OAI21_X1  g503(.A(KEYINPUT107), .B1(new_n471), .B2(new_n484), .ZN(new_n705));
  INV_X1    g504(.A(KEYINPUT107), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n613), .A2(new_n706), .A3(new_n615), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n705), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n699), .A2(KEYINPUT44), .ZN(new_n709));
  AOI22_X1  g508(.A1(new_n704), .A2(KEYINPUT44), .B1(new_n708), .B2(new_n709), .ZN(new_n710));
  XNOR2_X1  g509(.A(new_n663), .B(KEYINPUT106), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n712), .A2(new_n639), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n710), .A2(new_n605), .A3(new_n714), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n715), .A2(new_n419), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n703), .B1(new_n716), .B2(new_n499), .ZN(G1328gat));
  NOR3_X1   g516(.A1(new_n701), .A2(G36gat), .A3(new_n389), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT46), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n715), .A2(new_n392), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n719), .B1(new_n720), .B2(new_n500), .ZN(G1329gat));
  NAND2_X1  g520(.A1(new_n469), .A2(new_n493), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n701), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(new_n723), .ZN(new_n724));
  NOR4_X1   g523(.A1(new_n710), .A2(new_n605), .A3(new_n470), .A4(new_n714), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n725), .B2(new_n493), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT108), .ZN(new_n727));
  AOI21_X1  g526(.A(KEYINPUT47), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n704), .A2(KEYINPUT44), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n708), .A2(new_n709), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n470), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n731), .A2(new_n606), .A3(new_n732), .A4(new_n713), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n723), .B1(new_n733), .B2(G43gat), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n734), .A2(KEYINPUT108), .A3(new_n735), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n728), .A2(new_n736), .ZN(G1330gat));
  NOR3_X1   g536(.A1(new_n701), .A2(G50gat), .A3(new_n245), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT48), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n731), .A2(new_n606), .A3(new_n246), .A4(new_n713), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G50gat), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n741), .A2(KEYINPUT109), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n740), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n232), .B1(new_n715), .B2(new_n246), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n739), .B1(new_n746), .B2(new_n738), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n745), .A2(new_n747), .ZN(G1331gat));
  AND4_X1   g547(.A1(new_n610), .A2(new_n708), .A3(new_n639), .A4(new_n712), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n419), .ZN(new_n750));
  XOR2_X1   g549(.A(KEYINPUT110), .B(G57gat), .Z(new_n751));
  XNOR2_X1  g550(.A(new_n750), .B(new_n751), .ZN(G1332gat));
  NAND2_X1  g551(.A1(new_n749), .A2(new_n392), .ZN(new_n753));
  OAI21_X1  g552(.A(new_n753), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(KEYINPUT49), .B(G64gat), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n749), .A2(new_n392), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT111), .ZN(new_n758));
  XNOR2_X1  g557(.A(new_n757), .B(new_n758), .ZN(G1333gat));
  NAND2_X1  g558(.A1(new_n749), .A2(new_n732), .ZN(new_n760));
  NOR2_X1   g559(.A1(new_n476), .A2(G71gat), .ZN(new_n761));
  AOI22_X1  g560(.A1(new_n760), .A2(G71gat), .B1(new_n749), .B2(new_n761), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g562(.A1(new_n749), .A2(new_n246), .ZN(new_n764));
  XNOR2_X1  g563(.A(KEYINPUT112), .B(G78gat), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n764), .B(new_n765), .ZN(G1335gat));
  OAI211_X1 g565(.A(new_n639), .B(new_n700), .C1(new_n471), .C2(new_n484), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT51), .ZN(new_n768));
  INV_X1    g567(.A(new_n663), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n770), .A2(new_n291), .A3(new_n419), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n639), .A2(new_n663), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n710), .A2(new_n605), .A3(new_n772), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n773), .A2(new_n419), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n771), .B1(new_n774), .B2(new_n291), .ZN(G1336gat));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n768), .A2(new_n711), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n777), .A2(new_n522), .A3(new_n392), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n773), .A2(new_n392), .ZN(new_n779));
  OAI211_X1 g578(.A(new_n776), .B(new_n778), .C1(new_n779), .C2(new_n522), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n522), .B1(new_n773), .B2(new_n392), .ZN(new_n781));
  INV_X1    g580(.A(new_n778), .ZN(new_n782));
  OAI21_X1  g581(.A(KEYINPUT52), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n780), .A2(new_n783), .ZN(G1337gat));
  INV_X1    g583(.A(G99gat), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n770), .A2(new_n785), .A3(new_n469), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n773), .A2(new_n732), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n786), .B1(new_n787), .B2(new_n785), .ZN(G1338gat));
  NOR2_X1   g587(.A1(new_n245), .A2(G106gat), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n777), .A2(new_n789), .ZN(new_n790));
  AND2_X1   g589(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(G106gat), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n773), .A2(new_n246), .ZN(new_n794));
  OAI211_X1 g593(.A(new_n791), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n793), .B1(new_n773), .B2(new_n246), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n790), .A2(KEYINPUT113), .ZN(new_n797));
  OAI21_X1  g596(.A(KEYINPUT53), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(G1339gat));
  INV_X1    g598(.A(KEYINPUT116), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n800), .B1(new_n619), .B2(new_n622), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n627), .A2(new_n629), .ZN(new_n802));
  OAI211_X1 g601(.A(KEYINPUT116), .B(new_n621), .C1(new_n617), .C2(new_n618), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n801), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n631), .A2(new_n637), .B1(new_n804), .B2(new_n636), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n663), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n651), .A2(new_n648), .A3(new_n653), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n655), .A2(KEYINPUT114), .A3(KEYINPUT54), .A4(new_n807), .ZN(new_n808));
  AND3_X1   g607(.A1(new_n651), .A2(new_n648), .A3(new_n653), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT54), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n648), .B1(new_n651), .B2(new_n653), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n810), .A2(KEYINPUT114), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n809), .A2(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n808), .A2(new_n813), .A3(KEYINPUT55), .A4(new_n659), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(new_n662), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT115), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n814), .A2(KEYINPUT115), .A3(new_n662), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n808), .A2(new_n813), .A3(new_n659), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT55), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n817), .A2(new_n818), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n806), .B1(new_n639), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n699), .A2(new_n823), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n817), .A2(new_n805), .A3(new_n818), .A4(new_n821), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n825), .B1(new_n567), .B2(new_n570), .ZN(new_n826));
  INV_X1    g625(.A(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n828), .A2(new_n606), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n638), .A2(new_n663), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n607), .A2(new_n609), .A3(new_n830), .ZN(new_n831));
  AOI211_X1 g630(.A(new_n246), .B(new_n468), .C1(new_n829), .C2(new_n831), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n392), .A2(new_n301), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n834), .A2(new_n251), .A3(new_n638), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n246), .B1(new_n829), .B2(new_n831), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n469), .A3(new_n833), .ZN(new_n837));
  OAI21_X1  g636(.A(G113gat), .B1(new_n837), .B2(new_n639), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n835), .A2(new_n838), .ZN(G1340gat));
  NAND3_X1  g638(.A1(new_n834), .A2(new_n253), .A3(new_n663), .ZN(new_n840));
  OAI21_X1  g639(.A(G120gat), .B1(new_n837), .B2(new_n711), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1341gat));
  NOR3_X1   g641(.A1(new_n837), .A2(new_n256), .A3(new_n606), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n834), .A2(new_n605), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n843), .B1(new_n844), .B2(new_n256), .ZN(G1342gat));
  AOI21_X1  g644(.A(new_n301), .B1(new_n829), .B2(new_n831), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n699), .A2(new_n392), .ZN(new_n847));
  NAND4_X1  g646(.A1(new_n846), .A2(new_n257), .A3(new_n482), .A4(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(new_n848), .B(KEYINPUT56), .Z(new_n849));
  OAI21_X1  g648(.A(G134gat), .B1(new_n837), .B2(new_n699), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(G1343gat));
  INV_X1    g650(.A(KEYINPUT57), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT55), .B1(new_n819), .B2(KEYINPUT117), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT117), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n808), .A2(new_n813), .A3(new_n855), .A4(new_n659), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n815), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n638), .B1(new_n857), .B2(KEYINPUT118), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n819), .A2(KEYINPUT117), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(new_n820), .A3(new_n856), .ZN(new_n860));
  INV_X1    g659(.A(new_n815), .ZN(new_n861));
  AND3_X1   g660(.A1(new_n860), .A2(KEYINPUT118), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n806), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n826), .B1(new_n863), .B2(new_n699), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n853), .B1(new_n864), .B2(new_n605), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n860), .A2(new_n861), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n857), .A2(KEYINPUT118), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n638), .A3(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n571), .B1(new_n870), .B2(new_n806), .ZN(new_n871));
  OAI211_X1 g670(.A(KEYINPUT119), .B(new_n606), .C1(new_n871), .C2(new_n826), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n865), .A2(new_n831), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n852), .B1(new_n873), .B2(new_n246), .ZN(new_n874));
  AND3_X1   g673(.A1(new_n607), .A2(new_n609), .A3(new_n830), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n605), .B1(new_n824), .B2(new_n827), .ZN(new_n876));
  OAI211_X1 g675(.A(new_n852), .B(new_n246), .C1(new_n875), .C2(new_n876), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n470), .A2(new_n833), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n874), .A2(new_n879), .A3(new_n639), .ZN(new_n880));
  INV_X1    g679(.A(G141gat), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT120), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n732), .A2(new_n245), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n846), .A2(new_n883), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n885), .A2(new_n881), .A3(new_n389), .A4(new_n638), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n886), .B1(new_n880), .B2(new_n881), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT58), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n882), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI221_X1 g688(.A(new_n886), .B1(KEYINPUT120), .B2(KEYINPUT58), .C1(new_n880), .C2(new_n881), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(G1344gat));
  INV_X1    g690(.A(KEYINPUT59), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n884), .A2(new_n392), .ZN(new_n893));
  AOI211_X1 g692(.A(new_n892), .B(G148gat), .C1(new_n893), .C2(new_n663), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n874), .A2(new_n879), .A3(new_n769), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n831), .B1(new_n605), .B2(new_n864), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n896), .A2(new_n852), .A3(new_n246), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n245), .B1(new_n829), .B2(new_n831), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n898), .B2(new_n852), .ZN(new_n899));
  XOR2_X1   g698(.A(new_n878), .B(KEYINPUT121), .Z(new_n900));
  OR3_X1    g699(.A1(new_n900), .A2(new_n892), .A3(new_n769), .ZN(new_n901));
  OAI22_X1  g700(.A1(new_n895), .A2(KEYINPUT59), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n894), .B1(new_n902), .B2(G148gat), .ZN(G1345gat));
  AOI21_X1  g702(.A(G155gat), .B1(new_n893), .B2(new_n605), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n874), .A2(new_n879), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n605), .A2(G155gat), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n904), .B1(new_n905), .B2(new_n906), .ZN(G1346gat));
  INV_X1    g706(.A(G162gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n885), .A2(new_n908), .A3(new_n847), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n874), .A2(new_n879), .A3(new_n699), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n908), .ZN(G1347gat));
  NOR2_X1   g710(.A1(new_n419), .A2(new_n389), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n832), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n913), .A2(new_n310), .A3(new_n638), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n469), .A2(new_n912), .ZN(new_n915));
  XOR2_X1   g714(.A(new_n915), .B(KEYINPUT122), .Z(new_n916));
  NAND2_X1  g715(.A1(new_n836), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT123), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n836), .A2(KEYINPUT123), .A3(new_n916), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n921), .A2(new_n638), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n914), .B1(new_n922), .B2(new_n310), .ZN(G1348gat));
  AOI21_X1  g722(.A(G176gat), .B1(new_n913), .B2(new_n663), .ZN(new_n924));
  NOR2_X1   g723(.A1(new_n711), .A2(new_n311), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n924), .B1(new_n921), .B2(new_n925), .ZN(G1349gat));
  NAND3_X1  g725(.A1(new_n919), .A2(new_n605), .A3(new_n920), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G183gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n336), .A2(new_n340), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n606), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g729(.A(KEYINPUT124), .B1(new_n913), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  XNOR2_X1  g731(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n928), .A2(new_n931), .A3(new_n933), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1350gat));
  NAND3_X1  g736(.A1(new_n919), .A2(new_n571), .A3(new_n920), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n938), .A2(G190gat), .ZN(new_n939));
  XNOR2_X1  g738(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n940));
  OR2_X1    g739(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n939), .A2(new_n940), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n913), .A2(new_n344), .A3(new_n571), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(G1351gat));
  NAND2_X1  g743(.A1(new_n470), .A2(new_n912), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n899), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g746(.A(G197gat), .B1(new_n947), .B2(new_n639), .ZN(new_n948));
  AOI211_X1 g747(.A(new_n245), .B(new_n945), .C1(new_n829), .C2(new_n831), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n949), .A2(new_n633), .A3(new_n638), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1352gat));
  INV_X1    g750(.A(G204gat), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n949), .A2(new_n952), .A3(new_n663), .ZN(new_n953));
  XOR2_X1   g752(.A(new_n953), .B(KEYINPUT62), .Z(new_n954));
  OAI21_X1  g753(.A(G204gat), .B1(new_n947), .B2(new_n711), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n954), .A2(new_n955), .ZN(G1353gat));
  NAND3_X1  g755(.A1(new_n949), .A2(new_n207), .A3(new_n605), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n946), .A2(new_n605), .ZN(new_n958));
  AND3_X1   g757(.A1(new_n958), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n959));
  AOI21_X1  g758(.A(KEYINPUT63), .B1(new_n958), .B2(G211gat), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n959), .B2(new_n960), .ZN(G1354gat));
  AOI21_X1  g760(.A(G218gat), .B1(new_n949), .B2(new_n571), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n699), .A2(new_n208), .ZN(new_n963));
  AOI21_X1  g762(.A(new_n962), .B1(new_n946), .B2(new_n963), .ZN(G1355gat));
endmodule


