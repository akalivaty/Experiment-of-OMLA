//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 0 0 1 0 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 0 0 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 0 0 1 1 1 0 1 0 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:43 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(G110), .B(G140), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(G227), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT77), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT11), .ZN(new_n196));
  INV_X1    g010(.A(G134), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n196), .B1(new_n197), .B2(G137), .ZN(new_n198));
  INV_X1    g012(.A(G137), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(KEYINPUT11), .A3(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n197), .A2(G137), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G131), .ZN(new_n203));
  INV_X1    g017(.A(G131), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n200), .A3(new_n204), .A4(new_n201), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT3), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(KEYINPUT3), .A3(G104), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n209), .A2(new_n211), .ZN(new_n212));
  XNOR2_X1  g026(.A(KEYINPUT79), .B(G101), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT78), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n214), .B1(new_n210), .B2(G104), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n208), .A2(KEYINPUT78), .A3(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n212), .A2(new_n213), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  OAI21_X1  g031(.A(KEYINPUT81), .B1(new_n210), .B2(G104), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT81), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n208), .A3(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n210), .A2(G104), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  XNOR2_X1  g037(.A(G143), .B(G146), .ZN(new_n224));
  INV_X1    g038(.A(G128), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  AOI21_X1  g041(.A(new_n226), .B1(G143), .B2(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n225), .B1(new_n228), .B2(KEYINPUT82), .ZN(new_n229));
  INV_X1    g043(.A(G143), .ZN(new_n230));
  OAI21_X1  g044(.A(KEYINPUT1), .B1(new_n230), .B2(G146), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT82), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n224), .B1(new_n229), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n227), .A2(G143), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n230), .A2(G146), .ZN(new_n236));
  NAND4_X1  g050(.A1(new_n235), .A2(new_n236), .A3(new_n226), .A4(G128), .ZN(new_n237));
  INV_X1    g051(.A(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n217), .B(new_n223), .C1(new_n234), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n217), .A2(new_n223), .ZN(new_n240));
  AOI22_X1  g054(.A1(new_n231), .A2(G128), .B1(new_n235), .B2(new_n236), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  AOI21_X1  g057(.A(new_n206), .B1(new_n239), .B2(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n203), .A2(new_n205), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT12), .B1(new_n245), .B2(KEYINPUT83), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n244), .B(new_n247), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT10), .ZN(new_n249));
  INV_X1    g063(.A(new_n240), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n242), .A2(new_n249), .ZN(new_n251));
  AOI22_X1  g065(.A1(new_n239), .A2(new_n249), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n217), .A2(KEYINPUT4), .ZN(new_n253));
  INV_X1    g067(.A(G101), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n215), .A2(new_n216), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n254), .B1(new_n255), .B2(new_n212), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n212), .A2(new_n215), .A3(new_n216), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT4), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n258), .A2(new_n259), .A3(G101), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n235), .A2(new_n236), .A3(KEYINPUT0), .A4(G128), .ZN(new_n261));
  XNOR2_X1  g075(.A(KEYINPUT0), .B(G128), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n224), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n260), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT80), .ZN(new_n266));
  NOR3_X1   g080(.A1(new_n257), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n263), .B1(new_n256), .B2(new_n259), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n258), .A2(G101), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n269), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT80), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n252), .B(new_n206), .C1(new_n267), .C2(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n195), .B1(new_n248), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n272), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT84), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n235), .A2(KEYINPUT82), .A3(KEYINPUT1), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n233), .A2(G128), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n235), .A2(new_n236), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n238), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n249), .B1(new_n279), .B2(new_n240), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n225), .B1(new_n235), .B2(KEYINPUT1), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n237), .B1(new_n281), .B2(new_n224), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n282), .A2(new_n217), .A3(new_n223), .A4(KEYINPUT10), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n280), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(new_n266), .B1(new_n257), .B2(new_n265), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n268), .A2(new_n270), .A3(KEYINPUT80), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n284), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n275), .B1(new_n287), .B2(new_n206), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n252), .B1(new_n267), .B2(new_n271), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT84), .A3(new_n245), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n274), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n273), .B1(new_n291), .B2(new_n193), .ZN(new_n292));
  OAI21_X1  g106(.A(G469), .B1(new_n292), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(G469), .ZN(new_n294));
  INV_X1    g108(.A(G902), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n288), .A2(new_n290), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n193), .B1(new_n296), .B2(new_n272), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n272), .A2(new_n193), .ZN(new_n298));
  XNOR2_X1  g112(.A(new_n244), .B(new_n246), .ZN(new_n299));
  OAI21_X1  g113(.A(KEYINPUT85), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT85), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n248), .A2(new_n301), .A3(new_n272), .A4(new_n193), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n294), .B(new_n295), .C1(new_n297), .C2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n189), .B1(new_n293), .B2(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(G478), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n306), .A2(KEYINPUT15), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n308), .A2(G128), .A3(new_n230), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n230), .A2(G128), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n225), .A2(G143), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI211_X1 g126(.A(new_n309), .B(G134), .C1(new_n312), .C2(new_n308), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n310), .A2(new_n311), .A3(new_n197), .ZN(new_n314));
  XNOR2_X1  g128(.A(G116), .B(G122), .ZN(new_n315));
  XNOR2_X1  g129(.A(new_n315), .B(new_n210), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n313), .A2(new_n314), .A3(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(G217), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n187), .A2(new_n318), .A3(G953), .ZN(new_n319));
  INV_X1    g133(.A(G122), .ZN(new_n320));
  OAI21_X1  g134(.A(KEYINPUT14), .B1(new_n320), .B2(G116), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT93), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g137(.A(G116), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G122), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n325), .A2(KEYINPUT93), .A3(KEYINPUT14), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n320), .A2(G116), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT14), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n328), .A2(new_n324), .A3(G122), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n323), .A2(new_n326), .A3(new_n327), .A4(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G107), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(G134), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n332), .A2(new_n314), .B1(new_n210), .B2(new_n315), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n331), .A2(KEYINPUT94), .A3(new_n333), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT94), .B1(new_n331), .B2(new_n333), .ZN(new_n335));
  OAI211_X1 g149(.A(new_n317), .B(new_n319), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT95), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n317), .B1(new_n334), .B2(new_n335), .ZN(new_n339));
  INV_X1    g153(.A(new_n319), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT94), .ZN(new_n342));
  AOI21_X1  g156(.A(KEYINPUT93), .B1(new_n325), .B2(KEYINPUT14), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n329), .A2(new_n327), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n210), .B1(new_n345), .B2(new_n326), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n315), .A2(new_n210), .ZN(new_n347));
  INV_X1    g161(.A(new_n314), .ZN(new_n348));
  AOI21_X1  g162(.A(new_n197), .B1(new_n310), .B2(new_n311), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n347), .B1(new_n348), .B2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n342), .B1(new_n346), .B2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n331), .A2(KEYINPUT94), .A3(new_n333), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(KEYINPUT95), .A3(new_n317), .A4(new_n319), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n338), .A2(new_n341), .A3(new_n354), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(KEYINPUT96), .A3(new_n295), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(KEYINPUT96), .B1(new_n355), .B2(new_n295), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n307), .B1(new_n357), .B2(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n358), .A2(new_n307), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  XNOR2_X1  g176(.A(G113), .B(G122), .ZN(new_n363));
  XNOR2_X1  g177(.A(new_n363), .B(new_n208), .ZN(new_n364));
  INV_X1    g178(.A(G237), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n191), .A3(G214), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n230), .ZN(new_n367));
  NOR2_X1   g181(.A1(G237), .A2(G953), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n368), .A2(G143), .A3(G214), .ZN(new_n369));
  NAND2_X1  g183(.A1(KEYINPUT18), .A2(G131), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n367), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G140), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G125), .ZN(new_n373));
  INV_X1    g187(.A(G125), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G140), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n373), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n376), .A2(G146), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n373), .A2(new_n375), .A3(new_n227), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n367), .A2(new_n369), .ZN(new_n380));
  INV_X1    g194(.A(new_n370), .ZN(new_n381));
  AOI21_X1  g195(.A(KEYINPUT91), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT91), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n383), .B(new_n370), .C1(new_n367), .C2(new_n369), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n371), .B(new_n379), .C1(new_n382), .C2(new_n384), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n368), .A2(G143), .A3(G214), .ZN(new_n386));
  AOI21_X1  g200(.A(G143), .B1(new_n368), .B2(G214), .ZN(new_n387));
  OAI21_X1  g201(.A(G131), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n367), .A2(new_n204), .A3(new_n369), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT16), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n372), .A3(G125), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT72), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT16), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n391), .A2(new_n372), .A3(KEYINPUT72), .A4(G125), .ZN(new_n396));
  NAND4_X1  g210(.A1(new_n394), .A2(new_n395), .A3(G146), .A4(new_n396), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n373), .A2(new_n375), .A3(KEYINPUT19), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT19), .B1(new_n373), .B2(new_n375), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n227), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n390), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n364), .B1(new_n385), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n379), .A2(new_n371), .ZN(new_n403));
  NOR2_X1   g217(.A1(new_n386), .A2(new_n387), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n383), .B1(new_n404), .B2(new_n370), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n380), .A2(KEYINPUT91), .A3(new_n381), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n403), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n227), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT73), .A3(new_n397), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT73), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n411), .A3(new_n227), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT17), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n388), .A2(new_n414), .A3(new_n389), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n380), .A2(KEYINPUT17), .A3(G131), .ZN(new_n416));
  AND2_X1   g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n407), .B1(new_n413), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n402), .B1(new_n418), .B2(new_n364), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT20), .B1(new_n419), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT20), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n415), .A2(new_n416), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n412), .B2(new_n410), .ZN(new_n425));
  INV_X1    g239(.A(new_n364), .ZN(new_n426));
  NOR3_X1   g240(.A1(new_n425), .A2(new_n426), .A3(new_n407), .ZN(new_n427));
  OAI211_X1 g241(.A(new_n423), .B(new_n420), .C1(new_n427), .C2(new_n402), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n422), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n413), .A2(new_n417), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n364), .B1(new_n430), .B2(new_n385), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n295), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G475), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n362), .A2(new_n434), .ZN(new_n435));
  AND2_X1   g249(.A1(new_n191), .A2(G952), .ZN(new_n436));
  NAND2_X1  g250(.A1(G234), .A2(G237), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(G898), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n437), .A2(G902), .A3(G953), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G214), .B1(G237), .B2(G902), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n242), .A2(new_n374), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n263), .A2(G125), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AND2_X1   g260(.A1(new_n191), .A2(G224), .ZN(new_n447));
  XNOR2_X1  g261(.A(new_n446), .B(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT86), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(G119), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n324), .A2(G119), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(KEYINPUT5), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n453), .A2(KEYINPUT5), .ZN(new_n458));
  INV_X1    g272(.A(G113), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(KEYINPUT2), .B(G113), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  AOI22_X1  g276(.A1(new_n457), .A2(new_n460), .B1(new_n456), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n250), .A2(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n455), .B(new_n461), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n465), .B(new_n260), .C1(new_n253), .C2(new_n256), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n451), .B1(new_n464), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT6), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n464), .A2(new_n466), .A3(new_n451), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n468), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT87), .B1(new_n467), .B2(new_n468), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n448), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n450), .B(KEYINPUT88), .ZN(new_n477));
  OR2_X1    g291(.A1(new_n477), .A2(KEYINPUT8), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(KEYINPUT8), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n464), .A2(KEYINPUT89), .ZN(new_n480));
  OR2_X1    g294(.A1(new_n250), .A2(new_n463), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n464), .A2(KEYINPUT89), .ZN(new_n483));
  OAI211_X1 g297(.A(new_n478), .B(new_n479), .C1(new_n482), .C2(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT7), .ZN(new_n485));
  OR2_X1    g299(.A1(new_n485), .A2(KEYINPUT90), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n444), .A2(new_n445), .A3(new_n486), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n485), .B2(new_n447), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n447), .A2(new_n485), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n444), .A2(new_n445), .A3(new_n489), .A4(new_n486), .ZN(new_n490));
  AND3_X1   g304(.A1(new_n488), .A2(new_n470), .A3(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(G902), .B1(new_n484), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(G210), .B1(G237), .B2(G902), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n476), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n476), .B2(new_n492), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n442), .B(new_n443), .C1(new_n494), .C2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  AND3_X1   g311(.A1(new_n305), .A2(new_n435), .A3(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT70), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n225), .B2(G119), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n452), .A2(KEYINPUT70), .A3(G128), .ZN(new_n501));
  AOI22_X1  g315(.A1(new_n500), .A2(new_n501), .B1(G119), .B2(new_n225), .ZN(new_n502));
  XOR2_X1   g316(.A(KEYINPUT24), .B(G110), .Z(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n225), .A2(G119), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n452), .A2(G128), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT71), .A4(KEYINPUT23), .ZN(new_n507));
  OR2_X1    g321(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT71), .A2(KEYINPUT23), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n508), .A2(G119), .A3(new_n225), .A4(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n510), .A3(G110), .ZN(new_n511));
  AND2_X1   g325(.A1(new_n504), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n410), .A2(new_n412), .A3(new_n512), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n502), .A2(new_n503), .ZN(new_n514));
  AOI21_X1  g328(.A(G110), .B1(new_n507), .B2(new_n510), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n378), .B(new_n397), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT22), .B(G137), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n517), .B(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n516), .A3(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n520), .A2(new_n295), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n513), .A2(new_n516), .ZN(new_n522));
  INV_X1    g336(.A(new_n519), .ZN(new_n523));
  AOI21_X1  g337(.A(KEYINPUT74), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT74), .ZN(new_n525));
  AOI211_X1 g339(.A(new_n525), .B(new_n519), .C1(new_n513), .C2(new_n516), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n521), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT25), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n529));
  OAI211_X1 g343(.A(new_n521), .B(new_n529), .C1(new_n524), .C2(new_n526), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n318), .B1(G234), .B2(new_n295), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n528), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(KEYINPUT75), .ZN(new_n533));
  INV_X1    g347(.A(new_n531), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n527), .B2(KEYINPUT25), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT75), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n536), .A3(new_n530), .ZN(new_n537));
  OR2_X1    g351(.A1(new_n524), .A2(new_n526), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n531), .A2(G902), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n520), .A3(new_n539), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n533), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n264), .A2(new_n245), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n199), .A2(G134), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n204), .B1(new_n544), .B2(new_n201), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(KEYINPUT65), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT65), .ZN(new_n547));
  AOI211_X1 g361(.A(new_n547), .B(new_n204), .C1(new_n544), .C2(new_n201), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n282), .B(new_n205), .C1(new_n546), .C2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n543), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n465), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n368), .A2(G210), .ZN(new_n553));
  XNOR2_X1  g367(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(KEYINPUT26), .B(G101), .ZN(new_n555));
  AND2_X1   g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n555), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT29), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n556), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT28), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n278), .B1(new_n228), .B2(new_n225), .ZN(new_n561));
  AND3_X1   g375(.A1(new_n198), .A2(new_n200), .A3(new_n201), .ZN(new_n562));
  AOI22_X1  g376(.A1(new_n237), .A2(new_n561), .B1(new_n562), .B2(new_n204), .ZN(new_n563));
  XNOR2_X1  g377(.A(new_n545), .B(KEYINPUT65), .ZN(new_n564));
  AOI22_X1  g378(.A1(new_n563), .A2(new_n564), .B1(new_n245), .B2(new_n264), .ZN(new_n565));
  INV_X1    g379(.A(new_n465), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n560), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n543), .A2(new_n549), .A3(new_n566), .A4(new_n560), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n551), .B(new_n559), .C1(new_n567), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT69), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n543), .A2(new_n549), .A3(new_n566), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(KEYINPUT28), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n568), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT69), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n574), .A2(new_n575), .A3(new_n551), .A4(new_n559), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n571), .A2(new_n295), .A3(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT64), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n264), .A2(new_n245), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n579), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n578), .B1(new_n264), .B2(new_n245), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n549), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n582), .A2(new_n465), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n556), .A2(new_n557), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n583), .A2(new_n574), .A3(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT68), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n583), .A2(new_n574), .A3(KEYINPUT68), .A4(new_n584), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n587), .A2(new_n558), .A3(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n565), .A2(KEYINPUT30), .ZN(new_n590));
  INV_X1    g404(.A(new_n549), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n543), .A2(KEYINPUT64), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(new_n579), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n465), .B(new_n590), .C1(new_n593), .C2(KEYINPUT30), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n584), .B1(new_n594), .B2(new_n572), .ZN(new_n595));
  OAI21_X1  g409(.A(new_n577), .B1(new_n589), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n596), .A2(G472), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n584), .B1(new_n583), .B2(new_n574), .ZN(new_n598));
  AND2_X1   g412(.A1(new_n584), .A2(new_n572), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT31), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n594), .A2(KEYINPUT31), .A3(new_n599), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n598), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g418(.A1(G472), .A2(G902), .ZN(new_n605));
  XNOR2_X1  g419(.A(new_n605), .B(KEYINPUT67), .ZN(new_n606));
  NOR3_X1   g420(.A1(new_n604), .A2(KEYINPUT32), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT32), .ZN(new_n608));
  AND3_X1   g422(.A1(new_n594), .A2(KEYINPUT31), .A3(new_n599), .ZN(new_n609));
  AOI21_X1  g423(.A(KEYINPUT31), .B1(new_n594), .B2(new_n599), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n583), .A2(new_n574), .ZN(new_n611));
  OAI22_X1  g425(.A1(new_n609), .A2(new_n610), .B1(new_n611), .B2(new_n584), .ZN(new_n612));
  INV_X1    g426(.A(new_n606), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n608), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n597), .B1(new_n607), .B2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT76), .B1(new_n542), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(KEYINPUT32), .B1(new_n604), .B2(new_n606), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n612), .A2(new_n608), .A3(new_n613), .ZN(new_n618));
  AOI22_X1  g432(.A1(new_n617), .A2(new_n618), .B1(new_n596), .B2(G472), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT76), .ZN(new_n620));
  NOR3_X1   g434(.A1(new_n619), .A2(new_n620), .A3(new_n541), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n498), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  XOR2_X1   g436(.A(new_n622), .B(new_n213), .Z(G3));
  INV_X1    g437(.A(G472), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n624), .B1(new_n612), .B2(new_n295), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT97), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n625), .A2(new_n626), .B1(new_n606), .B2(new_n604), .ZN(new_n627));
  AOI211_X1 g441(.A(KEYINPUT97), .B(new_n624), .C1(new_n612), .C2(new_n295), .ZN(new_n628));
  NOR3_X1   g442(.A1(new_n627), .A2(new_n541), .A3(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT99), .ZN(new_n630));
  AND2_X1   g444(.A1(new_n429), .A2(new_n433), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n341), .A2(KEYINPUT33), .A3(new_n336), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n306), .A2(G902), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT98), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT33), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n355), .A2(new_n634), .A3(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n634), .B1(new_n355), .B2(new_n635), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n632), .B(new_n633), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n355), .A2(new_n295), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n639), .A2(new_n306), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n631), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n630), .B1(new_n497), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n638), .A2(new_n640), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n434), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n644), .A2(new_n496), .A3(KEYINPUT99), .ZN(new_n645));
  OAI211_X1 g459(.A(new_n305), .B(new_n629), .C1(new_n642), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT34), .B(G104), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G6));
  NAND2_X1  g462(.A1(new_n293), .A2(new_n304), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n497), .A2(new_n649), .A3(new_n188), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n650), .A2(new_n629), .A3(new_n362), .A4(new_n631), .ZN(new_n651));
  XOR2_X1   g465(.A(KEYINPUT35), .B(G107), .Z(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G9));
  NOR2_X1   g467(.A1(new_n627), .A2(new_n628), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n523), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n522), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n539), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n533), .A2(new_n537), .A3(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n533), .A2(KEYINPUT100), .A3(new_n537), .A4(new_n657), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n650), .A2(new_n654), .A3(new_n662), .A4(new_n435), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT37), .B(G110), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G12));
  AND4_X1   g479(.A1(new_n536), .A2(new_n528), .A3(new_n530), .A4(new_n531), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n536), .B1(new_n535), .B2(new_n530), .ZN(new_n667));
  NOR2_X1   g481(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(KEYINPUT100), .B1(new_n668), .B2(new_n657), .ZN(new_n669));
  INV_X1    g483(.A(new_n661), .ZN(new_n670));
  OAI211_X1 g484(.A(new_n305), .B(new_n615), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n438), .B1(G900), .B2(new_n441), .ZN(new_n672));
  AND3_X1   g486(.A1(new_n429), .A2(new_n433), .A3(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n307), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT96), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n639), .A2(new_n675), .ZN(new_n676));
  AOI21_X1  g490(.A(new_n674), .B1(new_n676), .B2(new_n356), .ZN(new_n677));
  OAI21_X1  g491(.A(new_n673), .B1(new_n677), .B2(new_n360), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT101), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n443), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n476), .A2(new_n492), .ZN(new_n682));
  INV_X1    g496(.A(new_n493), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n476), .A2(new_n492), .A3(new_n493), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n681), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g500(.A(new_n673), .B(KEYINPUT101), .C1(new_n677), .C2(new_n360), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n680), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT102), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT102), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n680), .A2(new_n690), .A3(new_n686), .A4(new_n687), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n671), .B1(new_n689), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n225), .ZN(G30));
  INV_X1    g507(.A(new_n594), .ZN(new_n694));
  INV_X1    g508(.A(new_n572), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n584), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n584), .ZN(new_n697));
  AOI21_X1  g511(.A(G902), .B1(new_n697), .B2(new_n551), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n624), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n617), .B2(new_n618), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT103), .ZN(new_n701));
  OR2_X1    g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n700), .A2(new_n701), .ZN(new_n703));
  AND2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n684), .A2(new_n685), .ZN(new_n706));
  XOR2_X1   g520(.A(new_n706), .B(KEYINPUT38), .Z(new_n707));
  NOR2_X1   g521(.A1(new_n631), .A2(new_n681), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n708), .A2(new_n362), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n707), .A2(new_n662), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n672), .B(KEYINPUT39), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n305), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n713));
  OR2_X1    g527(.A1(new_n712), .A2(KEYINPUT40), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n705), .A2(new_n710), .A3(new_n713), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G143), .ZN(G45));
  AND3_X1   g530(.A1(new_n641), .A2(new_n686), .A3(new_n672), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n662), .A2(new_n717), .A3(new_n305), .A4(new_n615), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  NOR2_X1   g533(.A1(new_n619), .A2(new_n541), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n295), .B1(new_n297), .B2(new_n303), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n721), .A2(G469), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n722), .A2(new_n188), .A3(new_n304), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  OAI211_X1 g538(.A(new_n720), .B(new_n724), .C1(new_n642), .C2(new_n645), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT41), .B(G113), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G15));
  AND3_X1   g541(.A1(new_n497), .A2(new_n362), .A3(new_n631), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n720), .A3(new_n724), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G116), .ZN(G18));
  NAND2_X1  g544(.A1(new_n497), .A2(new_n435), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n731), .A2(new_n723), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n619), .B1(new_n660), .B2(new_n661), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n732), .A2(KEYINPUT104), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(KEYINPUT104), .B1(new_n732), .B2(new_n733), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(new_n452), .ZN(G21));
  NAND4_X1  g551(.A1(new_n722), .A2(new_n188), .A3(new_n304), .A4(new_n442), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n708), .A2(new_n362), .A3(new_n706), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(new_n625), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n609), .A2(new_n610), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n584), .B1(new_n574), .B2(new_n551), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n613), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n741), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n745), .A2(new_n541), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n740), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G122), .ZN(G24));
  AOI21_X1  g562(.A(new_n745), .B1(new_n660), .B2(new_n661), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n641), .A2(new_n672), .ZN(new_n750));
  INV_X1    g564(.A(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n722), .A2(new_n686), .A3(new_n188), .A4(new_n304), .ZN(new_n752));
  INV_X1    g566(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(new_n751), .A3(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G125), .ZN(G27));
  NOR2_X1   g569(.A1(new_n706), .A2(new_n681), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n305), .A2(new_n542), .A3(new_n615), .A4(new_n756), .ZN(new_n757));
  OAI21_X1  g571(.A(KEYINPUT105), .B1(new_n757), .B2(new_n750), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT42), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(KEYINPUT105), .B(KEYINPUT42), .C1(new_n757), .C2(new_n750), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n762), .B(new_n204), .ZN(G33));
  INV_X1    g577(.A(new_n757), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n680), .A2(new_n687), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(KEYINPUT107), .ZN(new_n768));
  NAND2_X1  g582(.A1(G469), .A2(G902), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n291), .A2(new_n193), .ZN(new_n770));
  INV_X1    g584(.A(new_n273), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT45), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n294), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT106), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n292), .A2(KEYINPUT45), .ZN(new_n776));
  AND3_X1   g590(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n775), .B1(new_n774), .B2(new_n776), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n769), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT46), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n768), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n774), .A2(new_n776), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT106), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n774), .A2(new_n775), .A3(new_n776), .ZN(new_n784));
  NAND2_X1  g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n785), .A2(KEYINPUT107), .A3(KEYINPUT46), .A4(new_n769), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n779), .A2(new_n780), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n781), .A2(new_n304), .A3(new_n786), .A4(new_n787), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(new_n188), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n434), .B1(new_n638), .B2(new_n640), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(KEYINPUT43), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n791), .B(new_n662), .C1(new_n628), .C2(new_n627), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT44), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n756), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n792), .B2(new_n793), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n789), .A2(new_n711), .A3(new_n794), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(G137), .ZN(G39));
  XOR2_X1   g612(.A(KEYINPUT108), .B(KEYINPUT47), .Z(new_n799));
  AND3_X1   g613(.A1(new_n788), .A2(new_n188), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT47), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n788), .A2(new_n188), .B1(KEYINPUT108), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  NOR4_X1   g617(.A1(new_n795), .A2(new_n750), .A3(new_n542), .A4(new_n615), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  NOR2_X1   g620(.A1(new_n700), .A2(new_n658), .ZN(new_n807));
  INV_X1    g621(.A(new_n739), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n808), .A3(new_n305), .A4(new_n672), .ZN(new_n809));
  AND2_X1   g623(.A1(new_n718), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n689), .A2(new_n691), .ZN(new_n811));
  AND3_X1   g625(.A1(new_n662), .A2(new_n305), .A3(new_n615), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n810), .A2(new_n813), .A3(new_n754), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT52), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n810), .A2(new_n813), .A3(KEYINPUT52), .A4(new_n754), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n542), .A2(new_n615), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n819), .A2(new_n723), .ZN(new_n820));
  AOI22_X1  g634(.A1(new_n820), .A2(new_n728), .B1(new_n740), .B2(new_n746), .ZN(new_n821));
  OAI211_X1 g635(.A(new_n821), .B(new_n725), .C1(new_n734), .C2(new_n735), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n644), .A2(KEYINPUT109), .ZN(new_n823));
  OAI21_X1  g637(.A(KEYINPUT110), .B1(new_n677), .B2(new_n360), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n359), .A2(new_n361), .A3(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n824), .A2(new_n826), .A3(new_n631), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT109), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n641), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n823), .A2(new_n827), .A3(new_n829), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n650), .A3(new_n629), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT111), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n622), .A2(new_n663), .A3(new_n831), .A4(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n622), .A2(new_n663), .A3(new_n831), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n834), .A2(KEYINPUT111), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n822), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n824), .A2(new_n826), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n615), .A3(new_n673), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n838), .B1(new_n750), .B2(new_n745), .ZN(new_n839));
  INV_X1    g653(.A(new_n305), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n840), .A2(new_n795), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n839), .A2(new_n662), .A3(new_n841), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n761), .A2(new_n760), .A3(new_n766), .A4(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n818), .A2(new_n836), .A3(KEYINPUT53), .A4(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n835), .A2(new_n833), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n725), .A2(new_n729), .A3(new_n747), .ZN(new_n847));
  INV_X1    g661(.A(new_n734), .ZN(new_n848));
  INV_X1    g662(.A(new_n735), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n846), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT115), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT53), .A4(new_n818), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n845), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n846), .A2(new_n843), .A3(new_n850), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n856));
  XNOR2_X1  g670(.A(KEYINPUT114), .B(KEYINPUT52), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n814), .A2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT113), .ZN(new_n859));
  INV_X1    g673(.A(new_n754), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n859), .B1(new_n692), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n813), .A2(KEYINPUT113), .A3(new_n754), .ZN(new_n862));
  AND3_X1   g676(.A1(new_n718), .A2(new_n809), .A3(KEYINPUT52), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n855), .A2(new_n856), .B1(new_n858), .B2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n836), .A2(KEYINPUT112), .A3(new_n843), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT53), .B1(new_n865), .B2(new_n866), .ZN(new_n867));
  OAI21_X1  g681(.A(KEYINPUT54), .B1(new_n854), .B2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT53), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n816), .A2(new_n817), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n855), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT54), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n864), .A2(new_n858), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n873), .A2(KEYINPUT53), .A3(new_n836), .A4(new_n843), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n868), .A2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(new_n438), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n791), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n724), .A2(new_n756), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  AND2_X1   g694(.A1(new_n880), .A2(KEYINPUT118), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n880), .A2(KEYINPUT118), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n749), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT50), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n443), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n707), .A2(new_n724), .A3(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n791), .A2(new_n877), .A3(new_n746), .ZN(new_n888));
  NOR2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n884), .A2(new_n885), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n879), .A2(new_n438), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n643), .A2(new_n434), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n542), .A3(new_n704), .A4(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT119), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n883), .B(new_n891), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n722), .A2(new_n304), .ZN(new_n899));
  OAI22_X1  g713(.A1(new_n800), .A2(new_n802), .B1(new_n188), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n888), .A2(new_n795), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(KEYINPUT116), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n903), .A2(KEYINPUT51), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n903), .A2(KEYINPUT51), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n705), .A2(new_n541), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n906), .A2(new_n641), .A3(new_n892), .ZN(new_n907));
  OAI211_X1 g721(.A(new_n907), .B(new_n436), .C1(new_n752), .C2(new_n888), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n881), .A2(new_n882), .ZN(new_n909));
  OR3_X1    g723(.A1(new_n909), .A2(KEYINPUT48), .A3(new_n819), .ZN(new_n910));
  OAI21_X1  g724(.A(KEYINPUT48), .B1(new_n909), .B2(new_n819), .ZN(new_n911));
  AOI21_X1  g725(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n904), .A2(new_n905), .A3(new_n912), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n876), .A2(new_n913), .B1(G952), .B2(G953), .ZN(new_n914));
  AND4_X1   g728(.A1(new_n188), .A2(new_n707), .A3(new_n443), .A4(new_n790), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n899), .B(KEYINPUT49), .Z(new_n916));
  NAND3_X1  g730(.A1(new_n906), .A2(new_n915), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n914), .A2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n191), .A2(G952), .ZN(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n295), .B1(new_n871), .B2(new_n874), .ZN(new_n921));
  AOI21_X1  g735(.A(KEYINPUT56), .B1(new_n921), .B2(G210), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT120), .Z(new_n924));
  XOR2_X1   g738(.A(new_n448), .B(KEYINPUT55), .Z(new_n925));
  XNOR2_X1  g739(.A(new_n924), .B(new_n925), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n920), .B1(new_n922), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n927), .B1(new_n922), .B2(new_n926), .ZN(G51));
  AND3_X1   g742(.A1(new_n871), .A2(new_n872), .A3(new_n874), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n872), .B1(new_n871), .B2(new_n874), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n769), .B(KEYINPUT57), .ZN(new_n932));
  OAI22_X1  g746(.A1(new_n931), .A2(new_n932), .B1(new_n297), .B2(new_n303), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n921), .A2(new_n784), .A3(new_n783), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n919), .B1(new_n933), .B2(new_n934), .ZN(G54));
  NAND3_X1  g749(.A1(new_n921), .A2(KEYINPUT58), .A3(G475), .ZN(new_n936));
  AND2_X1   g750(.A1(new_n936), .A2(new_n419), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n419), .ZN(new_n938));
  NOR3_X1   g752(.A1(new_n937), .A2(new_n938), .A3(new_n919), .ZN(G60));
  INV_X1    g753(.A(KEYINPUT122), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n632), .B1(new_n636), .B2(new_n637), .ZN(new_n941));
  XNOR2_X1  g755(.A(new_n941), .B(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(G478), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT59), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n942), .A2(new_n944), .ZN(new_n945));
  AOI21_X1  g759(.A(KEYINPUT53), .B1(new_n851), .B2(new_n818), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n864), .A2(new_n858), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n846), .A2(new_n843), .A3(new_n850), .A4(KEYINPUT53), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT54), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n945), .B1(new_n950), .B2(new_n875), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n940), .B1(new_n951), .B2(new_n919), .ZN(new_n952));
  INV_X1    g766(.A(new_n945), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n953), .B1(new_n929), .B2(new_n930), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n954), .A2(KEYINPUT122), .A3(new_n920), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n952), .A2(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n942), .B1(new_n876), .B2(new_n944), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G63));
  XNOR2_X1  g772(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n318), .A2(new_n295), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n959), .B(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n961), .B1(new_n946), .B2(new_n949), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n538), .A2(new_n520), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n919), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g778(.A(new_n961), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n965), .B1(new_n871), .B2(new_n874), .ZN(new_n966));
  AND3_X1   g780(.A1(new_n966), .A2(KEYINPUT124), .A3(new_n656), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT124), .B1(new_n966), .B2(new_n656), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT125), .ZN(new_n970));
  AOI21_X1  g784(.A(KEYINPUT61), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI221_X1 g786(.A(new_n964), .B1(new_n970), .B2(KEYINPUT61), .C1(new_n967), .C2(new_n968), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n972), .A2(new_n973), .ZN(G66));
  AOI21_X1  g788(.A(new_n191), .B1(new_n440), .B2(G224), .ZN(new_n975));
  INV_X1    g789(.A(new_n836), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n975), .B1(new_n976), .B2(new_n191), .ZN(new_n977));
  INV_X1    g791(.A(G898), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n924), .B1(new_n978), .B2(G953), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n977), .B(new_n979), .ZN(G69));
  INV_X1    g794(.A(G227), .ZN(new_n981));
  INV_X1    g795(.A(G900), .ZN(new_n982));
  MUX2_X1   g796(.A(new_n593), .B(new_n550), .S(KEYINPUT30), .Z(new_n983));
  OR2_X1    g797(.A1(new_n398), .A2(new_n399), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI221_X1 g800(.A(G953), .B1(new_n981), .B2(new_n982), .C1(new_n986), .C2(KEYINPUT127), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n861), .A2(new_n862), .ZN(new_n989));
  AND2_X1   g803(.A1(new_n989), .A2(new_n718), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT62), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n990), .A2(new_n991), .A3(new_n715), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n989), .A2(new_n715), .A3(new_n718), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n992), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n712), .A2(new_n795), .ZN(new_n996));
  OAI211_X1 g810(.A(new_n996), .B(new_n830), .C1(new_n616), .C2(new_n621), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n805), .A2(new_n797), .A3(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n995), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n985), .B1(new_n1000), .B2(new_n191), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n986), .B1(G900), .B2(G953), .ZN(new_n1002));
  INV_X1    g816(.A(new_n1002), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n762), .B1(new_n765), .B2(new_n764), .ZN(new_n1004));
  NAND4_X1  g818(.A1(new_n805), .A2(new_n797), .A3(new_n1004), .A4(new_n990), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n819), .A2(new_n739), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n789), .A2(new_n711), .A3(new_n1006), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT126), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NOR2_X1   g823(.A1(new_n1005), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n1003), .B1(new_n1010), .B2(new_n191), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n988), .B1(new_n1001), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1007), .B(KEYINPUT126), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n990), .A2(new_n1004), .ZN(new_n1014));
  NAND4_X1  g828(.A1(new_n1013), .A2(new_n797), .A3(new_n805), .A4(new_n1014), .ZN(new_n1015));
  OAI21_X1  g829(.A(new_n1002), .B1(new_n1015), .B2(G953), .ZN(new_n1016));
  AOI21_X1  g830(.A(G953), .B1(new_n995), .B2(new_n999), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n1016), .B(new_n987), .C1(new_n1017), .C2(new_n985), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1012), .A2(new_n1018), .ZN(G72));
  NAND2_X1  g833(.A1(new_n594), .A2(new_n697), .ZN(new_n1020));
  NOR3_X1   g834(.A1(new_n1005), .A2(new_n1009), .A3(new_n1020), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n992), .A2(new_n994), .ZN(new_n1022));
  NOR3_X1   g836(.A1(new_n1022), .A2(new_n998), .A3(new_n696), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n836), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n696), .A2(new_n1020), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XNOR2_X1  g840(.A(new_n1026), .B(KEYINPUT63), .ZN(new_n1027));
  NOR2_X1   g841(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1028), .B1(new_n854), .B2(new_n867), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n919), .B1(new_n1025), .B2(new_n1027), .ZN(new_n1030));
  AND3_X1   g844(.A1(new_n1024), .A2(new_n1029), .A3(new_n1030), .ZN(G57));
endmodule


