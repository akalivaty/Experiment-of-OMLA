//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 0 0 0 1 1 0 0 0 1 0 0 0 1 0 0 1 1 1 0 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1 0 0 1 1 0 1 1 1 0 0 1 1 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:05 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n544, new_n545,
    new_n546, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n571, new_n572, new_n573, new_n574, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G2106), .ZN(new_n455));
  INV_X1    g030(.A(G567), .ZN(new_n456));
  OAI22_X1  g031(.A1(new_n451), .A2(new_n455), .B1(new_n456), .B2(new_n452), .ZN(new_n457));
  XNOR2_X1  g032(.A(new_n457), .B(KEYINPUT65), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  NOR2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  OAI21_X1  g036(.A(KEYINPUT66), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT66), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n462), .A2(new_n468), .A3(G125), .ZN(new_n469));
  NAND2_X1  g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  AOI21_X1  g045(.A(new_n459), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(G2105), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(G101), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n474));
  INV_X1    g049(.A(G137), .ZN(new_n475));
  OAI21_X1  g050(.A(new_n473), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n471), .A2(new_n476), .ZN(G160));
  AOI21_X1  g052(.A(G2105), .B1(new_n465), .B2(new_n467), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n459), .B1(new_n465), .B2(new_n467), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  OAI211_X1 g060(.A(G126), .B(G2105), .C1(new_n460), .C2(new_n461), .ZN(new_n486));
  OR2_X1    g061(.A1(G102), .A2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(G114), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n487), .A2(new_n489), .A3(G2104), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  NOR3_X1   g067(.A1(new_n492), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n462), .A2(new_n468), .A3(new_n493), .ZN(new_n494));
  OAI211_X1 g069(.A(G138), .B(new_n459), .C1(new_n460), .C2(new_n461), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n491), .B1(new_n494), .B2(new_n496), .ZN(G164));
  INV_X1    g072(.A(G543), .ZN(new_n498));
  OAI21_X1  g073(.A(KEYINPUT68), .B1(new_n498), .B2(KEYINPUT5), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT5), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n500), .A2(new_n501), .A3(G543), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n499), .A2(new_n502), .B1(KEYINPUT5), .B2(new_n498), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT67), .B1(new_n504), .B2(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT67), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n506), .A2(new_n507), .A3(G651), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n505), .A2(new_n508), .B1(KEYINPUT6), .B2(new_n504), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI22_X1  g089(.A1(new_n503), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n515), .A2(new_n504), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n514), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n519), .B(KEYINPUT70), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  AND2_X1   g096(.A1(new_n503), .A2(new_n509), .ZN(new_n522));
  NAND2_X1  g097(.A1(new_n522), .A2(G89), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n509), .A2(G543), .ZN(new_n524));
  XOR2_X1   g099(.A(KEYINPUT69), .B(G51), .Z(new_n525));
  NAND2_X1  g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND3_X1  g101(.A1(new_n503), .A2(G63), .A3(G651), .ZN(new_n527));
  NAND4_X1  g102(.A1(new_n521), .A2(new_n523), .A3(new_n526), .A4(new_n527), .ZN(G286));
  INV_X1    g103(.A(G286), .ZN(G168));
  XOR2_X1   g104(.A(KEYINPUT71), .B(G90), .Z(new_n530));
  NAND2_X1  g105(.A1(new_n522), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n524), .A2(G52), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AOI22_X1  g108(.A1(new_n503), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n504), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n533), .A2(new_n535), .ZN(G171));
  NAND2_X1  g111(.A1(new_n522), .A2(G81), .ZN(new_n537));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n503), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n539));
  OAI221_X1 g114(.A(new_n537), .B1(new_n538), .B2(new_n512), .C1(new_n504), .C2(new_n539), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT72), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G860), .ZN(G153));
  NAND4_X1  g117(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g118(.A1(G1), .A2(G3), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT8), .ZN(new_n545));
  NAND4_X1  g120(.A1(G319), .A2(G483), .A3(G661), .A4(new_n545), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT73), .ZN(G188));
  INV_X1    g122(.A(KEYINPUT74), .ZN(new_n548));
  AOI22_X1  g123(.A1(new_n503), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n549));
  OAI21_X1  g124(.A(new_n548), .B1(new_n549), .B2(new_n504), .ZN(new_n550));
  NAND2_X1  g125(.A1(G78), .A2(G543), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n498), .A2(KEYINPUT5), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n500), .B1(new_n501), .B2(G543), .ZN(new_n553));
  NOR3_X1   g128(.A1(new_n498), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  INV_X1    g130(.A(G65), .ZN(new_n556));
  OAI21_X1  g131(.A(new_n551), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n557), .A2(KEYINPUT74), .A3(G651), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n550), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(G53), .ZN(new_n560));
  OAI21_X1  g135(.A(KEYINPUT9), .B1(new_n512), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(KEYINPUT9), .ZN(new_n562));
  NAND4_X1  g137(.A1(new_n509), .A2(new_n562), .A3(G53), .A4(G543), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n561), .A2(new_n563), .B1(G91), .B2(new_n522), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n559), .A2(new_n564), .ZN(G299));
  OAI21_X1  g140(.A(KEYINPUT75), .B1(new_n533), .B2(new_n535), .ZN(new_n566));
  INV_X1    g141(.A(new_n535), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  NAND4_X1  g143(.A1(new_n567), .A2(new_n568), .A3(new_n532), .A4(new_n531), .ZN(new_n569));
  AND2_X1   g144(.A1(new_n566), .A2(new_n569), .ZN(G301));
  NAND2_X1  g145(.A1(new_n522), .A2(G87), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n524), .A2(G49), .ZN(new_n572));
  OAI21_X1  g147(.A(G651), .B1(new_n503), .B2(G74), .ZN(new_n573));
  AND3_X1   g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G288));
  AOI22_X1  g150(.A1(new_n503), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n576));
  OAI21_X1  g151(.A(KEYINPUT76), .B1(new_n576), .B2(new_n504), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n503), .A2(new_n509), .A3(G86), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n509), .A2(G48), .A3(G543), .ZN(new_n579));
  AND2_X1   g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(G73), .A2(G543), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n555), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n583), .A2(new_n584), .A3(G651), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n577), .A2(new_n580), .A3(new_n585), .ZN(G305));
  INV_X1    g161(.A(G85), .ZN(new_n587));
  XOR2_X1   g162(.A(KEYINPUT77), .B(G47), .Z(new_n588));
  OAI22_X1  g163(.A1(new_n510), .A2(new_n587), .B1(new_n512), .B2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n503), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n590), .A2(new_n504), .ZN(new_n591));
  OR2_X1    g166(.A1(new_n589), .A2(new_n591), .ZN(G290));
  NAND2_X1  g167(.A1(new_n522), .A2(G92), .ZN(new_n593));
  INV_X1    g168(.A(KEYINPUT10), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g170(.A1(G79), .A2(G543), .ZN(new_n596));
  INV_X1    g171(.A(G66), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n555), .B2(new_n597), .ZN(new_n598));
  AOI22_X1  g173(.A1(new_n598), .A2(G651), .B1(new_n524), .B2(G54), .ZN(new_n599));
  NAND2_X1  g174(.A1(new_n595), .A2(new_n599), .ZN(new_n600));
  MUX2_X1   g175(.A(new_n600), .B(G301), .S(G868), .Z(G284));
  MUX2_X1   g176(.A(new_n600), .B(G301), .S(G868), .Z(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  INV_X1    g178(.A(G299), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G280));
  INV_X1    g181(.A(new_n600), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n541), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g188(.A1(new_n462), .A2(new_n468), .A3(new_n472), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n615), .B(KEYINPUT13), .ZN(new_n616));
  XOR2_X1   g191(.A(KEYINPUT78), .B(G2100), .Z(new_n617));
  OR2_X1    g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n616), .A2(new_n617), .ZN(new_n619));
  OAI21_X1  g194(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n620));
  INV_X1    g195(.A(KEYINPUT79), .ZN(new_n621));
  INV_X1    g196(.A(G111), .ZN(new_n622));
  AOI22_X1  g197(.A1(new_n620), .A2(new_n621), .B1(new_n622), .B2(G2105), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(new_n621), .B2(new_n620), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n478), .A2(G135), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n480), .A2(G123), .ZN(new_n626));
  AND3_X1   g201(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2096), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n618), .A2(new_n619), .A3(new_n628), .ZN(G156));
  XNOR2_X1  g204(.A(G2427), .B(G2438), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(KEYINPUT15), .B(G2435), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n633), .A2(KEYINPUT14), .A3(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT80), .B(KEYINPUT16), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G2451), .B(G2454), .Z(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n637), .B(new_n640), .ZN(new_n641));
  XOR2_X1   g216(.A(G1341), .B(G1348), .Z(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(KEYINPUT81), .ZN(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n641), .B2(new_n642), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2072), .B(G2078), .Z(new_n647));
  XOR2_X1   g222(.A(G2084), .B(G2090), .Z(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g225(.A(new_n647), .B1(new_n650), .B2(KEYINPUT18), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT82), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n652), .B(G2100), .ZN(new_n653));
  INV_X1    g228(.A(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n650), .A2(KEYINPUT17), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n648), .A2(new_n649), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(G2096), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n653), .B(new_n658), .ZN(G227));
  XNOR2_X1  g234(.A(G1971), .B(G1976), .ZN(new_n660));
  INV_X1    g235(.A(KEYINPUT19), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  AND2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(KEYINPUT83), .B(KEYINPUT20), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n663), .A2(new_n664), .ZN(new_n669));
  NOR2_X1   g244(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  MUX2_X1   g245(.A(new_n670), .B(new_n669), .S(new_n662), .Z(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  XOR2_X1   g249(.A(G1991), .B(G1996), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1981), .B(G1986), .ZN(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n676), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G229));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n681), .A2(G22), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n682), .B(KEYINPUT86), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n681), .ZN(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(G1971), .ZN(new_n685));
  OR2_X1    g260(.A1(G6), .A2(G16), .ZN(new_n686));
  OAI21_X1  g261(.A(new_n686), .B1(G305), .B2(new_n681), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT32), .B(G1981), .ZN(new_n688));
  INV_X1    g263(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n685), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n681), .A2(G23), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(new_n574), .B2(new_n681), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT33), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(G1976), .ZN(new_n694));
  OAI211_X1 g269(.A(new_n690), .B(new_n694), .C1(new_n687), .C2(new_n689), .ZN(new_n695));
  OR2_X1    g270(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n696));
  NAND2_X1  g271(.A1(new_n695), .A2(KEYINPUT34), .ZN(new_n697));
  INV_X1    g272(.A(G29), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n698), .A2(G25), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n478), .A2(G131), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n480), .A2(G119), .ZN(new_n701));
  OR2_X1    g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n700), .A2(new_n701), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n699), .B1(new_n705), .B2(new_n698), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT35), .B(G1991), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n681), .A2(G24), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT84), .Z(new_n710));
  INV_X1    g285(.A(G290), .ZN(new_n711));
  OAI21_X1  g286(.A(new_n710), .B1(new_n711), .B2(new_n681), .ZN(new_n712));
  XOR2_X1   g287(.A(KEYINPUT85), .B(G1986), .Z(new_n713));
  OAI21_X1  g288(.A(new_n708), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  AOI21_X1  g289(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n696), .A2(new_n697), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT36), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n681), .A2(G20), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT23), .Z(new_n719));
  AOI21_X1  g294(.A(new_n719), .B1(G299), .B2(G16), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT95), .Z(new_n721));
  INV_X1    g296(.A(G1956), .ZN(new_n722));
  OR2_X1    g297(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n698), .A2(G35), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n724), .B1(G162), .B2(new_n698), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT29), .Z(new_n726));
  INV_X1    g301(.A(G2090), .ZN(new_n727));
  OR2_X1    g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n721), .A2(new_n722), .ZN(new_n729));
  NAND3_X1  g304(.A1(new_n723), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT96), .ZN(new_n731));
  NOR2_X1   g306(.A1(G171), .A2(new_n681), .ZN(new_n732));
  AOI21_X1  g307(.A(new_n732), .B1(G5), .B2(new_n681), .ZN(new_n733));
  INV_X1    g308(.A(G1961), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n698), .A2(G26), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(KEYINPUT28), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n478), .A2(G140), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n480), .A2(G128), .ZN(new_n738));
  OR2_X1    g313(.A1(G104), .A2(G2105), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n739), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n740));
  NAND3_X1  g315(.A1(new_n737), .A2(new_n738), .A3(new_n740), .ZN(new_n741));
  AND3_X1   g316(.A1(new_n741), .A2(KEYINPUT87), .A3(G29), .ZN(new_n742));
  AOI21_X1  g317(.A(KEYINPUT87), .B1(new_n741), .B2(G29), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n736), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  XOR2_X1   g319(.A(KEYINPUT88), .B(G2067), .Z(new_n745));
  OAI22_X1  g320(.A1(new_n733), .A2(new_n734), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n681), .A2(G21), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G168), .B2(new_n681), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n746), .B1(G1966), .B2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(G164), .A2(G29), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G27), .B2(G29), .ZN(new_n751));
  INV_X1    g326(.A(G2078), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT31), .B(G11), .Z(new_n754));
  INV_X1    g329(.A(G28), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n755), .B2(KEYINPUT30), .ZN(new_n756));
  OR2_X1    g331(.A1(new_n756), .A2(KEYINPUT93), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n756), .A2(KEYINPUT93), .ZN(new_n758));
  OR3_X1    g333(.A1(new_n755), .A2(KEYINPUT92), .A3(KEYINPUT30), .ZN(new_n759));
  OAI21_X1  g334(.A(KEYINPUT92), .B1(new_n755), .B2(KEYINPUT30), .ZN(new_n760));
  AND4_X1   g335(.A1(new_n757), .A2(new_n758), .A3(new_n759), .A4(new_n760), .ZN(new_n761));
  AOI211_X1 g336(.A(new_n754), .B(new_n761), .C1(new_n627), .C2(G29), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n753), .A2(new_n762), .ZN(new_n763));
  AND2_X1   g338(.A1(new_n698), .A2(G32), .ZN(new_n764));
  AND2_X1   g339(.A1(new_n472), .A2(G105), .ZN(new_n765));
  NAND3_X1  g340(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n766));
  XNOR2_X1  g341(.A(new_n766), .B(KEYINPUT26), .ZN(new_n767));
  AOI211_X1 g342(.A(new_n765), .B(new_n767), .C1(G129), .C2(new_n480), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n478), .A2(G141), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n769), .B(KEYINPUT90), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n764), .B1(new_n771), .B2(G29), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT27), .B(G1996), .ZN(new_n773));
  OAI22_X1  g348(.A1(new_n772), .A2(new_n773), .B1(new_n752), .B2(new_n751), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n681), .A2(G4), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(new_n607), .B2(new_n681), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n763), .B(new_n774), .C1(new_n776), .C2(G1348), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n733), .A2(new_n734), .ZN(new_n778));
  NAND2_X1  g353(.A1(new_n726), .A2(new_n727), .ZN(new_n779));
  OR2_X1    g354(.A1(new_n748), .A2(G1966), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n744), .A2(new_n745), .ZN(new_n781));
  AND4_X1   g356(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n781), .ZN(new_n782));
  OR2_X1    g357(.A1(new_n776), .A2(G1348), .ZN(new_n783));
  NAND4_X1  g358(.A1(new_n749), .A2(new_n777), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n698), .A2(G33), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT25), .Z(new_n787));
  INV_X1    g362(.A(G139), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n474), .B2(new_n788), .ZN(new_n789));
  NAND3_X1  g364(.A1(new_n462), .A2(new_n468), .A3(G127), .ZN(new_n790));
  INV_X1    g365(.A(G115), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n791), .B2(new_n464), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n789), .B1(new_n792), .B2(G2105), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n785), .B1(new_n793), .B2(new_n698), .ZN(new_n794));
  XOR2_X1   g369(.A(new_n794), .B(G2072), .Z(new_n795));
  INV_X1    g370(.A(KEYINPUT24), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G34), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n698), .B1(new_n796), .B2(G34), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(KEYINPUT89), .ZN(new_n799));
  AOI21_X1  g374(.A(new_n799), .B1(KEYINPUT89), .B2(new_n798), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n800), .B1(G160), .B2(G29), .ZN(new_n801));
  AOI22_X1  g376(.A1(new_n772), .A2(new_n773), .B1(G2084), .B2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n795), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT91), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n681), .A2(G19), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n805), .B1(new_n541), .B2(new_n681), .ZN(new_n806));
  NOR2_X1   g381(.A1(new_n806), .A2(G1341), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(G1341), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n801), .A2(G2084), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT94), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NOR4_X1   g386(.A1(new_n784), .A2(new_n804), .A3(new_n807), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n731), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT97), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g390(.A1(new_n731), .A2(KEYINPUT97), .A3(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n717), .A2(new_n817), .ZN(G150));
  INV_X1    g393(.A(G150), .ZN(G311));
  NAND2_X1  g394(.A1(new_n607), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  INV_X1    g396(.A(G93), .ZN(new_n822));
  INV_X1    g397(.A(G55), .ZN(new_n823));
  OAI22_X1  g398(.A1(new_n510), .A2(new_n822), .B1(new_n512), .B2(new_n823), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n503), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  NOR2_X1   g400(.A1(new_n825), .A2(new_n504), .ZN(new_n826));
  OR2_X1    g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n541), .A2(new_n827), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n827), .A2(KEYINPUT98), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n824), .A2(new_n826), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT98), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(new_n540), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  XOR2_X1   g410(.A(new_n821), .B(new_n835), .Z(new_n836));
  INV_X1    g411(.A(KEYINPUT39), .ZN(new_n837));
  AOI21_X1  g412(.A(G860), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  OR2_X1    g415(.A1(new_n829), .A2(new_n832), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n841), .A2(G860), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(KEYINPUT37), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n840), .A2(new_n843), .ZN(G145));
  NAND2_X1  g419(.A1(new_n480), .A2(G130), .ZN(new_n845));
  OR2_X1    g420(.A1(G106), .A2(G2105), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n846), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G142), .B2(new_n478), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n615), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n850), .A2(new_n704), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n850), .A2(new_n704), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n793), .B(new_n771), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(new_n741), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n856), .B(G164), .ZN(new_n857));
  XNOR2_X1  g432(.A(KEYINPUT100), .B(KEYINPUT101), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n857), .B(new_n858), .Z(new_n859));
  INV_X1    g434(.A(new_n854), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n851), .A2(new_n860), .A3(new_n852), .ZN(new_n861));
  AND3_X1   g436(.A1(new_n855), .A2(new_n859), .A3(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n859), .B1(new_n855), .B2(new_n861), .ZN(new_n863));
  XNOR2_X1  g438(.A(G160), .B(G162), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n864), .B(new_n627), .Z(new_n865));
  OR3_X1    g440(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(G37), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n865), .B1(new_n862), .B2(new_n863), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  OR2_X1    g444(.A1(new_n869), .A2(KEYINPUT102), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(KEYINPUT102), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g448(.A(G868), .ZN(new_n874));
  NAND2_X1  g449(.A1(new_n841), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n600), .B(G299), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(KEYINPUT103), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n600), .B(new_n604), .ZN(new_n878));
  INV_X1    g453(.A(KEYINPUT41), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n876), .A2(KEYINPUT41), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n835), .B(new_n610), .ZN(new_n883));
  MUX2_X1   g458(.A(new_n877), .B(new_n882), .S(new_n883), .Z(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G305), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(new_n574), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(KEYINPUT42), .Z(new_n888));
  XNOR2_X1  g463(.A(new_n884), .B(new_n888), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n875), .B1(new_n889), .B2(new_n874), .ZN(G295));
  OAI21_X1  g465(.A(new_n875), .B1(new_n889), .B2(new_n874), .ZN(G331));
  NOR2_X1   g466(.A1(G301), .A2(G286), .ZN(new_n892));
  NOR2_X1   g467(.A1(G168), .A2(G171), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n835), .A2(new_n894), .ZN(new_n895));
  OAI211_X1 g470(.A(new_n828), .B(new_n834), .C1(new_n892), .C2(new_n893), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n897), .A2(new_n882), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n895), .A2(new_n878), .A3(new_n896), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n887), .ZN(new_n901));
  INV_X1    g476(.A(new_n887), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n901), .A2(new_n867), .A3(new_n903), .ZN(new_n904));
  XOR2_X1   g479(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n904), .A2(new_n906), .ZN(new_n907));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n880), .A2(KEYINPUT105), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n897), .A2(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT105), .B1(new_n880), .B2(new_n881), .ZN(new_n911));
  OAI221_X1 g486(.A(new_n887), .B1(new_n877), .B2(new_n897), .C1(new_n910), .C2(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n912), .A2(new_n867), .A3(new_n903), .A4(new_n905), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n907), .A2(new_n908), .A3(new_n913), .ZN(new_n914));
  OR2_X1    g489(.A1(new_n904), .A2(new_n906), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n887), .B1(new_n897), .B2(new_n877), .ZN(new_n917));
  OAI211_X1 g492(.A(new_n867), .B(new_n903), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n918), .A2(KEYINPUT43), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n918), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n915), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n914), .B1(new_n923), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g499(.A1(G303), .A2(G8), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT55), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n925), .B(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n494), .A2(new_n496), .ZN(new_n929));
  INV_X1    g504(.A(new_n491), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g506(.A(G1384), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n931), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G40), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n471), .A2(new_n934), .A3(new_n476), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT45), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n936), .B1(G164), .B2(G1384), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n933), .A2(new_n935), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(G1971), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  INV_X1    g516(.A(new_n476), .ZN(new_n942));
  AND2_X1   g517(.A1(new_n469), .A2(new_n470), .ZN(new_n943));
  OAI211_X1 g518(.A(G40), .B(new_n942), .C1(new_n943), .C2(new_n459), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT50), .ZN(new_n945));
  NOR2_X1   g520(.A1(G164), .A2(G1384), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT110), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n948), .B1(new_n931), .B2(new_n932), .ZN(new_n949));
  NOR3_X1   g524(.A1(G164), .A2(KEYINPUT110), .A3(G1384), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT50), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n947), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g527(.A(G2090), .B1(new_n952), .B2(KEYINPUT115), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n931), .A2(new_n948), .A3(new_n932), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT110), .B1(G164), .B2(G1384), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n945), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n931), .A2(new_n932), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n935), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n958));
  OR3_X1    g533(.A1(new_n956), .A2(new_n958), .A3(KEYINPUT115), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n941), .B1(new_n953), .B2(new_n959), .ZN(new_n960));
  INV_X1    g535(.A(G8), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n928), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n945), .B1(new_n931), .B2(new_n932), .ZN(new_n963));
  NOR2_X1   g538(.A1(new_n963), .A2(new_n944), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n954), .A2(new_n955), .A3(new_n945), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n964), .A2(new_n965), .A3(new_n727), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n966), .A2(new_n940), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT111), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n966), .A2(KEYINPUT111), .A3(new_n940), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n969), .A2(new_n927), .A3(G8), .A4(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT49), .ZN(new_n972));
  NAND2_X1  g547(.A1(G305), .A2(G1981), .ZN(new_n973));
  INV_X1    g548(.A(G1981), .ZN(new_n974));
  NAND4_X1  g549(.A1(new_n577), .A2(new_n580), .A3(new_n585), .A4(new_n974), .ZN(new_n975));
  NAND2_X1  g550(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT113), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AOI211_X1 g553(.A(KEYINPUT113), .B(KEYINPUT49), .C1(new_n973), .C2(new_n975), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n954), .A2(new_n935), .A3(new_n955), .ZN(new_n981));
  INV_X1    g556(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n961), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n574), .A2(G1976), .ZN(new_n984));
  NAND3_X1  g559(.A1(new_n984), .A2(G8), .A3(new_n981), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT112), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT52), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n985), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n574), .A2(KEYINPUT52), .A3(G1976), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n989), .B1(new_n985), .B2(new_n987), .ZN(new_n990));
  AOI22_X1  g565(.A1(new_n980), .A2(new_n983), .B1(new_n988), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(G2084), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n964), .A2(new_n992), .A3(new_n965), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n936), .B1(new_n949), .B2(new_n950), .ZN(new_n994));
  NOR3_X1   g569(.A1(G164), .A2(new_n936), .A3(G1384), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n944), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(G1966), .B1(new_n994), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(G8), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  NOR2_X1   g573(.A1(new_n998), .A2(G286), .ZN(new_n999));
  NAND4_X1  g574(.A1(new_n962), .A2(new_n971), .A3(new_n991), .A4(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT63), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT116), .ZN(new_n1003));
  AND2_X1   g578(.A1(new_n970), .A2(G8), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n927), .B1(new_n1004), .B2(new_n969), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n976), .A2(new_n977), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(KEYINPUT49), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n976), .A2(new_n977), .A3(new_n972), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n1007), .A2(new_n983), .A3(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n988), .A2(new_n990), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1003), .B1(new_n1005), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n970), .A2(G8), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT111), .B1(new_n966), .B2(new_n940), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n928), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n991), .A2(new_n1015), .A3(KEYINPUT116), .ZN(new_n1016));
  AND3_X1   g591(.A1(new_n999), .A2(new_n971), .A3(KEYINPUT63), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n1012), .A2(new_n1016), .A3(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1002), .A2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n722), .B1(new_n956), .B2(new_n958), .ZN(new_n1020));
  XNOR2_X1  g595(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1021));
  XNOR2_X1  g596(.A(new_n1021), .B(G2072), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n996), .A2(new_n937), .A3(new_n1022), .ZN(new_n1023));
  OR2_X1    g598(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1024));
  NAND2_X1  g599(.A1(KEYINPUT117), .A2(KEYINPUT57), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n559), .A2(new_n564), .A3(new_n1024), .A4(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(G299), .A2(KEYINPUT117), .A3(KEYINPUT57), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(G1348), .B1(new_n964), .B2(new_n965), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  NOR2_X1   g605(.A1(new_n981), .A2(G2067), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n600), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g608(.A1(new_n1020), .A2(new_n1023), .B1(new_n1027), .B2(new_n1026), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1028), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT61), .ZN(new_n1036));
  AND4_X1   g611(.A1(new_n1020), .A2(new_n1023), .A3(new_n1026), .A4(new_n1027), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1036), .B1(new_n1037), .B2(new_n1034), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n1032), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT60), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n1040), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1039), .A2(new_n607), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1020), .A2(new_n1023), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1027), .A2(new_n1026), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1045), .A2(KEYINPUT61), .A3(new_n1028), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1030), .A2(KEYINPUT60), .A3(new_n1032), .A4(new_n600), .ZN(new_n1047));
  NAND4_X1  g622(.A1(new_n1038), .A2(new_n1042), .A3(new_n1046), .A4(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1049));
  NOR2_X1   g624(.A1(KEYINPUT121), .A2(KEYINPUT59), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT120), .ZN(new_n1051));
  XOR2_X1   g626(.A(KEYINPUT58), .B(G1341), .Z(new_n1052));
  AND3_X1   g627(.A1(new_n981), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1051), .B1(new_n981), .B2(new_n1052), .ZN(new_n1054));
  XNOR2_X1  g629(.A(KEYINPUT119), .B(G1996), .ZN(new_n1055));
  NOR2_X1   g630(.A1(new_n938), .A2(new_n1055), .ZN(new_n1056));
  NOR3_X1   g631(.A1(new_n1053), .A2(new_n1054), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(new_n541), .ZN(new_n1058));
  OAI21_X1  g633(.A(new_n1050), .B1(new_n1057), .B2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(new_n1050), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n938), .A2(new_n1055), .ZN(new_n1061));
  AND2_X1   g636(.A1(new_n981), .A2(new_n1052), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1061), .B1(new_n1062), .B2(new_n1051), .ZN(new_n1063));
  OAI211_X1 g638(.A(new_n541), .B(new_n1060), .C1(new_n1063), .C2(new_n1053), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1049), .B1(new_n1059), .B2(new_n1064), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1035), .B1(new_n1048), .B2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(G286), .A2(G8), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT122), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT51), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n998), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT45), .B1(new_n954), .B2(new_n955), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n933), .A2(new_n935), .ZN(new_n1073));
  NOR2_X1   g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n964), .A2(new_n965), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1074), .A2(G1966), .B1(new_n1075), .B2(G2084), .ZN(new_n1076));
  OAI211_X1 g651(.A(G8), .B(new_n1069), .C1(new_n1076), .C2(G286), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1076), .A2(G8), .A3(G286), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1071), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n954), .A2(new_n955), .A3(new_n945), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n935), .B1(new_n946), .B2(new_n945), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n734), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND4_X1  g657(.A1(new_n933), .A2(new_n935), .A3(new_n937), .A4(new_n752), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n1084));
  NAND2_X1  g659(.A1(new_n1083), .A2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1084), .A2(G2078), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n933), .A2(new_n935), .A3(new_n937), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT123), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  OAI21_X1  g665(.A(G171), .B1(new_n1086), .B2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n994), .A2(new_n996), .A3(new_n1087), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n1082), .A2(new_n1092), .A3(G301), .A4(new_n1085), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1093), .A2(KEYINPUT124), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1075), .A2(new_n734), .B1(new_n1084), .B2(new_n1083), .ZN(new_n1095));
  INV_X1    g670(.A(KEYINPUT124), .ZN(new_n1096));
  NAND4_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(G301), .A4(new_n1092), .ZN(new_n1097));
  NAND4_X1  g672(.A1(new_n1091), .A2(new_n1094), .A3(KEYINPUT54), .A4(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  NAND4_X1  g674(.A1(new_n996), .A2(new_n1089), .A3(new_n937), .A4(new_n1087), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1088), .A2(KEYINPUT123), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1095), .A2(new_n1102), .A3(G301), .ZN(new_n1103));
  AOI21_X1  g678(.A(G301), .B1(new_n1095), .B2(new_n1092), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1099), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  AND3_X1   g680(.A1(new_n1079), .A2(new_n1098), .A3(new_n1105), .ZN(new_n1106));
  AND3_X1   g681(.A1(new_n962), .A2(new_n971), .A3(new_n991), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1066), .A2(new_n1106), .A3(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n983), .ZN(new_n1109));
  NOR2_X1   g684(.A1(G288), .A2(G1976), .ZN(new_n1110));
  OAI21_X1  g685(.A(new_n1110), .B1(new_n978), .B2(new_n979), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n1109), .B1(new_n1111), .B2(new_n975), .ZN(new_n1112));
  INV_X1    g687(.A(new_n1112), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n1113), .B(KEYINPUT114), .C1(new_n971), .C2(new_n1011), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1011), .A2(new_n971), .ZN(new_n1116));
  OAI21_X1  g691(.A(new_n1115), .B1(new_n1116), .B2(new_n1112), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1114), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1019), .A2(new_n1108), .A3(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT125), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1019), .A2(new_n1108), .A3(new_n1118), .A4(KEYINPUT125), .ZN(new_n1122));
  OR2_X1    g697(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1079), .A2(KEYINPUT62), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1123), .A2(new_n1107), .A3(new_n1104), .A4(new_n1124), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1121), .A2(new_n1122), .A3(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(KEYINPUT107), .B1(new_n944), .B2(new_n937), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT107), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n935), .A2(new_n957), .A3(new_n1128), .A4(new_n936), .ZN(new_n1129));
  AND2_X1   g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  NAND3_X1  g705(.A1(new_n1130), .A2(G1996), .A3(new_n771), .ZN(new_n1131));
  XOR2_X1   g706(.A(new_n1131), .B(KEYINPUT108), .Z(new_n1132));
  INV_X1    g707(.A(G2067), .ZN(new_n1133));
  XNOR2_X1  g708(.A(new_n741), .B(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1134), .B1(new_n771), .B2(G1996), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1132), .B1(new_n1130), .B2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n704), .B(new_n707), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n1137), .B(KEYINPUT109), .Z(new_n1138));
  NAND2_X1  g713(.A1(new_n1138), .A2(new_n1130), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  XNOR2_X1  g715(.A(G290), .B(G1986), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n1130), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1126), .A2(new_n1142), .ZN(new_n1143));
  INV_X1    g718(.A(G1996), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1130), .A2(new_n1144), .ZN(new_n1145));
  XNOR2_X1  g720(.A(new_n1145), .B(KEYINPUT46), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1130), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n1134), .A2(new_n770), .A3(new_n768), .ZN(new_n1148));
  OAI21_X1  g723(.A(new_n1146), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(KEYINPUT47), .ZN(new_n1150));
  NOR3_X1   g725(.A1(new_n1147), .A2(G1986), .A3(G290), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT48), .ZN(new_n1152));
  OAI21_X1  g727(.A(new_n1150), .B1(new_n1140), .B2(new_n1152), .ZN(new_n1153));
  AND2_X1   g728(.A1(new_n705), .A2(new_n707), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1136), .A2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g730(.A1(new_n856), .A2(new_n1133), .ZN(new_n1156));
  AOI21_X1  g731(.A(new_n1147), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  OR3_X1    g732(.A1(new_n1153), .A2(new_n1157), .A3(KEYINPUT126), .ZN(new_n1158));
  OAI21_X1  g733(.A(KEYINPUT126), .B1(new_n1153), .B2(new_n1157), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1143), .A2(new_n1160), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g736(.A(KEYINPUT127), .ZN(new_n1163));
  INV_X1    g737(.A(G319), .ZN(new_n1164));
  NOR2_X1   g738(.A1(G227), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g739(.A1(new_n679), .A2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g740(.A(new_n1163), .B1(new_n1166), .B2(G401), .ZN(new_n1167));
  OR2_X1    g741(.A1(new_n644), .A2(new_n645), .ZN(new_n1168));
  NAND4_X1  g742(.A1(new_n1168), .A2(KEYINPUT127), .A3(new_n679), .A4(new_n1165), .ZN(new_n1169));
  AOI22_X1  g743(.A1(new_n870), .A2(new_n871), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g744(.A1(new_n907), .A2(new_n913), .ZN(new_n1171));
  NAND2_X1  g745(.A1(new_n1170), .A2(new_n1171), .ZN(G225));
  INV_X1    g746(.A(G225), .ZN(G308));
endmodule


